//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n572, new_n574,
    new_n575, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT67), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  XOR2_X1   g014(.A(KEYINPUT68), .B(G69), .Z(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  AND2_X1   g018(.A1(G2072), .A2(G2078), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT69), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR3_X1   g028(.A1(G218), .A2(G219), .A3(G221), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n437), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT71), .ZN(new_n456));
  XNOR2_X1  g031(.A(KEYINPUT70), .B(KEYINPUT2), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n456), .B(new_n457), .ZN(new_n458));
  OR4_X1    g033(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  NAND2_X1  g036(.A1(new_n458), .A2(G2106), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT72), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT72), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n466), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT73), .B1(new_n469), .B2(KEYINPUT3), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT73), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(new_n467), .A3(G2104), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n478), .A2(new_n480), .A3(new_n481), .A4(new_n470), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT74), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n483), .A2(new_n484), .A3(G137), .ZN(new_n485));
  INV_X1    g060(.A(G137), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT74), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n469), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G101), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n477), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G160));
  NAND2_X1  g067(.A1(new_n483), .A2(G136), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT75), .B1(G100), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NOR3_X1   g070(.A1(KEYINPUT75), .A2(G100), .A3(G2105), .ZN(new_n496));
  OAI221_X1 g071(.A(G2104), .B1(G112), .B2(new_n481), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G124), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n478), .A2(new_n480), .A3(new_n470), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n493), .B(new_n497), .C1(new_n498), .C2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G162));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT76), .ZN(new_n504));
  OR3_X1    g079(.A1(new_n504), .A2(new_n481), .A3(G114), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n481), .B2(G114), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n499), .A2(G2105), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G126), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n510));
  INV_X1    g085(.A(G138), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n511), .A2(G2105), .ZN(new_n512));
  INV_X1    g087(.A(new_n474), .ZN(new_n513));
  AOI21_X1  g088(.A(KEYINPUT72), .B1(new_n468), .B2(new_n470), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n510), .B(new_n512), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n478), .A2(new_n480), .A3(new_n470), .A4(new_n512), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n516), .A2(KEYINPUT77), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT4), .B1(new_n516), .B2(KEYINPUT77), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n509), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(G164));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G62), .ZN(new_n526));
  NAND2_X1  g101(.A1(G75), .A2(G543), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT79), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n522), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT80), .ZN(new_n530));
  AND2_X1   g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  NOR2_X1   g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n529), .A2(KEYINPUT80), .B1(G50), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G88), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n523), .A2(new_n524), .ZN(new_n538));
  OAI21_X1  g113(.A(KEYINPUT78), .B1(new_n538), .B2(new_n533), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT78), .ZN(new_n540));
  OAI221_X1 g115(.A(new_n540), .B1(new_n523), .B2(new_n524), .C1(new_n532), .C2(new_n531), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n530), .B(new_n536), .C1(new_n537), .C2(new_n542), .ZN(G303));
  INV_X1    g118(.A(G303), .ZN(G166));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  INV_X1    g121(.A(G89), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(KEYINPUT81), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT81), .ZN(new_n550));
  OAI211_X1 g125(.A(new_n550), .B(new_n546), .C1(new_n542), .C2(new_n547), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n538), .A2(new_n522), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n552), .A2(G63), .B1(new_n535), .B2(G51), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n549), .A2(new_n551), .A3(new_n553), .ZN(G286));
  INV_X1    g129(.A(G286), .ZN(G168));
  AOI22_X1  g130(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n522), .ZN(new_n557));
  INV_X1    g132(.A(G52), .ZN(new_n558));
  INV_X1    g133(.A(new_n535), .ZN(new_n559));
  INV_X1    g134(.A(G90), .ZN(new_n560));
  OAI221_X1 g135(.A(new_n557), .B1(new_n558), .B2(new_n559), .C1(new_n542), .C2(new_n560), .ZN(G301));
  INV_X1    g136(.A(G301), .ZN(G171));
  AOI22_X1  g137(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(new_n522), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(KEYINPUT82), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n564), .A2(KEYINPUT82), .B1(G43), .B2(new_n535), .ZN(new_n566));
  INV_X1    g141(.A(new_n542), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G81), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT83), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND4_X1  g150(.A1(G319), .A2(G483), .A3(G661), .A4(new_n575), .ZN(G188));
  NAND2_X1  g151(.A1(new_n535), .A2(G53), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT9), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n567), .A2(G91), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n522), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(G299));
  OAI21_X1  g157(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n583));
  XOR2_X1   g158(.A(new_n583), .B(KEYINPUT85), .Z(new_n584));
  NAND2_X1  g159(.A1(new_n567), .A2(G87), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n535), .A2(G49), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT84), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n584), .A2(new_n585), .A3(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n538), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(new_n535), .B2(G48), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n539), .A2(new_n541), .A3(G86), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n567), .A2(G85), .ZN(new_n597));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G60), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n538), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(new_n535), .B2(G47), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n567), .A2(G92), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n538), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(new_n535), .B2(G54), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n603), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n603), .B1(new_n612), .B2(G868), .ZN(G321));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(G299), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G168), .B2(new_n615), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(G168), .B2(new_n615), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n569), .A2(new_n615), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n611), .A2(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n615), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g199(.A(new_n489), .B1(new_n513), .B2(new_n514), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  AND2_X1   g202(.A1(new_n627), .A2(KEYINPUT13), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n627), .A2(KEYINPUT13), .ZN(new_n629));
  OAI22_X1  g204(.A1(new_n628), .A2(new_n629), .B1(KEYINPUT87), .B2(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(KEYINPUT87), .A2(G2100), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n630), .B(new_n631), .Z(new_n632));
  INV_X1    g207(.A(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n481), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI22_X1  g210(.A1(new_n500), .A2(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(G135), .B2(new_n483), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT88), .ZN(new_n638));
  INV_X1    g213(.A(G2096), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n632), .A2(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  OAI21_X1  g228(.A(G14), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT89), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n652), .A2(KEYINPUT89), .A3(new_n653), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n661), .B(KEYINPUT17), .Z(new_n665));
  INV_X1    g240(.A(new_n660), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n666), .A2(new_n662), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n664), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n662), .B1(new_n661), .B2(KEYINPUT90), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(KEYINPUT90), .B2(new_n661), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n670), .A2(KEYINPUT91), .A3(new_n666), .ZN(new_n671));
  INV_X1    g246(.A(new_n662), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n671), .B1(new_n672), .B2(new_n665), .ZN(new_n673));
  AOI21_X1  g248(.A(KEYINPUT91), .B1(new_n670), .B2(new_n666), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n668), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n639), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT92), .B(G2100), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n682), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n680), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n680), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n689), .B(new_n690), .Z(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  OR2_X1    g271(.A1(G4), .A2(G16), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n611), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G1348), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT96), .B(KEYINPUT28), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT97), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G26), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n703), .B(new_n705), .Z(new_n706));
  INV_X1    g281(.A(G128), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n481), .A2(G116), .ZN(new_n708));
  OAI21_X1  g283(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n709));
  OAI22_X1  g284(.A1(new_n500), .A2(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n483), .A2(G140), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n706), .B1(new_n712), .B2(new_n704), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G2067), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n698), .A2(G20), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT23), .Z(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G299), .B2(G16), .ZN(new_n717));
  INV_X1    g292(.A(G1956), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NOR3_X1   g294(.A1(new_n701), .A2(new_n714), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(G168), .A2(new_n698), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n698), .B2(G21), .ZN(new_n722));
  INV_X1    g297(.A(G1966), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  NOR2_X1   g300(.A1(G29), .A2(G35), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G162), .B2(G29), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT29), .B(G2090), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n698), .A2(G19), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n569), .B2(G16), .ZN(new_n731));
  INV_X1    g306(.A(G1341), .ZN(new_n732));
  OAI221_X1 g307(.A(new_n729), .B1(new_n731), .B2(new_n732), .C1(new_n704), .C2(new_n638), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n725), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n698), .A2(G5), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G171), .B2(new_n698), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(G1961), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT103), .B(KEYINPUT31), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G11), .ZN(new_n739));
  INV_X1    g314(.A(G28), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(KEYINPUT30), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT104), .ZN(new_n742));
  AOI21_X1  g317(.A(G29), .B1(new_n740), .B2(KEYINPUT30), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI211_X1 g319(.A(new_n739), .B(new_n744), .C1(new_n736), .C2(G1961), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n731), .A2(new_n732), .B1(new_n727), .B2(new_n728), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT24), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n747), .A2(G34), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(G34), .ZN(new_n749));
  AOI21_X1  g324(.A(G29), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n491), .B2(G29), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2084), .ZN(new_n752));
  AND4_X1   g327(.A1(new_n737), .A2(new_n745), .A3(new_n746), .A4(new_n752), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n720), .A2(new_n724), .A3(new_n734), .A4(new_n753), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n704), .A2(G32), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n483), .A2(G141), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT26), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n759), .A2(new_n760), .B1(G105), .B2(new_n489), .ZN(new_n761));
  AND3_X1   g336(.A1(new_n499), .A2(G129), .A3(G2105), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT101), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n756), .B(new_n761), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT102), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n755), .B1(new_n768), .B2(G29), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT27), .B(G1996), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n704), .A2(G33), .ZN(new_n772));
  OAI21_X1  g347(.A(G127), .B1(new_n513), .B2(new_n514), .ZN(new_n773));
  INV_X1    g348(.A(G115), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(new_n469), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n481), .B1(new_n775), .B2(KEYINPUT98), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(KEYINPUT98), .B2(new_n775), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT25), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n483), .B2(G139), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n772), .B1(new_n781), .B2(new_n704), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G2072), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(KEYINPUT99), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(KEYINPUT99), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n769), .A2(new_n770), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n771), .A2(new_n784), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n782), .A2(G2072), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT100), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n704), .A2(G27), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT105), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n520), .B2(G29), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2078), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT106), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n754), .A2(new_n787), .A3(new_n789), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n698), .A2(G23), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n584), .A2(new_n588), .A3(new_n585), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n698), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT33), .B(G1976), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(KEYINPUT94), .ZN(new_n801));
  NOR2_X1   g376(.A1(G6), .A2(G16), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n595), .B2(G16), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT32), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1981), .ZN(new_n805));
  NOR2_X1   g380(.A1(G16), .A2(G22), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G166), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1971), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n800), .A2(KEYINPUT94), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n801), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT34), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n809), .A2(new_n801), .A3(new_n813), .A4(new_n810), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n508), .A2(G119), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT93), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n817));
  INV_X1    g392(.A(G107), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(G2105), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n483), .B2(G131), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  MUX2_X1   g396(.A(G25), .B(new_n821), .S(G29), .Z(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n822), .A2(new_n824), .ZN(new_n826));
  MUX2_X1   g401(.A(G24), .B(G290), .S(G16), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1986), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n812), .A2(new_n814), .A3(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT95), .B(KEYINPUT36), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n831), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n812), .A2(new_n833), .A3(new_n814), .A4(new_n829), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n795), .A2(new_n832), .A3(new_n834), .ZN(G150));
  INV_X1    g410(.A(KEYINPUT107), .ZN(new_n836));
  XNOR2_X1  g411(.A(G150), .B(new_n836), .ZN(G311));
  NAND2_X1  g412(.A1(new_n612), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n535), .A2(G55), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT108), .B(G93), .ZN(new_n842));
  OAI221_X1 g417(.A(new_n840), .B1(new_n841), .B2(new_n522), .C1(new_n542), .C2(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n569), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n569), .A2(new_n843), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n839), .B(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n849), .A2(new_n850), .A3(G860), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n843), .A2(G860), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n851), .A2(new_n853), .ZN(G145));
  XNOR2_X1  g429(.A(KEYINPUT111), .B(G37), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n515), .B(KEYINPUT109), .C1(new_n517), .C2(new_n518), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n480), .A2(new_n470), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT77), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n858), .A2(new_n859), .A3(new_n478), .A4(new_n512), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n516), .A2(KEYINPUT77), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(KEYINPUT4), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT109), .B1(new_n862), .B2(new_n515), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n509), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n781), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n712), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n767), .B(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n868), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(G130), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n481), .A2(G118), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  OAI22_X1  g449(.A1(new_n500), .A2(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(G142), .B2(new_n483), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(new_n627), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n821), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT110), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n871), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n638), .B(new_n501), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G160), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT110), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n870), .A2(new_n869), .A3(new_n883), .A4(new_n878), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n880), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n882), .B1(new_n880), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n855), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g463(.A1(new_n843), .A2(new_n615), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n846), .B(KEYINPUT112), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n622), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n611), .A2(G299), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n611), .A2(G299), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT41), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n896), .B1(new_n894), .B2(new_n891), .ZN(new_n897));
  XOR2_X1   g472(.A(G290), .B(KEYINPUT113), .Z(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(G288), .ZN(new_n899));
  XNOR2_X1  g474(.A(G303), .B(G305), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n898), .B(new_n797), .ZN(new_n902));
  INV_X1    g477(.A(new_n900), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT42), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT114), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n902), .A2(new_n903), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n899), .A2(new_n900), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n901), .A2(new_n904), .A3(KEYINPUT114), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n905), .B1(new_n911), .B2(KEYINPUT42), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n897), .B(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n889), .B1(new_n913), .B2(new_n615), .ZN(G295));
  OAI21_X1  g489(.A(new_n889), .B1(new_n913), .B2(new_n615), .ZN(G331));
  NAND2_X1  g490(.A1(G168), .A2(G171), .ZN(new_n916));
  NAND2_X1  g491(.A1(G286), .A2(G301), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n846), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT115), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n916), .A2(new_n844), .A3(new_n845), .A4(new_n917), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n847), .A2(KEYINPUT115), .A3(new_n917), .A4(new_n916), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n894), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT116), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n919), .A2(new_n921), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n895), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(KEYINPUT116), .A3(new_n925), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n932), .B2(new_n911), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n901), .A2(new_n904), .A3(KEYINPUT114), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT114), .B1(new_n901), .B2(new_n904), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n936), .A2(new_n928), .A3(new_n930), .A4(new_n931), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT43), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n855), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n894), .B(new_n940), .ZN(new_n941));
  OAI22_X1  g516(.A1(new_n941), .A2(new_n924), .B1(new_n894), .B2(new_n929), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n939), .B1(new_n911), .B2(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n937), .A2(new_n943), .A3(KEYINPUT43), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT44), .B1(new_n938), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n933), .B2(new_n937), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n937), .A2(new_n943), .A3(new_n947), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n945), .A2(new_n950), .ZN(G397));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT45), .B1(new_n864), .B2(new_n952), .ZN(new_n953));
  AND4_X1   g528(.A1(G40), .A2(new_n477), .A3(new_n488), .A4(new_n490), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT117), .B1(new_n955), .B2(G1996), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n957));
  INV_X1    g532(.A(new_n507), .ZN(new_n958));
  INV_X1    g533(.A(G126), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n958), .B1(new_n500), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n519), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n960), .B1(new_n962), .B2(new_n856), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n957), .B1(new_n963), .B2(G1384), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n477), .A2(new_n488), .A3(G40), .A4(new_n490), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT117), .ZN(new_n967));
  INV_X1    g542(.A(G1996), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n956), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT46), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n970), .B(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n712), .B(G2067), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n966), .B1(new_n768), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT47), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n970), .A2(new_n767), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n974), .B1(new_n768), .B2(G1996), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n978), .B1(new_n955), .B2(new_n979), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n980), .A2(new_n821), .A3(new_n824), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n867), .A2(G2067), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n966), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n821), .B(new_n824), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n980), .B1(new_n966), .B2(new_n984), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n955), .A2(G1986), .A3(G290), .ZN(new_n986));
  XOR2_X1   g561(.A(new_n986), .B(KEYINPUT48), .Z(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n977), .A2(new_n983), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT63), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n512), .A2(new_n510), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n992), .B1(new_n473), .B2(new_n474), .ZN(new_n993));
  AND4_X1   g568(.A1(new_n478), .A2(new_n480), .A3(new_n470), .A4(new_n512), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n510), .B1(new_n994), .B2(new_n859), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n993), .B1(new_n995), .B2(new_n861), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT45), .B(new_n952), .C1(new_n996), .C2(new_n960), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT119), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n520), .A2(KEYINPUT119), .A3(KEYINPUT45), .A4(new_n952), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n954), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n723), .B1(new_n1001), .B2(new_n953), .ZN(new_n1002));
  INV_X1    g577(.A(G2084), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n520), .A2(new_n952), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n965), .B1(new_n1004), .B2(KEYINPUT50), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n864), .A2(new_n952), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1003), .B(new_n1005), .C1(new_n1006), .C2(KEYINPUT50), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1002), .A2(new_n1007), .ZN(new_n1008));
  AND4_X1   g583(.A1(KEYINPUT120), .A2(new_n1008), .A3(G8), .A4(G168), .ZN(new_n1009));
  INV_X1    g584(.A(G8), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n1002), .B2(new_n1007), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT120), .B1(new_n1011), .B2(G168), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(G303), .A2(G8), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT55), .ZN(new_n1015));
  INV_X1    g590(.A(G1971), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n864), .A2(KEYINPUT45), .A3(new_n952), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1004), .A2(new_n957), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(new_n954), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n520), .A2(new_n1020), .A3(new_n952), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n954), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n1006), .B2(KEYINPUT50), .ZN(new_n1023));
  INV_X1    g598(.A(G2090), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n1016), .A2(new_n1019), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1015), .B1(new_n1025), .B2(new_n1010), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n962), .A2(new_n856), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1384), .B1(new_n1027), .B2(new_n509), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1010), .B1(new_n1028), .B2(new_n954), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n797), .A2(G1976), .ZN(new_n1030));
  INV_X1    g605(.A(G1976), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(G288), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1028), .A2(new_n954), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT118), .B(G1981), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n595), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1981), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1036), .B1(new_n1037), .B2(new_n595), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT49), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1036), .B(KEYINPUT49), .C1(new_n1037), .C2(new_n595), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1034), .A2(G8), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1033), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1015), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n965), .B1(new_n1028), .B2(KEYINPUT45), .ZN(new_n1048));
  AOI21_X1  g623(.A(G1971), .B1(new_n1048), .B2(new_n1018), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n963), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1384), .B1(new_n509), .B2(new_n519), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n954), .B1(new_n1051), .B2(new_n1020), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1050), .A2(G2090), .A3(new_n1052), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1047), .B(G8), .C1(new_n1049), .C2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1026), .A2(new_n1046), .A3(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n991), .B1(new_n1013), .B2(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1046), .A2(new_n1054), .ZN(new_n1057));
  OAI21_X1  g632(.A(G8), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n991), .B1(new_n1058), .B2(new_n1015), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1057), .B(new_n1059), .C1(new_n1009), .C2(new_n1012), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1062), .B(G8), .C1(new_n1008), .C2(G286), .ZN(new_n1063));
  NAND2_X1  g638(.A1(G286), .A2(G8), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT126), .B1(new_n1008), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT126), .ZN(new_n1067));
  AOI211_X1 g642(.A(new_n1067), .B(new_n1064), .C1(new_n1002), .C2(new_n1007), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1063), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1011), .A2(new_n1062), .A3(new_n1065), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT62), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n964), .A2(new_n954), .A3(new_n999), .A4(new_n1000), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1052), .B1(new_n1028), .B2(new_n1020), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1072), .A2(new_n723), .B1(new_n1073), .B2(new_n1003), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1067), .B1(new_n1074), .B2(new_n1064), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1008), .A2(KEYINPUT126), .A3(new_n1065), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT62), .ZN(new_n1078));
  OAI211_X1 g653(.A(KEYINPUT51), .B(new_n1064), .C1(new_n1074), .C2(new_n1010), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .A4(new_n1063), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1082));
  INV_X1    g657(.A(G1961), .ZN(new_n1083));
  OAI211_X1 g658(.A(KEYINPUT122), .B(new_n1005), .C1(new_n1006), .C2(KEYINPUT50), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1019), .B2(G2078), .ZN(new_n1087));
  INV_X1    g662(.A(G2078), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT53), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1085), .B(new_n1087), .C1(new_n1089), .C2(new_n1072), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G171), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1055), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1071), .A2(new_n1080), .A3(new_n1092), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1054), .A2(new_n1045), .A3(new_n1043), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1042), .A2(new_n1031), .A3(new_n797), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1036), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1094), .B1(new_n1029), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1061), .A2(new_n1093), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1082), .A2(new_n700), .A3(new_n1084), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1034), .A2(G2067), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(new_n611), .ZN(new_n1102));
  XOR2_X1   g677(.A(G299), .B(KEYINPUT57), .Z(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT56), .B(G2072), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1048), .A2(new_n1018), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT50), .B1(new_n963), .B2(G1384), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n965), .B1(new_n1051), .B2(new_n1020), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT121), .B1(new_n1108), .B2(new_n718), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n1110));
  AOI211_X1 g685(.A(new_n1110), .B(G1956), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1103), .B(new_n1105), .C1(new_n1109), .C2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1102), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1105), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1103), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n1112), .A3(KEYINPUT61), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT124), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1116), .A2(new_n1112), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT58), .B(G1341), .Z(new_n1124));
  NAND2_X1  g699(.A1(new_n1034), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1017), .A2(new_n968), .A3(new_n954), .A4(new_n1018), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1123), .B1(new_n1127), .B2(new_n570), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1123), .A3(new_n570), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  AOI211_X1 g707(.A(KEYINPUT123), .B(new_n569), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT59), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1116), .A2(new_n1112), .A3(new_n1136), .A4(KEYINPUT61), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1119), .A2(new_n1122), .A3(new_n1135), .A4(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1101), .A2(KEYINPUT60), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1099), .A2(KEYINPUT60), .A3(new_n1100), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n612), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1140), .A2(new_n1141), .A3(new_n611), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1101), .A2(KEYINPUT125), .A3(KEYINPUT60), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1139), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1117), .B1(new_n1138), .B2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1048), .A2(KEYINPUT53), .A3(new_n1088), .A4(new_n964), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1085), .A2(new_n1087), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(G171), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1151), .B(KEYINPUT54), .C1(G171), .C2(new_n1090), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1152), .A2(new_n1026), .A3(new_n1057), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1150), .A2(G171), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT54), .B1(new_n1155), .B2(new_n1091), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1153), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1098), .B1(new_n1148), .B2(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(G290), .B(G1986), .Z(new_n1159));
  OAI21_X1  g734(.A(new_n985), .B1(new_n955), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n990), .B1(new_n1158), .B2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g736(.A1(G227), .A2(new_n464), .ZN(new_n1163));
  OAI21_X1  g737(.A(KEYINPUT127), .B1(new_n1163), .B2(G401), .ZN(new_n1164));
  NAND2_X1  g738(.A1(new_n695), .A2(new_n1164), .ZN(new_n1165));
  NOR3_X1   g739(.A1(new_n1163), .A2(G401), .A3(KEYINPUT127), .ZN(new_n1166));
  NOR2_X1   g740(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g741(.A(new_n887), .B(new_n1167), .C1(new_n948), .C2(new_n949), .ZN(G225));
  INV_X1    g742(.A(G225), .ZN(G308));
endmodule


