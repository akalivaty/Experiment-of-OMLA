//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n531, new_n532, new_n534, new_n535, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n563, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n579, new_n580, new_n583,
    new_n585, new_n586, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1080, new_n1081, new_n1082,
    new_n1083;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G236), .A3(G238), .A4(G235), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  XNOR2_X1  g029(.A(G325), .B(KEYINPUT66), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G125), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT68), .ZN(new_n464));
  OAI21_X1  g039(.A(G2105), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G101), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n460), .A2(G2105), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n469), .B1(new_n470), .B2(G137), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n465), .A2(new_n471), .ZN(G160));
  OR2_X1    g047(.A1(G100), .A2(G2105), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n473), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G124), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n478), .B1(G136), .B2(new_n470), .ZN(G162));
  AND2_X1   g054(.A1(KEYINPUT70), .A2(G138), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n466), .B(new_n480), .C1(new_n458), .C2(new_n459), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT69), .B(G114), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(new_n466), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n466), .A2(KEYINPUT70), .A3(KEYINPUT4), .A4(G138), .ZN(new_n488));
  NAND2_X1  g063(.A1(G126), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(new_n475), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n483), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G164));
  INV_X1    g068(.A(G50), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT6), .A2(G651), .ZN(new_n495));
  NOR2_X1   g070(.A1(KEYINPUT6), .A2(G651), .ZN(new_n496));
  OR2_X1    g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G543), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G88), .ZN(new_n501));
  OAI22_X1  g076(.A1(new_n494), .A2(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n502), .A2(new_n505), .ZN(G166));
  NAND3_X1  g081(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n507));
  XNOR2_X1  g082(.A(new_n507), .B(KEYINPUT7), .ZN(new_n508));
  INV_X1    g083(.A(G89), .ZN(new_n509));
  INV_X1    g084(.A(G51), .ZN(new_n510));
  OAI221_X1 g085(.A(new_n508), .B1(new_n500), .B2(new_n509), .C1(new_n510), .C2(new_n498), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n499), .A2(G63), .A3(G651), .ZN(new_n512));
  XOR2_X1   g087(.A(new_n512), .B(KEYINPUT71), .Z(new_n513));
  NOR2_X1   g088(.A1(new_n511), .A2(new_n513), .ZN(G168));
  INV_X1    g089(.A(G90), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT72), .B(G52), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n515), .A2(new_n500), .B1(new_n498), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n499), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n518), .A2(new_n504), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n517), .A2(new_n519), .ZN(G301));
  INV_X1    g095(.A(G301), .ZN(G171));
  AOI22_X1  g096(.A1(new_n499), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n522), .A2(new_n504), .ZN(new_n523));
  XOR2_X1   g098(.A(new_n523), .B(KEYINPUT73), .Z(new_n524));
  INV_X1    g099(.A(new_n500), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n497), .A2(G543), .ZN(new_n526));
  AOI22_X1  g101(.A1(G81), .A2(new_n525), .B1(new_n526), .B2(G43), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G860), .ZN(G153));
  AND3_X1   g105(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G36), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT74), .ZN(G176));
  NAND2_X1  g108(.A1(G1), .A2(G3), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT8), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n531), .A2(new_n535), .ZN(G188));
  XNOR2_X1  g111(.A(KEYINPUT75), .B(G65), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n499), .A2(new_n537), .B1(G78), .B2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G91), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n538), .A2(new_n504), .B1(new_n500), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g115(.A(G53), .B(G543), .C1(new_n495), .C2(new_n496), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT9), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(G299));
  INV_X1    g120(.A(G168), .ZN(G286));
  INV_X1    g121(.A(G166), .ZN(G303));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n525), .B2(G87), .ZN(new_n549));
  INV_X1    g124(.A(G87), .ZN(new_n550));
  NOR3_X1   g125(.A1(new_n500), .A2(KEYINPUT76), .A3(new_n550), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n499), .A2(G74), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n526), .A2(G49), .B1(new_n553), .B2(G651), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(G288));
  INV_X1    g130(.A(G48), .ZN(new_n556));
  INV_X1    g131(.A(G86), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n556), .A2(new_n498), .B1(new_n500), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n499), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n504), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(G305));
  XOR2_X1   g137(.A(KEYINPUT77), .B(G47), .Z(new_n563));
  AOI22_X1  g138(.A1(G85), .A2(new_n525), .B1(new_n526), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n504), .B2(new_n565), .ZN(G290));
  NAND2_X1  g141(.A1(G301), .A2(G868), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n525), .A2(G92), .ZN(new_n568));
  XOR2_X1   g143(.A(new_n568), .B(KEYINPUT10), .Z(new_n569));
  NAND2_X1  g144(.A1(G79), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(new_n499), .ZN(new_n571));
  XOR2_X1   g146(.A(KEYINPUT78), .B(G66), .Z(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(G651), .A2(new_n573), .B1(new_n526), .B2(G54), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n567), .B1(new_n576), .B2(G868), .ZN(G284));
  OAI21_X1  g152(.A(new_n567), .B1(new_n576), .B2(G868), .ZN(G321));
  INV_X1    g153(.A(G868), .ZN(new_n579));
  NAND2_X1  g154(.A1(G299), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n580), .B1(new_n579), .B2(G168), .ZN(G297));
  OAI21_X1  g156(.A(new_n580), .B1(new_n579), .B2(G168), .ZN(G280));
  INV_X1    g157(.A(G559), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n576), .B1(new_n583), .B2(G860), .ZN(G148));
  NAND2_X1  g159(.A1(new_n528), .A2(new_n579), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n575), .A2(G559), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n586), .B2(new_n579), .ZN(G323));
  XNOR2_X1  g162(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g163(.A1(new_n470), .A2(G2104), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT12), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT13), .ZN(new_n591));
  INV_X1    g166(.A(G2100), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  INV_X1    g169(.A(new_n476), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G123), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n470), .A2(G135), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n466), .A2(G111), .ZN(new_n598));
  OAI21_X1  g173(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n596), .B(new_n597), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  XOR2_X1   g175(.A(new_n600), .B(G2096), .Z(new_n601));
  NAND3_X1  g176(.A1(new_n593), .A2(new_n594), .A3(new_n601), .ZN(G156));
  INV_X1    g177(.A(KEYINPUT14), .ZN(new_n603));
  XNOR2_X1  g178(.A(G2427), .B(G2438), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(G2430), .ZN(new_n605));
  XNOR2_X1  g180(.A(KEYINPUT15), .B(G2435), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(new_n606), .B2(new_n605), .ZN(new_n608));
  XNOR2_X1  g183(.A(G2451), .B(G2454), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT16), .ZN(new_n610));
  XNOR2_X1  g185(.A(G1341), .B(G1348), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n608), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(G2443), .B(G2446), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n615), .A2(G14), .A3(new_n616), .ZN(G401));
  XNOR2_X1  g192(.A(G2067), .B(G2678), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT79), .Z(new_n619));
  XNOR2_X1  g194(.A(G2072), .B(G2078), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT80), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(G2084), .B(G2090), .Z(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n620), .B(KEYINPUT17), .Z(new_n625));
  OAI211_X1 g200(.A(new_n622), .B(new_n624), .C1(new_n619), .C2(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n623), .A2(new_n618), .A3(new_n620), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT18), .Z(new_n628));
  NAND3_X1  g203(.A1(new_n619), .A2(new_n625), .A3(new_n623), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n626), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2096), .B(G2100), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(G227));
  XOR2_X1   g207(.A(G1971), .B(G1976), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT19), .ZN(new_n634));
  XOR2_X1   g209(.A(G1956), .B(G2474), .Z(new_n635));
  XOR2_X1   g210(.A(G1961), .B(G1966), .Z(new_n636));
  AND2_X1   g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT20), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n635), .A2(new_n636), .ZN(new_n640));
  NOR3_X1   g215(.A1(new_n634), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n634), .B2(new_n640), .ZN(new_n642));
  AND2_X1   g217(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT81), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1991), .B(G1996), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT82), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1981), .B(G1986), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(G229));
  MUX2_X1   g226(.A(G23), .B(G288), .S(G16), .Z(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT33), .B(G1976), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n652), .B(new_n653), .Z(new_n654));
  NOR2_X1   g229(.A1(G6), .A2(G16), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n561), .B2(G16), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT32), .B(G1981), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(G16), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(G22), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(G166), .B2(new_n660), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G1971), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  OR3_X1    g240(.A1(new_n654), .A2(KEYINPUT34), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(KEYINPUT34), .B1(new_n654), .B2(new_n665), .ZN(new_n667));
  MUX2_X1   g242(.A(G24), .B(G290), .S(G16), .Z(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(G1986), .Z(new_n669));
  INV_X1    g244(.A(G29), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(G25), .ZN(new_n671));
  OR2_X1    g246(.A1(G95), .A2(G2105), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n672), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n475), .A2(new_n466), .ZN(new_n674));
  INV_X1    g249(.A(G131), .ZN(new_n675));
  INV_X1    g250(.A(G119), .ZN(new_n676));
  OAI221_X1 g251(.A(new_n673), .B1(new_n674), .B2(new_n675), .C1(new_n676), .C2(new_n476), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n671), .B1(new_n682), .B2(new_n670), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT35), .B(G1991), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND4_X1  g260(.A1(new_n666), .A2(new_n667), .A3(new_n669), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT36), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT31), .B(G11), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT88), .B(G28), .Z(new_n689));
  AOI21_X1  g264(.A(G29), .B1(new_n689), .B2(KEYINPUT30), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(KEYINPUT30), .B2(new_n689), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n688), .B(new_n691), .C1(new_n600), .C2(new_n670), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n660), .A2(G21), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G168), .B2(new_n660), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT87), .B(G1966), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n692), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n660), .A2(G5), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G171), .B2(new_n660), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT89), .Z(new_n700));
  INV_X1    g275(.A(G1961), .ZN(new_n701));
  OAI221_X1 g276(.A(new_n697), .B1(new_n694), .B2(new_n696), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT90), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n576), .A2(new_n660), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G4), .B2(new_n660), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT84), .B(G1348), .Z(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n595), .A2(G128), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n470), .A2(G140), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n466), .A2(G116), .ZN(new_n711));
  OAI21_X1  g286(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n709), .B(new_n710), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n670), .A2(G26), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G2067), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n707), .A2(new_n708), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n595), .A2(G129), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n466), .A2(G105), .A3(G2104), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n470), .A2(G141), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT26), .Z(new_n725));
  NAND4_X1  g300(.A1(new_n721), .A2(new_n722), .A3(new_n723), .A4(new_n725), .ZN(new_n726));
  MUX2_X1   g301(.A(G32), .B(new_n726), .S(G29), .Z(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT27), .B(G1996), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G27), .A2(G29), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G164), .B2(G29), .ZN(new_n731));
  INV_X1    g306(.A(G2078), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(G29), .A2(G35), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G162), .B2(G29), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G2090), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n729), .B(new_n733), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n670), .A2(G33), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n470), .A2(G139), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n475), .A2(G127), .ZN(new_n743));
  NAND2_X1  g318(.A1(G115), .A2(G2104), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n466), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT25), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n742), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT85), .Z(new_n749));
  OAI21_X1  g324(.A(new_n740), .B1(new_n749), .B2(new_n670), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G2072), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT24), .ZN(new_n753));
  INV_X1    g328(.A(G34), .ZN(new_n754));
  AOI21_X1  g329(.A(G29), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n753), .B2(new_n754), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G160), .B2(new_n670), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT86), .Z(new_n758));
  OAI21_X1  g333(.A(new_n751), .B1(new_n752), .B2(new_n758), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n720), .A2(new_n739), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n660), .A2(G19), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n529), .B2(new_n660), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n700), .A2(new_n701), .B1(G1341), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G2072), .B2(new_n750), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n660), .A2(G20), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT92), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT23), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n544), .B2(new_n660), .ZN(new_n768));
  INV_X1    g343(.A(G1956), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n758), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(G2084), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n737), .A2(new_n738), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n762), .B2(G1341), .ZN(new_n774));
  NOR3_X1   g349(.A1(new_n764), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n687), .A2(new_n703), .A3(new_n760), .A4(new_n775), .ZN(G150));
  INV_X1    g351(.A(G150), .ZN(G311));
  AOI22_X1  g352(.A1(G93), .A2(new_n525), .B1(new_n526), .B2(G55), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(new_n504), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT93), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G860), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT95), .B(KEYINPUT37), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n783), .A2(new_n528), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n529), .A2(new_n781), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT38), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n575), .A2(new_n583), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(KEYINPUT39), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT94), .Z(new_n795));
  INV_X1    g370(.A(G860), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n793), .B2(KEYINPUT39), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n786), .B1(new_n795), .B2(new_n797), .ZN(G145));
  XNOR2_X1  g373(.A(new_n681), .B(new_n590), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n595), .A2(G130), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n466), .A2(G118), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n803));
  AND3_X1   g378(.A1(new_n470), .A2(new_n803), .A3(G142), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n470), .B2(G142), .ZN(new_n805));
  OAI221_X1 g380(.A(new_n800), .B1(new_n801), .B2(new_n802), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n799), .B(new_n806), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n713), .B(new_n492), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(new_n726), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n809), .A2(KEYINPUT96), .A3(new_n749), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n749), .B(KEYINPUT96), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n809), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT98), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n812), .B2(new_n807), .ZN(new_n816));
  XNOR2_X1  g391(.A(G160), .B(new_n600), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G162), .ZN(new_n818));
  AOI21_X1  g393(.A(G37), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n807), .B1(KEYINPUT99), .B2(new_n812), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(KEYINPUT99), .B2(new_n812), .ZN(new_n821));
  INV_X1    g396(.A(new_n818), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n815), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT40), .Z(G395));
  NOR2_X1   g400(.A1(new_n783), .A2(G868), .ZN(new_n826));
  XNOR2_X1  g401(.A(G288), .B(G290), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  XNOR2_X1  g405(.A(G166), .B(KEYINPUT100), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n561), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n830), .A2(new_n832), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT42), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n787), .A2(new_n788), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n586), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n575), .B(new_n544), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n839), .B(KEYINPUT41), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n841), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n836), .B1(new_n844), .B2(KEYINPUT102), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(KEYINPUT102), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n845), .B(new_n846), .Z(new_n847));
  AOI21_X1  g422(.A(new_n826), .B1(new_n847), .B2(G868), .ZN(G295));
  AOI21_X1  g423(.A(new_n826), .B1(new_n847), .B2(G868), .ZN(G331));
  XNOR2_X1  g424(.A(G168), .B(G301), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n789), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n850), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n837), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n854), .A2(new_n842), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n851), .A2(KEYINPUT104), .A3(new_n853), .ZN(new_n856));
  OR3_X1    g431(.A1(new_n837), .A2(KEYINPUT104), .A3(new_n852), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n840), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR3_X1   g433(.A1(new_n855), .A2(new_n858), .A3(new_n835), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n859), .A2(G37), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n835), .B1(new_n855), .B2(new_n858), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n843), .A2(new_n857), .A3(new_n856), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n854), .A2(new_n839), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n867), .A2(new_n868), .B1(new_n834), .B2(new_n833), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n859), .A2(new_n869), .A3(G37), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n863), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n865), .A2(new_n866), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n862), .B2(new_n864), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n860), .A2(KEYINPUT105), .A3(new_n863), .A4(new_n861), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT43), .B1(new_n870), .B2(new_n876), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n874), .B(new_n875), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n872), .B1(new_n879), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g455(.A(G1384), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n492), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT45), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(KEYINPUT107), .B(G40), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n465), .A2(new_n471), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT108), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n681), .B(new_n684), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(KEYINPUT109), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(KEYINPUT109), .B2(new_n889), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n713), .B(G2067), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(G1996), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n887), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n888), .A2(new_n726), .ZN(new_n896));
  OAI221_X1 g471(.A(new_n893), .B1(new_n726), .B2(new_n895), .C1(new_n896), .C2(new_n894), .ZN(new_n897));
  NOR2_X1   g472(.A1(G290), .A2(G1986), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n887), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(KEYINPUT48), .Z(new_n900));
  NOR3_X1   g475(.A1(new_n891), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n895), .B(KEYINPUT46), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(new_n896), .A3(new_n893), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n903), .B(KEYINPUT47), .Z(new_n904));
  NAND2_X1  g479(.A1(new_n682), .A2(new_n684), .ZN(new_n905));
  OAI22_X1  g480(.A1(new_n897), .A2(new_n905), .B1(G2067), .B2(new_n713), .ZN(new_n906));
  AOI211_X1 g481(.A(new_n901), .B(new_n904), .C1(new_n888), .C2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT126), .ZN(new_n908));
  OAI21_X1  g483(.A(G8), .B1(new_n886), .B2(new_n882), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n554), .B(G1976), .C1(new_n549), .C2(new_n551), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(G1976), .B1(new_n552), .B2(new_n554), .ZN(new_n913));
  OR3_X1    g488(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT52), .ZN(new_n914));
  INV_X1    g489(.A(new_n560), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n525), .A2(G86), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n526), .A2(G48), .ZN(new_n917));
  INV_X1    g492(.A(G1981), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n915), .A2(new_n916), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(G1981), .B1(new_n558), .B2(new_n560), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT49), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(new_n909), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(KEYINPUT49), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT114), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n912), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT113), .B1(new_n912), .B2(KEYINPUT52), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n914), .B(new_n927), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT110), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n492), .A2(KEYINPUT45), .A3(new_n881), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT45), .B1(new_n492), .B2(new_n881), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n932), .A2(new_n933), .A3(new_n886), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n931), .B1(new_n934), .B2(G1971), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n882), .A2(KEYINPUT50), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n465), .A2(new_n471), .A3(new_n885), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT50), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n492), .A2(new_n938), .A3(new_n881), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT111), .B1(new_n940), .B2(G2090), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n886), .B1(KEYINPUT50), .B2(new_n882), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n942), .A2(new_n943), .A3(new_n738), .A4(new_n939), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n492), .A2(KEYINPUT45), .A3(new_n881), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n884), .A2(new_n937), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1971), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(KEYINPUT110), .A3(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n935), .A2(new_n941), .A3(new_n944), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(G303), .A2(G8), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT55), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(G8), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT112), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n949), .A2(new_n955), .A3(new_n952), .A4(G8), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n930), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n952), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT117), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT117), .ZN(new_n961));
  AOI21_X1  g536(.A(G2090), .B1(new_n940), .B2(new_n961), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n960), .A2(new_n962), .B1(new_n947), .B2(new_n946), .ZN(new_n963));
  INV_X1    g538(.A(G8), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n958), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n959), .A2(new_n752), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT118), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n946), .A2(new_n967), .A3(new_n695), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT118), .B1(new_n934), .B2(new_n696), .ZN(new_n971));
  AOI211_X1 g546(.A(new_n964), .B(G286), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n957), .A2(KEYINPUT119), .A3(new_n965), .A4(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT63), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n954), .A2(new_n956), .ZN(new_n976));
  INV_X1    g551(.A(new_n930), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n976), .A2(new_n965), .A3(new_n977), .A4(new_n972), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT119), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n972), .A2(KEYINPUT63), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n952), .B1(new_n949), .B2(G8), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n975), .A2(new_n980), .B1(new_n957), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n909), .B(KEYINPUT115), .ZN(new_n985));
  NOR2_X1   g560(.A1(G288), .A2(G1976), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT116), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n987), .A2(new_n927), .ZN(new_n988));
  INV_X1    g563(.A(new_n919), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n976), .B2(new_n930), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT120), .B1(new_n984), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n980), .A2(new_n974), .A3(new_n973), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n983), .A2(new_n957), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT120), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT56), .B(G2072), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n934), .A2(new_n998), .B1(new_n940), .B2(new_n769), .ZN(new_n999));
  NAND3_X1  g574(.A1(G299), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT57), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT121), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1001), .B1(new_n544), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n886), .A2(new_n882), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n940), .A2(new_n706), .B1(new_n718), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(new_n575), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n934), .A2(new_n998), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n959), .A2(G1956), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT61), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1012), .A2(new_n1014), .A3(new_n1004), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1014), .B1(new_n1012), .B2(new_n1004), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1006), .A2(new_n575), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT60), .B1(new_n1018), .B2(new_n1007), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT60), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n576), .A2(new_n1020), .A3(new_n1006), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(G1341), .ZN(new_n1023));
  OAI22_X1  g598(.A1(new_n946), .A2(G1996), .B1(new_n1005), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(new_n529), .A3(KEYINPUT123), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1025), .A2(KEYINPUT59), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(KEYINPUT59), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1019), .B(new_n1021), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1013), .B1(new_n1017), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n934), .A2(KEYINPUT53), .A3(new_n732), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n946), .B2(G2078), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n940), .A2(new_n701), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1030), .A2(new_n1032), .A3(G301), .A4(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT125), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n471), .A2(KEYINPUT53), .A3(G40), .A4(new_n732), .ZN(new_n1037));
  INV_X1    g612(.A(new_n462), .ZN(new_n1038));
  INV_X1    g613(.A(new_n464), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT124), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1040), .A2(new_n466), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1039), .A3(KEYINPUT124), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1037), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(new_n884), .A3(new_n945), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1032), .A2(new_n1044), .A3(new_n1033), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(G171), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1036), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT54), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1050));
  AOI21_X1  g625(.A(G301), .B1(new_n1050), .B2(new_n1030), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1045), .B2(G171), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1049), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n971), .A2(new_n966), .A3(G168), .A4(new_n968), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G8), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(KEYINPUT51), .ZN(new_n1057));
  INV_X1    g632(.A(new_n971), .ZN(new_n1058));
  OAI21_X1  g633(.A(G286), .B1(new_n969), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(G8), .A3(new_n1055), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1057), .B1(KEYINPUT51), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1029), .A2(new_n1054), .A3(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(KEYINPUT62), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT62), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1051), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1063), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n957), .A2(new_n965), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n992), .A2(new_n997), .A3(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(G290), .B(G1986), .ZN(new_n1071));
  AOI211_X1 g646(.A(new_n897), .B(new_n891), .C1(new_n887), .C2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n908), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1069), .B1(new_n995), .B2(new_n996), .ZN(new_n1074));
  AOI211_X1 g649(.A(KEYINPUT120), .B(new_n991), .C1(new_n993), .C2(new_n994), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n908), .B(new_n1072), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n907), .B1(new_n1073), .B2(new_n1077), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g653(.A(G319), .ZN(new_n1080));
  OR3_X1    g654(.A1(G401), .A2(new_n1080), .A3(G227), .ZN(new_n1081));
  NOR3_X1   g655(.A1(new_n824), .A2(G229), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g656(.A1(new_n865), .A2(new_n871), .ZN(new_n1083));
  AND2_X1   g657(.A1(new_n1082), .A2(new_n1083), .ZN(G308));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(G225));
endmodule


