//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G22gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(KEYINPUT81), .A2(G22gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(new_n204), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G141gat), .B(G148gat), .Z(new_n210));
  XNOR2_X1  g009(.A(G155gat), .B(G162gat), .ZN(new_n211));
  INV_X1    g010(.A(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G162gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT2), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n210), .A2(KEYINPUT77), .A3(new_n211), .A4(new_n214), .ZN(new_n218));
  INV_X1    g017(.A(new_n211), .ZN(new_n219));
  XOR2_X1   g018(.A(KEYINPUT76), .B(KEYINPUT2), .Z(new_n220));
  NAND2_X1  g019(.A1(new_n210), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n217), .A2(new_n218), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G197gat), .B(G204gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT71), .B(G211gat), .ZN(new_n224));
  INV_X1    g023(.A(G218gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n223), .B1(new_n226), .B2(KEYINPUT22), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n227), .A2(KEYINPUT72), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(KEYINPUT72), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G211gat), .B(G218gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT29), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n222), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G228gat), .A2(G233gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n233), .A2(new_n235), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT73), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n233), .A2(KEYINPUT73), .A3(new_n235), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n217), .A2(new_n218), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n221), .A2(new_n219), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(KEYINPUT29), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n240), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n234), .B1(new_n249), .B2(KEYINPUT3), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n241), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n239), .B1(new_n238), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n209), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n252), .A2(new_n255), .A3(new_n209), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G113gat), .B(G120gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n261));
  XNOR2_X1  g060(.A(G127gat), .B(G134gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT69), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n262), .A2(KEYINPUT68), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT1), .B1(new_n260), .B2(KEYINPUT69), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(KEYINPUT68), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n264), .B(new_n265), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n222), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT78), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n222), .A2(KEYINPUT78), .A3(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT4), .ZN(new_n274));
  INV_X1    g073(.A(new_n269), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(KEYINPUT4), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n279));
  NAND2_X1  g078(.A1(G225gat), .A2(G233gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n268), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(new_n222), .B2(new_n237), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n279), .B(new_n280), .C1(new_n250), .C2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT79), .B1(new_n278), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n276), .B1(new_n273), .B2(KEYINPUT4), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT79), .ZN(new_n286));
  INV_X1    g085(.A(new_n283), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n271), .B(new_n272), .C1(new_n222), .C2(new_n268), .ZN(new_n290));
  INV_X1    g089(.A(new_n280), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n279), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OR2_X1    g091(.A1(new_n250), .A2(new_n282), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n275), .A2(KEYINPUT4), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(new_n294), .A3(new_n280), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n273), .A2(KEYINPUT4), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n289), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G1gat), .B(G29gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT0), .ZN(new_n300));
  XNOR2_X1  g099(.A(G57gat), .B(G85gat), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n300), .B(new_n301), .Z(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n298), .A2(KEYINPUT6), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT80), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n278), .A2(KEYINPUT79), .A3(new_n283), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n286), .B1(new_n285), .B2(new_n287), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n302), .B(new_n297), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT6), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n302), .B1(new_n289), .B2(new_n297), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(new_n306), .A3(new_n310), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n305), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n241), .ZN(new_n316));
  INV_X1    g115(.A(G226gat), .ZN(new_n317));
  INV_X1    g116(.A(G233gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n321));
  INV_X1    g120(.A(G183gat), .ZN(new_n322));
  INV_X1    g121(.A(G190gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT65), .ZN(new_n327));
  NOR2_X1   g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT23), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n330), .B1(G169gat), .B2(G176gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n331), .B2(new_n328), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT66), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n326), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT25), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n337), .A2(new_n338), .A3(new_n332), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT27), .B(G183gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n323), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT28), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  NOR3_X1   g144(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n346), .B1(G169gat), .B2(G176gat), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n347), .A2(new_n348), .B1(G183gat), .B2(G190gat), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n345), .A2(KEYINPUT67), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT67), .B1(new_n345), .B2(new_n349), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n341), .A2(KEYINPUT74), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n345), .A2(new_n349), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT67), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n345), .A2(KEYINPUT67), .A3(new_n349), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n339), .B1(new_n334), .B2(new_n335), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n354), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n320), .B1(new_n353), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n360), .B1(new_n345), .B2(new_n349), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n319), .A2(KEYINPUT29), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n316), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n353), .A2(new_n361), .A3(new_n364), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n363), .A2(new_n319), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n245), .A3(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G8gat), .B(G36gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(G64gat), .B(G92gat), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n371), .B(new_n372), .Z(new_n373));
  NAND3_X1  g172(.A1(new_n367), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n374), .A2(KEYINPUT30), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT30), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n367), .A2(new_n376), .A3(new_n370), .A4(new_n373), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT75), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n367), .A2(new_n370), .ZN(new_n380));
  INV_X1    g179(.A(new_n373), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AOI211_X1 g181(.A(KEYINPUT75), .B(new_n373), .C1(new_n367), .C2(new_n370), .ZN(new_n383));
  OAI22_X1  g182(.A1(new_n375), .A2(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n259), .B1(new_n315), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G15gat), .B(G43gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(G71gat), .B(G99gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n341), .A2(new_n281), .A3(new_n352), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n268), .B1(new_n359), .B2(new_n360), .ZN(new_n390));
  INV_X1    g189(.A(G227gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(new_n318), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n388), .B1(new_n393), .B2(KEYINPUT32), .ZN(new_n394));
  INV_X1    g193(.A(new_n393), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n394), .B1(KEYINPUT33), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n388), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n397), .A2(KEYINPUT70), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(KEYINPUT70), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(KEYINPUT33), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n393), .A2(KEYINPUT32), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT34), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n389), .A2(new_n390), .ZN(new_n404));
  INV_X1    g203(.A(new_n392), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI211_X1 g205(.A(KEYINPUT34), .B(new_n392), .C1(new_n389), .C2(new_n390), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n402), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n396), .A2(new_n401), .A3(new_n408), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n410), .A2(KEYINPUT36), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT36), .B1(new_n410), .B2(new_n411), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n384), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n374), .A2(KEYINPUT30), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n377), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n419), .B(KEYINPUT82), .C1(new_n382), .C2(new_n383), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT83), .B(KEYINPUT40), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n274), .A2(new_n293), .A3(new_n277), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n291), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n290), .A2(new_n291), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT39), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n303), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n422), .A2(new_n425), .A3(new_n291), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n421), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n423), .A2(new_n426), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n430), .A2(KEYINPUT40), .A3(new_n302), .A4(new_n428), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT84), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n427), .A2(KEYINPUT84), .A3(KEYINPUT40), .A4(new_n428), .ZN(new_n434));
  AOI211_X1 g233(.A(new_n312), .B(new_n429), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n417), .A2(new_n420), .A3(new_n435), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n252), .A2(new_n255), .A3(new_n209), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n437), .A2(new_n256), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n380), .A2(new_n381), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT37), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n373), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n439), .A2(new_n442), .B1(KEYINPUT37), .B2(new_n380), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT38), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n245), .B1(new_n368), .B2(new_n369), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n353), .A2(new_n361), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n319), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n363), .A2(new_n365), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n241), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT85), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n445), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n447), .A2(KEYINPUT85), .A3(new_n241), .A4(new_n448), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n440), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n373), .B1(new_n367), .B2(new_n370), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n444), .B1(new_n454), .B2(new_n441), .ZN(new_n455));
  OAI22_X1  g254(.A1(new_n443), .A2(new_n444), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n309), .A2(new_n310), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n304), .B(new_n374), .C1(new_n457), .C2(new_n312), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n438), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n385), .B(new_n415), .C1(new_n436), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n417), .A2(new_n420), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n457), .A2(new_n312), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(new_n305), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT35), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n438), .A2(new_n410), .A3(new_n464), .A4(new_n411), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n438), .A2(new_n410), .A3(new_n411), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n315), .A2(new_n384), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n469), .B2(new_n464), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n460), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(G229gat), .A2(G233gat), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(G29gat), .A2(G36gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT14), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(G29gat), .A2(G36gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(KEYINPUT87), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT15), .ZN(new_n480));
  INV_X1    g279(.A(G43gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G50gat), .ZN(new_n482));
  INV_X1    g281(.A(G50gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G43gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n480), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n484), .A3(KEYINPUT86), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT88), .B(G43gat), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n482), .B1(new_n490), .B2(G50gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n480), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n479), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT89), .ZN(new_n494));
  INV_X1    g293(.A(new_n479), .ZN(new_n495));
  INV_X1    g294(.A(new_n489), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n493), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n479), .A2(new_n489), .A3(new_n492), .A4(KEYINPUT89), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G15gat), .B(G22gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT16), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n500), .B1(new_n501), .B2(G1gat), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(G1gat), .B2(new_n500), .ZN(new_n503));
  XOR2_X1   g302(.A(new_n503), .B(G8gat), .Z(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT90), .B1(new_n499), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT90), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n497), .A2(new_n510), .A3(KEYINPUT17), .A4(new_n498), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT17), .B1(new_n497), .B2(new_n498), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(new_n505), .ZN(new_n514));
  AOI211_X1 g313(.A(new_n473), .B(new_n507), .C1(new_n512), .C2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT91), .B1(new_n515), .B2(KEYINPUT18), .ZN(new_n516));
  XNOR2_X1  g315(.A(G113gat), .B(G141gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(G197gat), .ZN(new_n518));
  XOR2_X1   g317(.A(KEYINPUT11), .B(G169gat), .Z(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n520), .B(KEYINPUT12), .Z(new_n521));
  XNOR2_X1  g320(.A(new_n499), .B(new_n505), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n472), .B(KEYINPUT13), .Z(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(new_n515), .B2(KEYINPUT18), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n512), .A2(new_n514), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(new_n472), .A3(new_n506), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT18), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n516), .B(new_n521), .C1(new_n525), .C2(new_n529), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n527), .A2(new_n528), .B1(new_n522), .B2(new_n523), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n515), .A2(KEYINPUT18), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT91), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(new_n527), .B2(new_n528), .ZN(new_n534));
  INV_X1    g333(.A(new_n521), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n531), .B(new_n532), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(G85gat), .ZN(new_n539));
  INV_X1    g338(.A(G92gat), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT7), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT7), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(G85gat), .A3(G92gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(new_n540), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G99gat), .ZN(new_n548));
  INV_X1    g347(.A(G106gat), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT8), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n544), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G99gat), .B(G106gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n544), .A2(new_n552), .A3(new_n547), .A4(new_n550), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT99), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n513), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n512), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n554), .A2(new_n555), .ZN(new_n562));
  AND2_X1   g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n499), .A2(new_n562), .B1(KEYINPUT41), .B2(new_n563), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n559), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n561), .B1(new_n559), .B2(new_n564), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT97), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n563), .A2(KEYINPUT41), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n569), .B(new_n570), .Z(new_n571));
  OAI211_X1 g370(.A(new_n567), .B(new_n571), .C1(KEYINPUT100), .C2(new_n566), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n571), .B1(new_n566), .B2(KEYINPUT100), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(new_n566), .B2(new_n565), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT92), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(KEYINPUT92), .A2(G71gat), .A3(G78gat), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n578), .B(new_n579), .C1(G71gat), .C2(G78gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT9), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G57gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(G64gat), .ZN(new_n584));
  INV_X1    g383(.A(G64gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(G57gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT93), .A2(new_n582), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT93), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n576), .A2(new_n588), .A3(new_n581), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n580), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G71gat), .B(G78gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n582), .A2(KEYINPUT93), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n584), .A2(new_n586), .ZN(new_n593));
  AND4_X1   g392(.A1(new_n591), .A2(new_n592), .A3(new_n589), .A4(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT94), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT94), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n592), .A2(new_n593), .A3(new_n591), .A4(new_n589), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n592), .A2(new_n589), .A3(new_n593), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n596), .B(new_n597), .C1(new_n598), .C2(new_n580), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT21), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n504), .B1(new_n600), .B2(new_n601), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G127gat), .B(G155gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT96), .ZN(new_n609));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT95), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n609), .B(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G183gat), .B(G211gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n604), .A2(new_n605), .ZN(new_n616));
  OR3_X1    g415(.A1(new_n607), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(new_n607), .B2(new_n616), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT101), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n595), .A2(new_n556), .A3(new_n599), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n554), .B(new_n555), .C1(new_n590), .C2(new_n594), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT10), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n562), .A2(new_n595), .A3(KEYINPUT10), .A4(new_n599), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n623), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(new_n622), .A3(new_n625), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT102), .ZN(new_n633));
  XNOR2_X1  g432(.A(G176gat), .B(G204gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(new_n635), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR4_X1   g438(.A1(new_n538), .A2(new_n575), .A3(new_n620), .A4(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n471), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n315), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G1gat), .ZN(G1324gat));
  INV_X1    g442(.A(new_n641), .ZN(new_n644));
  OAI21_X1  g443(.A(G8gat), .B1(new_n644), .B2(new_n461), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT42), .ZN(new_n646));
  INV_X1    g445(.A(new_n461), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT16), .B(G8gat), .Z(new_n648));
  NAND3_X1  g447(.A1(new_n641), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n646), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n650), .A2(KEYINPUT103), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(KEYINPUT103), .ZN(new_n652));
  OAI221_X1 g451(.A(new_n645), .B1(new_n646), .B2(new_n649), .C1(new_n651), .C2(new_n652), .ZN(G1325gat));
  NAND2_X1  g452(.A1(new_n410), .A2(new_n411), .ZN(new_n654));
  OR3_X1    g453(.A1(new_n644), .A2(G15gat), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(G15gat), .B1(new_n644), .B2(new_n415), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(G1326gat));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n259), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT104), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT43), .B(G22gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  NAND2_X1  g460(.A1(new_n451), .A2(new_n452), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT37), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT38), .B1(new_n439), .B2(new_n442), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n380), .A2(KEYINPUT37), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(new_n454), .B2(new_n441), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n663), .A2(new_n664), .B1(new_n666), .B2(KEYINPUT38), .ZN(new_n667));
  INV_X1    g466(.A(new_n458), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n259), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n417), .A2(new_n435), .A3(new_n420), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n414), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n654), .A2(new_n259), .ZN(new_n672));
  INV_X1    g471(.A(new_n384), .ZN(new_n673));
  INV_X1    g472(.A(new_n314), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n674), .A2(new_n311), .A3(new_n312), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n672), .B(new_n673), .C1(new_n675), .C2(new_n305), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT35), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n671), .A2(new_n385), .B1(new_n677), .B2(new_n467), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n572), .A2(new_n574), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n538), .A2(new_n619), .A3(new_n639), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n315), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n682), .A2(G29gat), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT45), .Z(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n678), .B2(new_n679), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n471), .A2(KEYINPUT44), .A3(new_n575), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(new_n315), .A3(new_n681), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G29gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n685), .A2(new_n691), .ZN(G1328gat));
  NOR2_X1   g491(.A1(new_n461), .A2(G36gat), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n680), .A2(new_n681), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT46), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n687), .A2(new_n688), .A3(new_n647), .A4(new_n681), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G36gat), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OR3_X1    g497(.A1(new_n695), .A2(new_n698), .A3(KEYINPUT105), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT105), .B1(new_n695), .B2(new_n698), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1329gat));
  NAND4_X1  g500(.A1(new_n687), .A2(new_n688), .A3(new_n414), .A4(new_n681), .ZN(new_n702));
  INV_X1    g501(.A(new_n490), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n654), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n680), .A2(new_n705), .A3(new_n490), .A4(new_n681), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT106), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1330gat));
  NAND4_X1  g508(.A1(new_n689), .A2(G50gat), .A3(new_n259), .A4(new_n681), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n483), .B1(new_n682), .B2(new_n438), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1331gat));
  NOR2_X1   g513(.A1(new_n575), .A2(new_n620), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n538), .A3(new_n639), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n678), .A2(KEYINPUT108), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT108), .B1(new_n678), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n683), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(new_n583), .ZN(G1332gat));
  INV_X1    g520(.A(new_n719), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n647), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT49), .B(G64gat), .Z(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n723), .B2(new_n725), .ZN(G1333gat));
  INV_X1    g525(.A(G71gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n722), .A2(new_n727), .A3(new_n705), .ZN(new_n728));
  OAI21_X1  g527(.A(G71gat), .B1(new_n719), .B2(new_n415), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n728), .A2(KEYINPUT50), .A3(new_n729), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1334gat));
  NAND2_X1  g533(.A1(new_n722), .A2(new_n259), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g535(.A1(new_n545), .A2(new_n546), .ZN(new_n737));
  INV_X1    g536(.A(new_n639), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n537), .A2(new_n619), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n689), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n737), .B1(new_n740), .B2(new_n683), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n678), .B2(new_n679), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n471), .A2(KEYINPUT109), .A3(new_n575), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n537), .A2(new_n619), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT51), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  INV_X1    g547(.A(new_n746), .ZN(new_n749));
  AOI211_X1 g548(.A(new_n748), .B(new_n749), .C1(new_n743), .C2(new_n744), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n315), .A2(new_n545), .A3(new_n546), .A4(new_n639), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n741), .B1(new_n751), .B2(new_n752), .ZN(G1336gat));
  NAND3_X1  g552(.A1(new_n647), .A2(new_n540), .A3(new_n639), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT110), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT109), .B1(new_n471), .B2(new_n575), .ZN(new_n756));
  AOI211_X1 g555(.A(new_n742), .B(new_n679), .C1(new_n460), .C2(new_n470), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n746), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n748), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n745), .A2(KEYINPUT51), .A3(new_n746), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n755), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n687), .A2(new_n688), .A3(new_n647), .A4(new_n739), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G92gat), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT52), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n766), .B(new_n763), .C1(new_n751), .C2(new_n755), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1337gat));
  OAI21_X1  g567(.A(G99gat), .B1(new_n740), .B2(new_n415), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n705), .A2(new_n548), .A3(new_n639), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT111), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n751), .B2(new_n771), .ZN(G1338gat));
  NOR3_X1   g571(.A1(new_n438), .A2(G106gat), .A3(new_n738), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n747), .B2(new_n750), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n687), .A2(new_n688), .A3(new_n259), .A4(new_n739), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G106gat), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n774), .B(new_n776), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n776), .B2(new_n777), .ZN(new_n780));
  INV_X1    g579(.A(new_n773), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n759), .B2(new_n760), .ZN(new_n782));
  INV_X1    g581(.A(new_n776), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n779), .A2(new_n784), .ZN(G1339gat));
  NAND2_X1  g584(.A1(KEYINPUT115), .A2(G113gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(KEYINPUT115), .B(G113gat), .ZN(new_n787));
  NOR4_X1   g586(.A1(new_n575), .A2(new_n537), .A3(new_n620), .A4(new_n639), .ZN(new_n788));
  INV_X1    g587(.A(new_n626), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(new_n622), .A3(new_n627), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n790), .A2(KEYINPUT54), .A3(new_n629), .ZN(new_n791));
  XNOR2_X1  g590(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n623), .B(new_n792), .C1(new_n626), .C2(new_n628), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n793), .A2(new_n794), .A3(new_n635), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n794), .B1(new_n793), .B2(new_n635), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n791), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n637), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n798), .B2(new_n797), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n527), .A2(new_n528), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n532), .A2(new_n801), .A3(new_n535), .A4(new_n524), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n507), .B1(new_n512), .B2(new_n514), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n803), .A2(new_n472), .B1(new_n522), .B2(new_n523), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n520), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n575), .A2(new_n800), .A3(new_n806), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n537), .A2(new_n800), .B1(new_n806), .B2(new_n639), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n808), .B2(new_n575), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n788), .B1(new_n809), .B2(new_n620), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(new_n468), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n647), .A2(new_n683), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n537), .ZN(new_n814));
  MUX2_X1   g613(.A(new_n786), .B(new_n787), .S(new_n814), .Z(G1340gat));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n639), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g616(.A1(new_n813), .A2(new_n619), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g618(.A1(new_n813), .A2(new_n575), .ZN(new_n820));
  OR3_X1    g619(.A1(new_n820), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT56), .B1(new_n820), .B2(G134gat), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(G134gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(G1343gat));
  INV_X1    g623(.A(new_n788), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n790), .A2(KEYINPUT54), .A3(new_n629), .ZN(new_n826));
  INV_X1    g625(.A(new_n796), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n793), .A2(new_n794), .A3(new_n635), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n636), .B1(new_n829), .B2(KEYINPUT55), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(KEYINPUT55), .B2(new_n829), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n802), .A2(new_n805), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n679), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n806), .A2(new_n639), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n538), .B2(new_n831), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n833), .B1(new_n835), .B2(new_n679), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n825), .B1(new_n836), .B2(new_n619), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n259), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n812), .A2(new_n415), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n537), .ZN(new_n841));
  INV_X1    g640(.A(G141gat), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n839), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n845), .B1(new_n810), .B2(new_n438), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n438), .A2(new_n845), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n797), .A2(KEYINPUT116), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n850), .B(new_n791), .C1(new_n795), .C2(new_n796), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n798), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n830), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT117), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(new_n830), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n537), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n575), .B1(new_n857), .B2(new_n834), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n620), .B1(new_n858), .B2(new_n833), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n848), .B1(new_n859), .B2(new_n825), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n846), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI211_X1 g661(.A(KEYINPUT118), .B(new_n848), .C1(new_n859), .C2(new_n825), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n844), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n538), .A2(new_n842), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n843), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT119), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT58), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n867), .A2(KEYINPUT119), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1344gat));
  NAND2_X1  g671(.A1(new_n838), .A2(KEYINPUT57), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n859), .A2(new_n825), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n845), .A3(new_n259), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n873), .A2(new_n875), .A3(new_n639), .A4(new_n844), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G148gat), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT59), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n639), .B(new_n844), .C1(new_n862), .C2(new_n863), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880));
  INV_X1    g679(.A(G148gat), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(KEYINPUT59), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n880), .B1(new_n879), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n878), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n840), .A2(new_n881), .A3(new_n639), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1345gat));
  OAI21_X1  g686(.A(G155gat), .B1(new_n864), .B2(new_n620), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n840), .A2(new_n212), .A3(new_n619), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1346gat));
  OAI21_X1  g689(.A(G162gat), .B1(new_n864), .B2(new_n679), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n840), .A2(new_n213), .A3(new_n575), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1347gat));
  NOR4_X1   g692(.A1(new_n810), .A2(new_n315), .A3(new_n468), .A4(new_n461), .ZN(new_n894));
  AOI21_X1  g693(.A(G169gat), .B1(new_n894), .B2(new_n537), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n461), .A2(new_n315), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n811), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT121), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n811), .A2(new_n899), .A3(new_n896), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n537), .A2(G169gat), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n895), .B1(new_n901), .B2(new_n902), .ZN(G1348gat));
  AOI21_X1  g702(.A(G176gat), .B1(new_n894), .B2(new_n639), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n904), .A2(KEYINPUT122), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(KEYINPUT122), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n639), .A2(G176gat), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n905), .A2(new_n906), .B1(new_n901), .B2(new_n907), .ZN(G1349gat));
  AND3_X1   g707(.A1(new_n894), .A2(new_n342), .A3(new_n619), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n898), .A2(new_n619), .A3(new_n900), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(G183gat), .ZN(new_n911));
  NAND2_X1  g710(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n911), .B(new_n912), .ZN(G1350gat));
  AOI21_X1  g712(.A(new_n323), .B1(new_n901), .B2(new_n575), .ZN(new_n914));
  XOR2_X1   g713(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n894), .A2(new_n323), .A3(new_n575), .ZN(new_n917));
  OR2_X1    g716(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n916), .B(new_n917), .C1(new_n914), .C2(new_n918), .ZN(G1351gat));
  NOR3_X1   g718(.A1(new_n461), .A2(new_n414), .A3(new_n438), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT125), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n810), .A2(new_n315), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  XOR2_X1   g723(.A(KEYINPUT126), .B(G197gat), .Z(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(new_n537), .A3(new_n925), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n873), .A2(new_n875), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n461), .A2(new_n414), .A3(new_n315), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n538), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n926), .B1(new_n930), .B2(new_n925), .ZN(G1352gat));
  NOR3_X1   g730(.A1(new_n923), .A2(G204gat), .A3(new_n738), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT62), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n927), .A2(new_n639), .A3(new_n928), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G204gat), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1353gat));
  NAND3_X1  g735(.A1(new_n924), .A2(new_n224), .A3(new_n619), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n927), .A2(new_n619), .A3(new_n928), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n938), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT63), .B1(new_n938), .B2(G211gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(G1354gat));
  OAI21_X1  g740(.A(G218gat), .B1(new_n929), .B2(new_n679), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n225), .A3(new_n575), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1355gat));
endmodule


