//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT15), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT83), .B(G36gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G29gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT84), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT84), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n213), .A3(G29gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(G29gat), .A2(G36gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT14), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT85), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n218), .B(new_n219), .C1(KEYINPUT15), .C2(new_n207), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n209), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n207), .B2(KEYINPUT15), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n216), .B(KEYINPUT14), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n224), .A2(new_n208), .A3(new_n214), .A4(new_n212), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(G1gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(G1gat), .B2(new_n227), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(G8gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT86), .B1(new_n226), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT86), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n221), .A2(new_n236), .A3(KEYINPUT17), .A4(new_n225), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n231), .B1(new_n226), .B2(new_n234), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n233), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT87), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(KEYINPUT18), .A3(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n226), .A2(new_n231), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n233), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n242), .B(KEYINPUT13), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT18), .B1(new_n240), .B2(new_n242), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n206), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n240), .A2(new_n242), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT18), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n206), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n253), .A2(new_n254), .A3(new_n243), .A4(new_n247), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(G15gat), .B(G43gat), .Z(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT69), .ZN(new_n259));
  XNOR2_X1  g058(.A(G71gat), .B(G99gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G227gat), .A2(G233gat), .ZN(new_n262));
  XOR2_X1   g061(.A(G127gat), .B(G134gat), .Z(new_n263));
  XNOR2_X1  g062(.A(G113gat), .B(G120gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(G113gat), .B(G120gat), .Z(new_n268));
  XNOR2_X1  g067(.A(G127gat), .B(G134gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n269), .A3(new_n265), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT25), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT23), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT23), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n280), .B1(G169gat), .B2(G176gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n278), .A2(new_n279), .A3(new_n281), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n276), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n278), .A2(new_n282), .A3(new_n281), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n285), .A2(KEYINPUT64), .ZN(new_n286));
  INV_X1    g085(.A(G183gat), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT27), .B1(new_n287), .B2(KEYINPUT66), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT66), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT27), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n290), .A3(G183gat), .ZN(new_n291));
  INV_X1    g090(.A(G190gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n288), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT27), .B(G183gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(G190gat), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n293), .A2(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n277), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT26), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n282), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n277), .A2(KEYINPUT26), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n273), .A3(new_n301), .ZN(new_n302));
  OAI22_X1  g101(.A1(new_n284), .A2(new_n286), .B1(new_n297), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT25), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT65), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n280), .A2(G169gat), .A3(G176gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n282), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n278), .A2(KEYINPUT65), .A3(new_n282), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n274), .A2(new_n275), .B1(new_n298), .B2(new_n280), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n304), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n271), .B1(new_n303), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n311), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT25), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n267), .A2(new_n270), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n293), .A2(new_n294), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n295), .A2(new_n296), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n302), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n285), .A2(KEYINPUT64), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(new_n283), .A3(new_n276), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n315), .A2(new_n316), .A3(new_n321), .A4(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n262), .B1(new_n313), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT68), .B(KEYINPUT33), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(KEYINPUT32), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n261), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT70), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g129(.A(KEYINPUT70), .B(new_n261), .C1(new_n325), .C2(new_n327), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n324), .A3(new_n262), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT34), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT34), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n313), .A2(new_n324), .A3(new_n336), .A4(new_n262), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n334), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n337), .A2(new_n335), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n326), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n261), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT32), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(new_n325), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n332), .A2(new_n340), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT72), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n344), .B1(new_n330), .B2(new_n331), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n349), .A2(KEYINPUT72), .A3(new_n340), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n332), .A2(new_n345), .ZN(new_n352));
  INV_X1    g151(.A(new_n340), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(KEYINPUT73), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT73), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n355), .B1(new_n349), .B2(new_n340), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT31), .B(G50gat), .ZN(new_n359));
  INV_X1    g158(.A(G106gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(G141gat), .B(G148gat), .Z(new_n363));
  INV_X1    g162(.A(G155gat), .ZN(new_n364));
  INV_X1    g163(.A(G162gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(KEYINPUT2), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n363), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G141gat), .B(G148gat), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n367), .B(new_n366), .C1(new_n371), .C2(KEYINPUT2), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G197gat), .B(G204gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT22), .ZN(new_n378));
  INV_X1    g177(.A(G211gat), .ZN(new_n379));
  INV_X1    g178(.A(G218gat), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G211gat), .B(G218gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n377), .A3(new_n381), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n376), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n370), .A2(new_n372), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT29), .B1(new_n385), .B2(new_n386), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n390), .B1(new_n391), .B2(KEYINPUT3), .ZN(new_n392));
  NAND2_X1  g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n389), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT79), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n389), .A2(new_n392), .A3(new_n397), .A4(new_n394), .ZN(new_n398));
  INV_X1    g197(.A(new_n373), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n390), .B1(new_n391), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n389), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n393), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n396), .A2(new_n398), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(G22gat), .ZN(new_n404));
  INV_X1    g203(.A(G78gat), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n395), .A2(KEYINPUT79), .B1(new_n401), .B2(new_n393), .ZN(new_n406));
  INV_X1    g205(.A(G22gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n407), .A3(new_n398), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n405), .B1(new_n404), .B2(new_n408), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n362), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n407), .B1(new_n406), .B2(new_n398), .ZN(new_n413));
  AND4_X1   g212(.A1(new_n407), .A2(new_n396), .A3(new_n398), .A4(new_n402), .ZN(new_n414));
  OAI21_X1  g213(.A(G78gat), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(new_n409), .A3(new_n361), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n358), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n390), .A2(KEYINPUT3), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(new_n374), .A3(new_n271), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n316), .A2(KEYINPUT4), .A3(new_n372), .A4(new_n370), .ZN(new_n421));
  NAND2_X1  g220(.A1(G225gat), .A2(G233gat), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n370), .A2(new_n267), .A3(new_n270), .A4(new_n372), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n420), .A2(new_n421), .A3(new_n422), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(KEYINPUT77), .A2(KEYINPUT5), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n428), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(G1gat), .B(G29gat), .Z(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT0), .ZN(new_n433));
  XNOR2_X1  g232(.A(G57gat), .B(G85gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n271), .A2(new_n390), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n437), .A2(new_n423), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT5), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n438), .A2(new_n439), .A3(new_n422), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(KEYINPUT78), .B(KEYINPUT6), .Z(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n431), .A2(new_n436), .A3(new_n441), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT81), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n440), .B1(new_n429), .B2(new_n430), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT81), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n446), .A2(new_n447), .A3(new_n436), .A4(new_n443), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n441), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n435), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n443), .B1(new_n446), .B2(new_n436), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n445), .A2(new_n448), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(G226gat), .A2(G233gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n375), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(new_n303), .B2(new_n312), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n315), .A2(new_n323), .A3(new_n321), .A4(new_n453), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n387), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n387), .B1(new_n455), .B2(new_n456), .ZN(new_n459));
  XNOR2_X1  g258(.A(G8gat), .B(G36gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(G64gat), .B(G92gat), .ZN(new_n461));
  XOR2_X1   g260(.A(new_n460), .B(new_n461), .Z(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n458), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(KEYINPUT74), .A3(KEYINPUT30), .ZN(new_n465));
  INV_X1    g264(.A(new_n459), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n466), .A2(new_n457), .A3(KEYINPUT30), .A4(new_n462), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT74), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n462), .B1(new_n466), .B2(new_n457), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n458), .A2(new_n459), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n462), .ZN(new_n473));
  XOR2_X1   g272(.A(KEYINPUT75), .B(KEYINPUT30), .Z(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n471), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT82), .B(KEYINPUT35), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n452), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n418), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n416), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n361), .B1(new_n415), .B2(new_n409), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n444), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(new_n450), .B2(new_n451), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n485), .A2(new_n477), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n349), .A2(new_n340), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n483), .A2(new_n486), .A3(new_n351), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT35), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n480), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n430), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n426), .A2(new_n428), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n436), .B(new_n441), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n442), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n446), .A2(new_n436), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n444), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n463), .B1(new_n458), .B2(new_n459), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(new_n464), .B2(new_n474), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(new_n469), .B2(new_n465), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n416), .A2(new_n412), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT40), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n420), .A2(new_n425), .A3(new_n421), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT39), .ZN(new_n504));
  INV_X1    g303(.A(new_n422), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n435), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n437), .A2(new_n422), .A3(new_n423), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT39), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n503), .B2(new_n505), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n502), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n503), .A2(new_n505), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n512), .A2(KEYINPUT39), .A3(new_n508), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n513), .A2(KEYINPUT40), .A3(new_n435), .A4(new_n506), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n514), .A3(new_n494), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n515), .B1(new_n470), .B2(new_n476), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n481), .A2(new_n516), .A3(new_n482), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT37), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n462), .B1(new_n472), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(new_n518), .B2(new_n472), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT38), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT80), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n472), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n518), .B1(new_n458), .B2(KEYINPUT80), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT38), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n464), .B1(new_n525), .B2(new_n519), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n452), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n501), .B1(new_n517), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n351), .A2(KEYINPUT36), .A3(new_n488), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n348), .A2(new_n350), .B1(new_n354), .B2(new_n356), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(KEYINPUT36), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n257), .B1(new_n491), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G85gat), .A2(G92gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT7), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(G85gat), .A3(G92gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT92), .ZN(new_n539));
  INV_X1    g338(.A(G85gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G92gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(KEYINPUT92), .A2(G85gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G99gat), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT8), .B1(new_n545), .B2(new_n360), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n538), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G99gat), .B(G106gat), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n538), .A2(new_n544), .A3(new_n548), .A4(new_n546), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n552), .B1(new_n226), .B2(new_n234), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n238), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n226), .A2(new_n552), .ZN(new_n555));
  AND2_X1   g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT41), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(KEYINPUT94), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT94), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n558), .B1(new_n238), .B2(new_n553), .ZN(new_n564));
  INV_X1    g363(.A(new_n561), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G134gat), .B(G162gat), .Z(new_n567));
  NOR2_X1   g366(.A1(new_n556), .A2(KEYINPUT41), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(new_n564), .B2(new_n565), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n562), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT95), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n562), .A2(new_n566), .A3(new_n570), .A4(KEYINPUT95), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT93), .B1(new_n560), .B2(new_n561), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n576), .B1(new_n561), .B2(new_n560), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n564), .A2(KEYINPUT93), .A3(new_n565), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n569), .B(KEYINPUT91), .Z(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(G57gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(G64gat), .ZN(new_n583));
  INV_X1    g382(.A(G64gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(G57gat), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT88), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n583), .A2(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT88), .B1(new_n590), .B2(KEYINPUT9), .ZN(new_n591));
  NOR2_X1   g390(.A1(G71gat), .A2(G78gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT89), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n589), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT89), .B1(new_n590), .B2(new_n592), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n588), .A2(new_n591), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n590), .A2(new_n592), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT9), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n589), .A2(new_n587), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n584), .A2(G57gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n582), .A2(G64gat), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n586), .A2(new_n587), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n598), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n597), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G127gat), .B(G155gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  AND2_X1   g409(.A1(new_n597), .A2(new_n605), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n231), .B1(KEYINPUT21), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n610), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT90), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G183gat), .B(G211gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n613), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n581), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G120gat), .B(G148gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(G176gat), .B(G204gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  INV_X1    g426(.A(KEYINPUT96), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n551), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n629), .A2(new_n605), .A3(new_n597), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n552), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n550), .A2(new_n551), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n632), .A2(new_n605), .A3(new_n597), .A4(new_n629), .ZN(new_n633));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n631), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n627), .B1(new_n636), .B2(KEYINPUT98), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n637), .B1(KEYINPUT98), .B2(new_n636), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n552), .A2(new_n630), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n632), .B1(new_n611), .B2(new_n629), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n632), .A2(new_n606), .A3(new_n639), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(KEYINPUT97), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT97), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT10), .B1(new_n631), .B2(new_n633), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n646), .B1(new_n647), .B2(new_n643), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n645), .A2(new_n648), .A3(new_n634), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n638), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n647), .A2(new_n643), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n636), .B1(new_n651), .B2(new_n635), .ZN(new_n652));
  INV_X1    g451(.A(new_n627), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n624), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n533), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n485), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT99), .B(G1gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(G1324gat));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n477), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT16), .B(G8gat), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT100), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n665), .A2(KEYINPUT42), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(KEYINPUT42), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(G8gat), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(G1325gat));
  INV_X1    g468(.A(new_n659), .ZN(new_n670));
  OAI21_X1  g469(.A(G15gat), .B1(new_n670), .B2(new_n531), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n358), .A2(G15gat), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(new_n670), .B2(new_n672), .ZN(G1326gat));
  NAND2_X1  g472(.A1(new_n659), .A2(new_n417), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT43), .B(G22gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  INV_X1    g475(.A(new_n581), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n677), .A2(new_n622), .A3(new_n655), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n533), .A2(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n679), .A2(G29gat), .A3(new_n497), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT45), .Z(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n418), .A2(new_n479), .B1(new_n489), .B2(KEYINPUT35), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT36), .B1(new_n351), .B2(new_n357), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT36), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n685), .B(new_n487), .C1(new_n348), .C2(new_n350), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n417), .B1(new_n485), .B2(new_n477), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n452), .A2(new_n521), .A3(new_n526), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n412), .B(new_n416), .C1(new_n500), .C2(new_n515), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT102), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT102), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n528), .A2(new_n531), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n683), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n682), .B1(new_n695), .B2(new_n677), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n491), .A2(new_n532), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(KEYINPUT44), .A3(new_n581), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n622), .B(KEYINPUT101), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n701), .A2(new_n257), .A3(new_n655), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G29gat), .B1(new_n703), .B2(new_n497), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n681), .A2(new_n704), .ZN(G1328gat));
  OAI21_X1  g504(.A(new_n210), .B1(new_n703), .B2(new_n500), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n679), .A2(new_n500), .A3(new_n210), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT46), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1329gat));
  NAND4_X1  g508(.A1(new_n696), .A2(new_n687), .A3(new_n698), .A4(new_n702), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G43gat), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT47), .B1(new_n711), .B2(KEYINPUT103), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n358), .A2(G43gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n679), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n712), .B(new_n714), .ZN(G1330gat));
  NAND3_X1  g514(.A1(new_n533), .A2(new_n417), .A3(new_n678), .ZN(new_n716));
  INV_X1    g515(.A(G50gat), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n716), .A2(new_n717), .B1(KEYINPUT104), .B2(KEYINPUT48), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n417), .A2(G50gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n703), .B2(new_n719), .ZN(new_n720));
  OR2_X1    g519(.A1(KEYINPUT104), .A2(KEYINPUT48), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1331gat));
  NAND3_X1  g521(.A1(new_n624), .A2(new_n257), .A3(new_n655), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n695), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n485), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G57gat), .ZN(G1332gat));
  INV_X1    g525(.A(new_n724), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n500), .ZN(new_n728));
  NOR2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  AND2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n728), .B2(new_n729), .ZN(G1333gat));
  NAND3_X1  g531(.A1(new_n724), .A2(G71gat), .A3(new_n687), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n727), .A2(new_n358), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n734), .B2(G71gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g535(.A1(new_n724), .A2(new_n417), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT105), .B(G78gat), .Z(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1335gat));
  NAND2_X1  g538(.A1(new_n541), .A2(new_n543), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n256), .A2(new_n622), .A3(new_n656), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n699), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n742), .B2(new_n497), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n528), .A2(new_n531), .A3(new_n693), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n693), .B1(new_n528), .B2(new_n531), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n491), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n256), .A2(new_n622), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n746), .A2(new_n581), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n748), .A2(new_n749), .A3(KEYINPUT51), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(KEYINPUT51), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT106), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n748), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n497), .A2(new_n656), .A3(new_n740), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT107), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n750), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n743), .A2(new_n757), .ZN(G1336gat));
  NAND4_X1  g557(.A1(new_n696), .A2(new_n477), .A3(new_n698), .A4(new_n741), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n759), .A2(G92gat), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(KEYINPUT52), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n500), .A2(new_n656), .A3(G92gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n750), .A2(new_n754), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n752), .A2(KEYINPUT108), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n748), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n746), .A2(new_n581), .A3(new_n747), .A4(new_n766), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n765), .B1(new_n770), .B2(new_n762), .ZN(new_n771));
  INV_X1    g570(.A(new_n762), .ZN(new_n772));
  AOI211_X1 g571(.A(KEYINPUT109), .B(new_n772), .C1(new_n768), .C2(new_n769), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n771), .A2(new_n773), .A3(new_n760), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n764), .B1(new_n774), .B2(new_n775), .ZN(G1337gat));
  OAI21_X1  g575(.A(G99gat), .B1(new_n742), .B2(new_n531), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n358), .A2(G99gat), .A3(new_n656), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n750), .A2(new_n754), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1338gat));
  NOR3_X1   g579(.A1(new_n483), .A2(G106gat), .A3(new_n656), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n770), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n696), .A2(new_n417), .A3(new_n698), .A4(new_n741), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n783), .A2(G106gat), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT53), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n783), .A2(KEYINPUT110), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n783), .A2(KEYINPUT110), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n786), .A2(new_n787), .A3(new_n360), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n750), .A2(new_n754), .A3(new_n781), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n785), .B1(new_n788), .B2(new_n791), .ZN(G1339gat));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n793), .B(new_n634), .C1(new_n647), .C2(new_n643), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n653), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n793), .B1(new_n651), .B2(new_n635), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n649), .B2(new_n796), .ZN(new_n797));
  AOI22_X1  g596(.A1(new_n797), .A2(KEYINPUT55), .B1(new_n649), .B2(new_n638), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT111), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n797), .A2(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n649), .A2(new_n796), .ZN(new_n801));
  INV_X1    g600(.A(new_n795), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(KEYINPUT55), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n650), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n800), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n245), .A2(new_n246), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n240), .B2(new_n242), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n205), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n255), .A2(new_n809), .ZN(new_n810));
  AND4_X1   g609(.A1(new_n581), .A2(new_n799), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n806), .A2(new_n256), .A3(new_n799), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n655), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n581), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n700), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n624), .A2(new_n257), .A3(new_n656), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n497), .A2(new_n477), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n351), .A2(new_n488), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n819), .A2(new_n820), .A3(new_n417), .ZN(new_n821));
  INV_X1    g620(.A(G113gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n822), .A3(new_n256), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n817), .A2(new_n818), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n418), .ZN(new_n825));
  OAI21_X1  g624(.A(G113gat), .B1(new_n825), .B2(new_n257), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(KEYINPUT112), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(KEYINPUT112), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n823), .B1(new_n827), .B2(new_n828), .ZN(G1340gat));
  AOI21_X1  g628(.A(G120gat), .B1(new_n821), .B2(new_n655), .ZN(new_n830));
  INV_X1    g629(.A(new_n825), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n655), .A2(G120gat), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(G1341gat));
  OAI21_X1  g632(.A(G127gat), .B1(new_n825), .B2(new_n700), .ZN(new_n834));
  INV_X1    g633(.A(G127gat), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n821), .A2(new_n835), .A3(new_n622), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(G1342gat));
  NOR2_X1   g636(.A1(new_n820), .A2(new_n417), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n677), .A2(G134gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n840), .A2(KEYINPUT56), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n819), .A2(new_n677), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n418), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(G134gat), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(KEYINPUT56), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n841), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT113), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n841), .A2(new_n848), .A3(new_n844), .A4(new_n845), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(G1343gat));
  NAND2_X1  g649(.A1(new_n531), .A2(new_n818), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n851), .B(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n483), .B1(new_n815), .B2(new_n816), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XOR2_X1   g655(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n797), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT116), .B1(new_n804), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n801), .A2(new_n802), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n857), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n798), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n860), .A2(new_n256), .A3(new_n864), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n865), .A2(KEYINPUT117), .A3(new_n813), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT117), .B1(new_n865), .B2(new_n813), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n866), .A2(new_n867), .A3(new_n581), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n623), .B1(new_n868), .B2(new_n811), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n483), .B1(new_n869), .B2(new_n816), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n256), .B(new_n856), .C1(new_n870), .C2(new_n855), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n867), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n865), .A2(new_n813), .A3(KEYINPUT117), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n677), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n811), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n622), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n816), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n417), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT57), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n881), .A2(KEYINPUT120), .A3(new_n256), .A4(new_n856), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n873), .A2(G141gat), .A3(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n854), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n257), .A2(G141gat), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n885), .B(KEYINPUT118), .Z(new_n886));
  NOR3_X1   g685(.A1(new_n884), .A2(new_n851), .A3(new_n886), .ZN(new_n887));
  XOR2_X1   g686(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n888));
  NOR2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n871), .A2(G141gat), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT58), .B1(new_n891), .B2(new_n887), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1344gat));
  NOR2_X1   g692(.A1(new_n884), .A2(new_n851), .ZN(new_n894));
  INV_X1    g693(.A(G148gat), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n895), .A3(new_n655), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n817), .A2(new_n855), .A3(new_n417), .ZN(new_n897));
  INV_X1    g696(.A(new_n853), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n899), .B1(KEYINPUT57), .B2(new_n880), .ZN(new_n900));
  AOI211_X1 g699(.A(KEYINPUT59), .B(new_n895), .C1(new_n900), .C2(new_n655), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n867), .A2(new_n581), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n811), .B1(new_n903), .B2(new_n875), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n816), .B1(new_n904), .B2(new_n622), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT57), .B1(new_n905), .B2(new_n417), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n884), .A2(new_n855), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n655), .B(new_n898), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n902), .B1(new_n908), .B2(G148gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n896), .B1(new_n901), .B2(new_n909), .ZN(G1345gat));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n364), .A3(new_n622), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n900), .A2(new_n701), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(new_n364), .ZN(G1346gat));
  NOR2_X1   g712(.A1(new_n687), .A2(new_n483), .ZN(new_n914));
  AOI21_X1  g713(.A(G162gat), .B1(new_n842), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n677), .A2(new_n365), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n900), .B2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n485), .A2(new_n500), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n817), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n418), .ZN(new_n920));
  OAI21_X1  g719(.A(G169gat), .B1(new_n920), .B2(new_n257), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n838), .ZN(new_n922));
  INV_X1    g721(.A(G169gat), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n256), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(new_n926), .ZN(G1348gat));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n655), .A2(G176gat), .ZN(new_n929));
  OR3_X1    g728(.A1(new_n920), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(G176gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n931), .B1(new_n922), .B2(new_n656), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n928), .B1(new_n920), .B2(new_n929), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n930), .A2(KEYINPUT123), .A3(new_n932), .A4(new_n933), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1349gat));
  OAI21_X1  g737(.A(G183gat), .B1(new_n920), .B2(new_n700), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n622), .A2(new_n295), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n922), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g741(.A(G190gat), .B1(new_n920), .B2(new_n677), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n581), .A2(new_n292), .ZN(new_n946));
  OAI22_X1  g745(.A1(new_n944), .A2(new_n945), .B1(new_n922), .B2(new_n946), .ZN(G1351gat));
  XNOR2_X1  g746(.A(KEYINPUT125), .B(G197gat), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n906), .A2(new_n907), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n531), .A2(new_n918), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT126), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n949), .B1(new_n954), .B2(new_n257), .ZN(new_n955));
  OR3_X1    g754(.A1(new_n884), .A2(KEYINPUT124), .A3(new_n951), .ZN(new_n956));
  OAI21_X1  g755(.A(KEYINPUT124), .B1(new_n884), .B2(new_n951), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n256), .A3(new_n948), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n955), .A2(new_n959), .ZN(G1352gat));
  NAND3_X1  g759(.A1(new_n950), .A2(new_n655), .A3(new_n953), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G204gat), .ZN(new_n962));
  NOR4_X1   g761(.A1(new_n884), .A2(G204gat), .A3(new_n656), .A4(new_n951), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT62), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(G1353gat));
  NOR2_X1   g764(.A1(new_n623), .A2(G211gat), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n956), .A2(new_n957), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT127), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n956), .A2(new_n969), .A3(new_n957), .A4(new_n966), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n622), .B(new_n953), .C1(new_n906), .C2(new_n907), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(G211gat), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(KEYINPUT63), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT63), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n972), .A2(new_n975), .A3(G211gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n971), .A2(new_n974), .A3(new_n976), .ZN(G1354gat));
  OAI21_X1  g776(.A(G218gat), .B1(new_n954), .B2(new_n677), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n958), .A2(new_n380), .A3(new_n581), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1355gat));
endmodule


