

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U549 ( .A1(n747), .A2(n746), .ZN(n748) );
  INV_X1 U550 ( .A(n720), .ZN(n713) );
  BUF_X1 U551 ( .A(n720), .Z(n729) );
  NAND2_X1 U552 ( .A1(G8), .A2(n720), .ZN(n810) );
  INV_X1 U553 ( .A(KEYINPUT17), .ZN(n516) );
  NOR2_X2 U554 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  NOR2_X2 U555 ( .A1(n521), .A2(G2105), .ZN(n890) );
  XNOR2_X2 U556 ( .A(KEYINPUT79), .B(n600), .ZN(n696) );
  XNOR2_X1 U557 ( .A(n728), .B(n727), .ZN(n741) );
  INV_X1 U558 ( .A(KEYINPUT31), .ZN(n727) );
  NOR2_X1 U559 ( .A1(n726), .A2(n725), .ZN(n728) );
  AND2_X1 U560 ( .A1(n741), .A2(n734), .ZN(n733) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n709) );
  NOR2_X1 U562 ( .A1(G164), .A2(G1384), .ZN(n784) );
  INV_X1 U563 ( .A(n810), .ZN(n758) );
  NOR2_X1 U564 ( .A1(n801), .A2(n515), .ZN(n802) );
  BUF_X1 U565 ( .A(n527), .Z(n889) );
  AND2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n893) );
  XOR2_X1 U567 ( .A(n707), .B(KEYINPUT28), .Z(n514) );
  XNOR2_X2 U568 ( .A(n683), .B(n682), .ZN(n782) );
  NAND2_X1 U569 ( .A1(n953), .A2(n800), .ZN(n515) );
  XNOR2_X1 U570 ( .A(KEYINPUT97), .B(KEYINPUT26), .ZN(n685) );
  XNOR2_X1 U571 ( .A(n686), .B(n685), .ZN(n687) );
  INV_X1 U572 ( .A(KEYINPUT98), .ZN(n690) );
  NOR2_X1 U573 ( .A1(G1966), .A2(n810), .ZN(n744) );
  INV_X1 U574 ( .A(KEYINPUT101), .ZN(n753) );
  NAND2_X1 U575 ( .A1(n681), .A2(G40), .ZN(n683) );
  XNOR2_X1 U576 ( .A(G2104), .B(KEYINPUT64), .ZN(n518) );
  XNOR2_X1 U577 ( .A(G543), .B(KEYINPUT0), .ZN(n538) );
  NAND2_X1 U578 ( .A1(n651), .A2(G56), .ZN(n580) );
  INV_X1 U579 ( .A(n518), .ZN(n521) );
  INV_X1 U580 ( .A(KEYINPUT1), .ZN(n546) );
  NOR2_X1 U581 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U582 ( .A(n591), .B(KEYINPUT77), .ZN(n961) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(n527) );
  NAND2_X1 U584 ( .A1(G138), .A2(n889), .ZN(n520) );
  NAND2_X1 U585 ( .A1(G102), .A2(n890), .ZN(n519) );
  NAND2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n526) );
  NAND2_X1 U587 ( .A1(G114), .A2(n893), .ZN(n524) );
  NAND2_X1 U588 ( .A1(G2105), .A2(n521), .ZN(n522) );
  XNOR2_X2 U589 ( .A(n522), .B(KEYINPUT65), .ZN(n895) );
  NAND2_X1 U590 ( .A1(G126), .A2(n895), .ZN(n523) );
  NAND2_X1 U591 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U592 ( .A1(n526), .A2(n525), .ZN(G164) );
  NAND2_X1 U593 ( .A1(n527), .A2(G137), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n528), .B(KEYINPUT66), .ZN(n530) );
  NAND2_X1 U595 ( .A1(G113), .A2(n893), .ZN(n529) );
  NAND2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n531), .B(KEYINPUT67), .ZN(n533) );
  NAND2_X1 U598 ( .A1(n895), .A2(G125), .ZN(n532) );
  NAND2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n536) );
  NAND2_X1 U600 ( .A1(G101), .A2(n890), .ZN(n534) );
  XNOR2_X1 U601 ( .A(KEYINPUT23), .B(n534), .ZN(n535) );
  NOR2_X2 U602 ( .A1(n536), .A2(n535), .ZN(n681) );
  BUF_X1 U603 ( .A(n681), .Z(G160) );
  XNOR2_X1 U604 ( .A(KEYINPUT9), .B(KEYINPUT73), .ZN(n543) );
  NOR2_X1 U605 ( .A1(G543), .A2(G651), .ZN(n639) );
  NAND2_X1 U606 ( .A1(n639), .A2(G90), .ZN(n541) );
  INV_X1 U607 ( .A(n538), .ZN(n539) );
  XNOR2_X1 U608 ( .A(KEYINPUT68), .B(n539), .ZN(n653) );
  XNOR2_X1 U609 ( .A(KEYINPUT69), .B(G651), .ZN(n545) );
  NOR2_X2 U610 ( .A1(n653), .A2(n545), .ZN(n637) );
  NAND2_X1 U611 ( .A1(G77), .A2(n637), .ZN(n540) );
  NAND2_X1 U612 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U613 ( .A(n543), .B(n542), .ZN(n552) );
  NOR2_X2 U614 ( .A1(G651), .A2(n653), .ZN(n647) );
  NAND2_X1 U615 ( .A1(G52), .A2(n647), .ZN(n544) );
  XNOR2_X1 U616 ( .A(n544), .B(KEYINPUT72), .ZN(n550) );
  NOR2_X1 U617 ( .A1(G543), .A2(n545), .ZN(n547) );
  XNOR2_X2 U618 ( .A(n547), .B(n546), .ZN(n651) );
  NAND2_X1 U619 ( .A1(G64), .A2(n651), .ZN(n548) );
  XOR2_X1 U620 ( .A(KEYINPUT71), .B(n548), .Z(n549) );
  NAND2_X1 U621 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U622 ( .A1(n552), .A2(n551), .ZN(G171) );
  AND2_X1 U623 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U624 ( .A1(n647), .A2(G53), .ZN(n554) );
  NAND2_X1 U625 ( .A1(G78), .A2(n637), .ZN(n553) );
  NAND2_X1 U626 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U627 ( .A1(n639), .A2(G91), .ZN(n556) );
  NAND2_X1 U628 ( .A1(G65), .A2(n651), .ZN(n555) );
  NAND2_X1 U629 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U630 ( .A1(n558), .A2(n557), .ZN(n706) );
  INV_X1 U631 ( .A(n706), .ZN(G299) );
  INV_X1 U632 ( .A(G57), .ZN(G237) );
  INV_X1 U633 ( .A(G132), .ZN(G219) );
  NAND2_X1 U634 ( .A1(G50), .A2(n647), .ZN(n560) );
  NAND2_X1 U635 ( .A1(G88), .A2(n639), .ZN(n559) );
  NAND2_X1 U636 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U637 ( .A1(G75), .A2(n637), .ZN(n562) );
  NAND2_X1 U638 ( .A1(G62), .A2(n651), .ZN(n561) );
  NAND2_X1 U639 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U640 ( .A1(n564), .A2(n563), .ZN(G166) );
  NAND2_X1 U641 ( .A1(G89), .A2(n639), .ZN(n565) );
  XNOR2_X1 U642 ( .A(n565), .B(KEYINPUT4), .ZN(n566) );
  XNOR2_X1 U643 ( .A(n566), .B(KEYINPUT80), .ZN(n568) );
  NAND2_X1 U644 ( .A1(G76), .A2(n637), .ZN(n567) );
  NAND2_X1 U645 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U646 ( .A(KEYINPUT5), .B(n569), .ZN(n575) );
  XNOR2_X1 U647 ( .A(KEYINPUT81), .B(KEYINPUT6), .ZN(n573) );
  NAND2_X1 U648 ( .A1(G51), .A2(n647), .ZN(n571) );
  NAND2_X1 U649 ( .A1(G63), .A2(n651), .ZN(n570) );
  NAND2_X1 U650 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U651 ( .A(n573), .B(n572), .ZN(n574) );
  NAND2_X1 U652 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U653 ( .A(KEYINPUT7), .B(n576), .ZN(G168) );
  XOR2_X1 U654 ( .A(G168), .B(KEYINPUT8), .Z(n577) );
  XNOR2_X1 U655 ( .A(KEYINPUT82), .B(n577), .ZN(G286) );
  NAND2_X1 U656 ( .A1(G7), .A2(G661), .ZN(n578) );
  XNOR2_X1 U657 ( .A(n578), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U658 ( .A(G223), .ZN(n836) );
  NAND2_X1 U659 ( .A1(n836), .A2(G567), .ZN(n579) );
  XOR2_X1 U660 ( .A(KEYINPUT11), .B(n579), .Z(G234) );
  XOR2_X1 U661 ( .A(KEYINPUT14), .B(n580), .Z(n590) );
  NAND2_X1 U662 ( .A1(n639), .A2(G81), .ZN(n581) );
  XNOR2_X1 U663 ( .A(n581), .B(KEYINPUT12), .ZN(n583) );
  NAND2_X1 U664 ( .A1(G68), .A2(n637), .ZN(n582) );
  NAND2_X1 U665 ( .A1(n583), .A2(n582), .ZN(n585) );
  XOR2_X1 U666 ( .A(KEYINPUT75), .B(KEYINPUT13), .Z(n584) );
  XNOR2_X1 U667 ( .A(n585), .B(n584), .ZN(n588) );
  NAND2_X1 U668 ( .A1(G43), .A2(n647), .ZN(n586) );
  XNOR2_X1 U669 ( .A(n586), .B(KEYINPUT76), .ZN(n587) );
  NAND2_X1 U670 ( .A1(n588), .A2(n587), .ZN(n589) );
  INV_X1 U671 ( .A(G860), .ZN(n622) );
  OR2_X1 U672 ( .A1(n961), .A2(n622), .ZN(G153) );
  INV_X1 U673 ( .A(G171), .ZN(G301) );
  NAND2_X1 U674 ( .A1(G868), .A2(G301), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n639), .A2(G92), .ZN(n593) );
  NAND2_X1 U676 ( .A1(G66), .A2(n651), .ZN(n592) );
  NAND2_X1 U677 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U678 ( .A(KEYINPUT78), .B(n594), .ZN(n598) );
  NAND2_X1 U679 ( .A1(n647), .A2(G54), .ZN(n596) );
  NAND2_X1 U680 ( .A1(G79), .A2(n637), .ZN(n595) );
  NAND2_X1 U681 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U682 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U683 ( .A(KEYINPUT15), .B(n599), .Z(n600) );
  INV_X1 U684 ( .A(G868), .ZN(n665) );
  NAND2_X1 U685 ( .A1(n696), .A2(n665), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n602), .A2(n601), .ZN(G284) );
  NAND2_X1 U687 ( .A1(G868), .A2(G286), .ZN(n604) );
  NAND2_X1 U688 ( .A1(G299), .A2(n665), .ZN(n603) );
  NAND2_X1 U689 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U690 ( .A1(n622), .A2(G559), .ZN(n605) );
  INV_X1 U691 ( .A(n696), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n605), .A2(n620), .ZN(n606) );
  XNOR2_X1 U693 ( .A(n606), .B(KEYINPUT16), .ZN(G148) );
  OR2_X1 U694 ( .A1(G559), .A2(n696), .ZN(n607) );
  NAND2_X1 U695 ( .A1(n607), .A2(G868), .ZN(n609) );
  NAND2_X1 U696 ( .A1(n961), .A2(n665), .ZN(n608) );
  NAND2_X1 U697 ( .A1(n609), .A2(n608), .ZN(G282) );
  NAND2_X1 U698 ( .A1(G111), .A2(n893), .ZN(n611) );
  NAND2_X1 U699 ( .A1(G135), .A2(n889), .ZN(n610) );
  NAND2_X1 U700 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U701 ( .A1(n895), .A2(G123), .ZN(n612) );
  XOR2_X1 U702 ( .A(KEYINPUT18), .B(n612), .Z(n613) );
  NOR2_X1 U703 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U704 ( .A1(n890), .A2(G99), .ZN(n615) );
  NAND2_X1 U705 ( .A1(n616), .A2(n615), .ZN(n1018) );
  XNOR2_X1 U706 ( .A(n1018), .B(G2096), .ZN(n617) );
  XNOR2_X1 U707 ( .A(n617), .B(KEYINPUT83), .ZN(n619) );
  INV_X1 U708 ( .A(G2100), .ZN(n618) );
  NAND2_X1 U709 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U710 ( .A1(G559), .A2(n620), .ZN(n621) );
  XOR2_X1 U711 ( .A(n961), .B(n621), .Z(n662) );
  NAND2_X1 U712 ( .A1(n622), .A2(n662), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n647), .A2(G55), .ZN(n624) );
  NAND2_X1 U714 ( .A1(G80), .A2(n637), .ZN(n623) );
  NAND2_X1 U715 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U716 ( .A1(n639), .A2(G93), .ZN(n626) );
  NAND2_X1 U717 ( .A1(G67), .A2(n651), .ZN(n625) );
  NAND2_X1 U718 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U719 ( .A1(n628), .A2(n627), .ZN(n664) );
  XOR2_X1 U720 ( .A(n629), .B(n664), .Z(G145) );
  NAND2_X1 U721 ( .A1(G47), .A2(n647), .ZN(n631) );
  NAND2_X1 U722 ( .A1(G85), .A2(n639), .ZN(n630) );
  NAND2_X1 U723 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U724 ( .A1(n637), .A2(G72), .ZN(n632) );
  XOR2_X1 U725 ( .A(KEYINPUT70), .B(n632), .Z(n633) );
  NOR2_X1 U726 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U727 ( .A1(G60), .A2(n651), .ZN(n635) );
  NAND2_X1 U728 ( .A1(n636), .A2(n635), .ZN(G290) );
  NAND2_X1 U729 ( .A1(n637), .A2(G73), .ZN(n638) );
  XOR2_X1 U730 ( .A(KEYINPUT2), .B(n638), .Z(n644) );
  NAND2_X1 U731 ( .A1(n639), .A2(G86), .ZN(n641) );
  NAND2_X1 U732 ( .A1(G61), .A2(n651), .ZN(n640) );
  NAND2_X1 U733 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U734 ( .A(KEYINPUT85), .B(n642), .Z(n643) );
  NOR2_X1 U735 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U736 ( .A1(n647), .A2(G48), .ZN(n645) );
  NAND2_X1 U737 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U738 ( .A1(G49), .A2(n647), .ZN(n649) );
  NAND2_X1 U739 ( .A1(G74), .A2(G651), .ZN(n648) );
  NAND2_X1 U740 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U741 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U742 ( .A(n652), .B(KEYINPUT84), .ZN(n655) );
  NAND2_X1 U743 ( .A1(G87), .A2(n653), .ZN(n654) );
  NAND2_X1 U744 ( .A1(n655), .A2(n654), .ZN(G288) );
  XOR2_X1 U745 ( .A(G305), .B(G288), .Z(n656) );
  XNOR2_X1 U746 ( .A(G290), .B(n656), .ZN(n659) );
  XNOR2_X1 U747 ( .A(G166), .B(KEYINPUT19), .ZN(n657) );
  XNOR2_X1 U748 ( .A(n657), .B(KEYINPUT86), .ZN(n658) );
  XOR2_X1 U749 ( .A(n659), .B(n658), .Z(n661) );
  XNOR2_X1 U750 ( .A(n706), .B(n664), .ZN(n660) );
  XNOR2_X1 U751 ( .A(n661), .B(n660), .ZN(n904) );
  XOR2_X1 U752 ( .A(n904), .B(n662), .Z(n663) );
  NOR2_X1 U753 ( .A1(n665), .A2(n663), .ZN(n667) );
  AND2_X1 U754 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U755 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U756 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U757 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U758 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U759 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U760 ( .A1(n671), .A2(G2072), .ZN(G158) );
  XOR2_X1 U761 ( .A(KEYINPUT74), .B(G82), .Z(G220) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U763 ( .A1(G220), .A2(G219), .ZN(n672) );
  XNOR2_X1 U764 ( .A(KEYINPUT22), .B(n672), .ZN(n673) );
  NAND2_X1 U765 ( .A1(n673), .A2(G96), .ZN(n674) );
  NOR2_X1 U766 ( .A1(n674), .A2(G218), .ZN(n675) );
  XNOR2_X1 U767 ( .A(n675), .B(KEYINPUT87), .ZN(n841) );
  NAND2_X1 U768 ( .A1(n841), .A2(G2106), .ZN(n679) );
  NAND2_X1 U769 ( .A1(G69), .A2(G120), .ZN(n676) );
  NOR2_X1 U770 ( .A1(G237), .A2(n676), .ZN(n677) );
  NAND2_X1 U771 ( .A1(G108), .A2(n677), .ZN(n842) );
  NAND2_X1 U772 ( .A1(n842), .A2(G567), .ZN(n678) );
  NAND2_X1 U773 ( .A1(n679), .A2(n678), .ZN(n861) );
  NAND2_X1 U774 ( .A1(G483), .A2(G661), .ZN(n680) );
  NOR2_X1 U775 ( .A1(n861), .A2(n680), .ZN(n840) );
  NAND2_X1 U776 ( .A1(n840), .A2(G36), .ZN(G176) );
  INV_X1 U777 ( .A(G166), .ZN(G303) );
  INV_X1 U778 ( .A(KEYINPUT88), .ZN(n682) );
  AND2_X1 U779 ( .A1(n784), .A2(G1996), .ZN(n684) );
  NAND2_X1 U780 ( .A1(n782), .A2(n684), .ZN(n686) );
  NOR2_X1 U781 ( .A1(n687), .A2(n961), .ZN(n689) );
  NAND2_X1 U782 ( .A1(n784), .A2(n782), .ZN(n720) );
  NAND2_X1 U783 ( .A1(G1341), .A2(n729), .ZN(n688) );
  NAND2_X1 U784 ( .A1(n689), .A2(n688), .ZN(n697) );
  NOR2_X1 U785 ( .A1(n697), .A2(n696), .ZN(n691) );
  XNOR2_X1 U786 ( .A(n691), .B(n690), .ZN(n695) );
  NOR2_X1 U787 ( .A1(G2067), .A2(n729), .ZN(n693) );
  NOR2_X1 U788 ( .A1(n713), .A2(G1348), .ZN(n692) );
  NOR2_X1 U789 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U790 ( .A1(n695), .A2(n694), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n704) );
  NAND2_X1 U793 ( .A1(n713), .A2(G2072), .ZN(n700) );
  XNOR2_X1 U794 ( .A(n700), .B(KEYINPUT27), .ZN(n702) );
  INV_X1 U795 ( .A(G1956), .ZN(n984) );
  NOR2_X1 U796 ( .A1(n984), .A2(n713), .ZN(n701) );
  NOR2_X1 U797 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n703) );
  NAND2_X1 U799 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U800 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n708), .A2(n514), .ZN(n710) );
  XNOR2_X1 U802 ( .A(n710), .B(n709), .ZN(n719) );
  XOR2_X1 U803 ( .A(G2078), .B(KEYINPUT25), .Z(n940) );
  NOR2_X1 U804 ( .A1(n940), .A2(n720), .ZN(n712) );
  INV_X1 U805 ( .A(KEYINPUT95), .ZN(n711) );
  XNOR2_X1 U806 ( .A(n712), .B(n711), .ZN(n715) );
  NOR2_X1 U807 ( .A1(n713), .A2(G1961), .ZN(n714) );
  NOR2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n717) );
  INV_X1 U809 ( .A(KEYINPUT96), .ZN(n716) );
  XNOR2_X1 U810 ( .A(n717), .B(n716), .ZN(n724) );
  NAND2_X1 U811 ( .A1(G171), .A2(n724), .ZN(n718) );
  NAND2_X1 U812 ( .A1(n719), .A2(n718), .ZN(n742) );
  NOR2_X1 U813 ( .A1(G2084), .A2(n729), .ZN(n743) );
  NOR2_X1 U814 ( .A1(n744), .A2(n743), .ZN(n721) );
  NAND2_X1 U815 ( .A1(n721), .A2(G8), .ZN(n722) );
  XNOR2_X1 U816 ( .A(n722), .B(KEYINPUT30), .ZN(n723) );
  NOR2_X1 U817 ( .A1(G168), .A2(n723), .ZN(n726) );
  NOR2_X1 U818 ( .A1(n724), .A2(G171), .ZN(n725) );
  NOR2_X1 U819 ( .A1(G1971), .A2(n810), .ZN(n731) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n729), .ZN(n730) );
  NOR2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U822 ( .A1(n732), .A2(G303), .ZN(n734) );
  NAND2_X1 U823 ( .A1(n742), .A2(n733), .ZN(n738) );
  INV_X1 U824 ( .A(n734), .ZN(n735) );
  OR2_X1 U825 ( .A1(n735), .A2(G286), .ZN(n736) );
  AND2_X1 U826 ( .A1(n736), .A2(G8), .ZN(n737) );
  NAND2_X1 U827 ( .A1(n738), .A2(n737), .ZN(n740) );
  XOR2_X1 U828 ( .A(KEYINPUT99), .B(KEYINPUT32), .Z(n739) );
  XNOR2_X1 U829 ( .A(n740), .B(n739), .ZN(n749) );
  AND2_X1 U830 ( .A1(n742), .A2(n741), .ZN(n747) );
  AND2_X1 U831 ( .A1(G8), .A2(n743), .ZN(n745) );
  OR2_X1 U832 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U833 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U834 ( .A(n750), .B(KEYINPUT100), .ZN(n808) );
  NOR2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n969) );
  NOR2_X1 U836 ( .A1(G1971), .A2(G303), .ZN(n751) );
  NOR2_X1 U837 ( .A1(n969), .A2(n751), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n808), .A2(n752), .ZN(n754) );
  XNOR2_X1 U839 ( .A(n754), .B(n753), .ZN(n755) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n966) );
  NAND2_X1 U841 ( .A1(n755), .A2(n966), .ZN(n756) );
  XNOR2_X1 U842 ( .A(n756), .B(KEYINPUT102), .ZN(n757) );
  INV_X1 U843 ( .A(n757), .ZN(n759) );
  NAND2_X1 U844 ( .A1(n759), .A2(n758), .ZN(n761) );
  INV_X1 U845 ( .A(KEYINPUT33), .ZN(n760) );
  NAND2_X1 U846 ( .A1(n761), .A2(n760), .ZN(n803) );
  NAND2_X1 U847 ( .A1(n969), .A2(KEYINPUT33), .ZN(n762) );
  NOR2_X1 U848 ( .A1(n762), .A2(n810), .ZN(n801) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n953) );
  NAND2_X1 U850 ( .A1(n893), .A2(G117), .ZN(n764) );
  NAND2_X1 U851 ( .A1(n889), .A2(G141), .ZN(n763) );
  NAND2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n890), .A2(G105), .ZN(n765) );
  XOR2_X1 U854 ( .A(KEYINPUT38), .B(n765), .Z(n766) );
  NOR2_X1 U855 ( .A1(n767), .A2(n766), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n895), .A2(G129), .ZN(n768) );
  NAND2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n882) );
  AND2_X1 U858 ( .A1(n882), .A2(G1996), .ZN(n781) );
  INV_X1 U859 ( .A(G1991), .ZN(n779) );
  NAND2_X1 U860 ( .A1(G107), .A2(n893), .ZN(n771) );
  NAND2_X1 U861 ( .A1(G95), .A2(n890), .ZN(n770) );
  NAND2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U863 ( .A1(G119), .A2(n895), .ZN(n772) );
  XNOR2_X1 U864 ( .A(KEYINPUT93), .B(n772), .ZN(n773) );
  NOR2_X1 U865 ( .A1(n774), .A2(n773), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n889), .A2(G131), .ZN(n775) );
  NAND2_X1 U867 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U868 ( .A(KEYINPUT94), .B(n777), .ZN(n886) );
  INV_X1 U869 ( .A(n886), .ZN(n778) );
  NOR2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n1009) );
  INV_X1 U872 ( .A(n782), .ZN(n783) );
  NOR2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U874 ( .A(n785), .B(KEYINPUT89), .ZN(n831) );
  NOR2_X1 U875 ( .A1(n1009), .A2(n831), .ZN(n825) );
  INV_X1 U876 ( .A(n825), .ZN(n799) );
  INV_X1 U877 ( .A(n831), .ZN(n797) );
  NAND2_X1 U878 ( .A1(n893), .A2(G116), .ZN(n786) );
  XNOR2_X1 U879 ( .A(n786), .B(KEYINPUT92), .ZN(n788) );
  NAND2_X1 U880 ( .A1(G128), .A2(n895), .ZN(n787) );
  NAND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U882 ( .A(KEYINPUT35), .B(n789), .ZN(n795) );
  NAND2_X1 U883 ( .A1(n890), .A2(G104), .ZN(n790) );
  XOR2_X1 U884 ( .A(KEYINPUT91), .B(n790), .Z(n792) );
  NAND2_X1 U885 ( .A1(n889), .A2(G140), .ZN(n791) );
  NAND2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U887 ( .A(KEYINPUT34), .B(n793), .Z(n794) );
  NAND2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U889 ( .A(KEYINPUT36), .B(n796), .Z(n880) );
  XNOR2_X1 U890 ( .A(G2067), .B(KEYINPUT37), .ZN(n822) );
  NOR2_X1 U891 ( .A1(n880), .A2(n822), .ZN(n1015) );
  NAND2_X1 U892 ( .A1(n797), .A2(n1015), .ZN(n798) );
  NAND2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n815) );
  INV_X1 U894 ( .A(n815), .ZN(n800) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n817) );
  NOR2_X1 U896 ( .A1(G1981), .A2(G305), .ZN(n804) );
  XOR2_X1 U897 ( .A(n804), .B(KEYINPUT24), .Z(n805) );
  OR2_X1 U898 ( .A1(n810), .A2(n805), .ZN(n813) );
  NOR2_X1 U899 ( .A1(G2090), .A2(G303), .ZN(n806) );
  XOR2_X1 U900 ( .A(KEYINPUT103), .B(n806), .Z(n807) );
  NAND2_X1 U901 ( .A1(G8), .A2(n807), .ZN(n809) );
  NAND2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n812) );
  AND2_X1 U904 ( .A1(n813), .A2(n812), .ZN(n814) );
  OR2_X1 U905 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U906 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U907 ( .A(n818), .B(KEYINPUT104), .ZN(n821) );
  XOR2_X1 U908 ( .A(G1986), .B(G290), .Z(n973) );
  NOR2_X1 U909 ( .A1(n973), .A2(n831), .ZN(n819) );
  XOR2_X1 U910 ( .A(KEYINPUT90), .B(n819), .Z(n820) );
  NAND2_X1 U911 ( .A1(n821), .A2(n820), .ZN(n834) );
  AND2_X1 U912 ( .A1(n880), .A2(n822), .ZN(n1017) );
  NOR2_X1 U913 ( .A1(G1996), .A2(n882), .ZN(n1012) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n823) );
  NOR2_X1 U915 ( .A1(n886), .A2(G1991), .ZN(n1016) );
  NOR2_X1 U916 ( .A1(n823), .A2(n1016), .ZN(n824) );
  NOR2_X1 U917 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U918 ( .A1(n1012), .A2(n826), .ZN(n827) );
  XOR2_X1 U919 ( .A(KEYINPUT39), .B(n827), .Z(n828) );
  NOR2_X1 U920 ( .A1(n1015), .A2(n828), .ZN(n829) );
  NOR2_X1 U921 ( .A1(n1017), .A2(n829), .ZN(n830) );
  NOR2_X1 U922 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U923 ( .A(KEYINPUT105), .B(n832), .ZN(n833) );
  NAND2_X1 U924 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U925 ( .A(n835), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U926 ( .A1(n836), .A2(G2106), .ZN(n837) );
  XNOR2_X1 U927 ( .A(n837), .B(KEYINPUT108), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U929 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U931 ( .A1(n840), .A2(n839), .ZN(G188) );
  INV_X1 U933 ( .A(G120), .ZN(G236) );
  INV_X1 U934 ( .A(G96), .ZN(G221) );
  INV_X1 U935 ( .A(G69), .ZN(G235) );
  NOR2_X1 U936 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  XOR2_X1 U938 ( .A(G2100), .B(G2096), .Z(n844) );
  XNOR2_X1 U939 ( .A(KEYINPUT42), .B(G2678), .ZN(n843) );
  XNOR2_X1 U940 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U941 ( .A(KEYINPUT43), .B(G2067), .Z(n846) );
  XNOR2_X1 U942 ( .A(G2090), .B(G2072), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U944 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U945 ( .A(G2078), .B(G2084), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n850), .B(n849), .ZN(G227) );
  XOR2_X1 U947 ( .A(G1986), .B(G1981), .Z(n852) );
  XNOR2_X1 U948 ( .A(G1961), .B(G1956), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U950 ( .A(G1976), .B(G1971), .Z(n854) );
  XNOR2_X1 U951 ( .A(G1991), .B(G1996), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U953 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U954 ( .A(G2474), .B(KEYINPUT109), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(n860) );
  XOR2_X1 U956 ( .A(G1966), .B(KEYINPUT41), .Z(n859) );
  XNOR2_X1 U957 ( .A(n860), .B(n859), .ZN(G229) );
  INV_X1 U958 ( .A(n861), .ZN(G319) );
  NAND2_X1 U959 ( .A1(G112), .A2(n893), .ZN(n863) );
  NAND2_X1 U960 ( .A1(G136), .A2(n889), .ZN(n862) );
  NAND2_X1 U961 ( .A1(n863), .A2(n862), .ZN(n868) );
  NAND2_X1 U962 ( .A1(G124), .A2(n895), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n864), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U964 ( .A1(n890), .A2(G100), .ZN(n865) );
  NAND2_X1 U965 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U966 ( .A1(n868), .A2(n867), .ZN(G162) );
  XOR2_X1 U967 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n879) );
  NAND2_X1 U968 ( .A1(G118), .A2(n893), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G130), .A2(n895), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n876) );
  NAND2_X1 U971 ( .A1(G142), .A2(n889), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G106), .A2(n890), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U974 ( .A(KEYINPUT110), .B(n873), .Z(n874) );
  XNOR2_X1 U975 ( .A(KEYINPUT45), .B(n874), .ZN(n875) );
  NOR2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n877), .B(KEYINPUT112), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n881), .B(n880), .ZN(n884) );
  XOR2_X1 U980 ( .A(n882), .B(G164), .Z(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n1018), .B(n885), .ZN(n888) );
  XNOR2_X1 U983 ( .A(n886), .B(G162), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n902) );
  NAND2_X1 U985 ( .A1(G139), .A2(n889), .ZN(n892) );
  NAND2_X1 U986 ( .A1(G103), .A2(n890), .ZN(n891) );
  NAND2_X1 U987 ( .A1(n892), .A2(n891), .ZN(n900) );
  NAND2_X1 U988 ( .A1(n893), .A2(G115), .ZN(n894) );
  XOR2_X1 U989 ( .A(KEYINPUT111), .B(n894), .Z(n897) );
  NAND2_X1 U990 ( .A1(n895), .A2(G127), .ZN(n896) );
  NAND2_X1 U991 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n898), .Z(n899) );
  NOR2_X1 U993 ( .A1(n900), .A2(n899), .ZN(n1020) );
  XOR2_X1 U994 ( .A(G160), .B(n1020), .Z(n901) );
  XNOR2_X1 U995 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U996 ( .A1(G37), .A2(n903), .ZN(G395) );
  XNOR2_X1 U997 ( .A(G171), .B(KEYINPUT113), .ZN(n907) );
  XNOR2_X1 U998 ( .A(n904), .B(n696), .ZN(n905) );
  XNOR2_X1 U999 ( .A(n905), .B(n961), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1001 ( .A(n908), .B(G286), .Z(n909) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n909), .ZN(G397) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n911), .B(n910), .ZN(n924) );
  XNOR2_X1 U1006 ( .A(G2443), .B(G2427), .ZN(n921) );
  XOR2_X1 U1007 ( .A(G2430), .B(KEYINPUT107), .Z(n913) );
  XNOR2_X1 U1008 ( .A(G2454), .B(G2435), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(n917) );
  XOR2_X1 U1010 ( .A(G2438), .B(KEYINPUT106), .Z(n915) );
  XNOR2_X1 U1011 ( .A(G1341), .B(G1348), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1013 ( .A(n917), .B(n916), .Z(n919) );
  XNOR2_X1 U1014 ( .A(G2451), .B(G2446), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(n919), .B(n918), .ZN(n920) );
  XNOR2_X1 U1016 ( .A(n921), .B(n920), .ZN(n922) );
  NAND2_X1 U1017 ( .A1(n922), .A2(G14), .ZN(n927) );
  NAND2_X1 U1018 ( .A1(G319), .A2(n927), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  INV_X1 U1023 ( .A(G108), .ZN(G238) );
  INV_X1 U1024 ( .A(n927), .ZN(G401) );
  INV_X1 U1025 ( .A(KEYINPUT55), .ZN(n1032) );
  XOR2_X1 U1026 ( .A(G2090), .B(G35), .Z(n930) );
  XOR2_X1 U1027 ( .A(KEYINPUT54), .B(G34), .Z(n928) );
  XNOR2_X1 U1028 ( .A(n928), .B(G2084), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n946) );
  XNOR2_X1 U1030 ( .A(G32), .B(G1996), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(n931), .B(KEYINPUT117), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(G1991), .B(G25), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(G33), .B(G2072), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1035 ( .A1(G28), .A2(n934), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(KEYINPUT116), .B(G2067), .ZN(n935) );
  XNOR2_X1 U1037 ( .A(G26), .B(n935), .ZN(n936) );
  NOR2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(G27), .B(n940), .ZN(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1042 ( .A(KEYINPUT118), .B(n943), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(KEYINPUT53), .B(n944), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(KEYINPUT119), .B(n947), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(n1032), .B(n948), .ZN(n950) );
  INV_X1 U1047 ( .A(G29), .ZN(n949) );
  NAND2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1049 ( .A1(G11), .A2(n951), .ZN(n1008) );
  XNOR2_X1 U1050 ( .A(G16), .B(KEYINPUT56), .ZN(n979) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G168), .ZN(n952) );
  XNOR2_X1 U1052 ( .A(n952), .B(KEYINPUT120), .ZN(n954) );
  NAND2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1054 ( .A(n955), .B(KEYINPUT57), .ZN(n960) );
  XOR2_X1 U1055 ( .A(G1348), .B(KEYINPUT121), .Z(n956) );
  XNOR2_X1 U1056 ( .A(n696), .B(n956), .ZN(n958) );
  XNOR2_X1 U1057 ( .A(G1961), .B(G301), .ZN(n957) );
  NOR2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n964) );
  XOR2_X1 U1060 ( .A(G1341), .B(n961), .Z(n962) );
  XNOR2_X1 U1061 ( .A(KEYINPUT125), .B(n962), .ZN(n963) );
  NOR2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n977) );
  XNOR2_X1 U1063 ( .A(G299), .B(G1956), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(G166), .B(G1971), .ZN(n965) );
  XNOR2_X1 U1065 ( .A(n965), .B(KEYINPUT122), .ZN(n967) );
  NAND2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1068 ( .A(KEYINPUT123), .B(n970), .ZN(n971) );
  NOR2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1071 ( .A(KEYINPUT124), .B(n975), .Z(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n1006) );
  INV_X1 U1074 ( .A(G16), .ZN(n1004) );
  XNOR2_X1 U1075 ( .A(G1966), .B(G21), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(G1961), .B(G5), .ZN(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n993) );
  XOR2_X1 U1078 ( .A(G4), .B(KEYINPUT126), .Z(n983) );
  XNOR2_X1 U1079 ( .A(G1348), .B(KEYINPUT59), .ZN(n982) );
  XNOR2_X1 U1080 ( .A(n983), .B(n982), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(G20), .B(n984), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(G1341), .B(G19), .ZN(n986) );
  XNOR2_X1 U1083 ( .A(G1981), .B(G6), .ZN(n985) );
  NOR2_X1 U1084 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1085 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1086 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1087 ( .A(n991), .B(KEYINPUT60), .ZN(n992) );
  NAND2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(G1971), .B(G22), .ZN(n995) );
  XNOR2_X1 U1090 ( .A(G24), .B(G1986), .ZN(n994) );
  NOR2_X1 U1091 ( .A1(n995), .A2(n994), .ZN(n997) );
  XOR2_X1 U1092 ( .A(G1976), .B(G23), .Z(n996) );
  NAND2_X1 U1093 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1094 ( .A(KEYINPUT58), .B(n998), .ZN(n999) );
  NOR2_X1 U1095 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1096 ( .A(n1001), .B(KEYINPUT61), .Z(n1002) );
  XNOR2_X1 U1097 ( .A(KEYINPUT127), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1098 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1099 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1036) );
  XNOR2_X1 U1101 ( .A(G160), .B(G2084), .ZN(n1010) );
  NAND2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1029) );
  XOR2_X1 U1103 ( .A(G2090), .B(G162), .Z(n1011) );
  NOR2_X1 U1104 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1105 ( .A(n1013), .B(KEYINPUT51), .ZN(n1014) );
  NOR2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1027) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1025) );
  XOR2_X1 U1109 ( .A(G2072), .B(n1020), .Z(n1022) );
  XOR2_X1 U1110 ( .A(G164), .B(G2078), .Z(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1112 ( .A(KEYINPUT50), .B(n1023), .Z(n1024) );
  NOR2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1116 ( .A(KEYINPUT52), .B(n1030), .Z(n1031) );
  XNOR2_X1 U1117 ( .A(KEYINPUT115), .B(n1031), .ZN(n1033) );
  NAND2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1119 ( .A1(n1034), .A2(G29), .ZN(n1035) );
  NAND2_X1 U1120 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XOR2_X1 U1121 ( .A(KEYINPUT62), .B(n1037), .Z(G311) );
  INV_X1 U1122 ( .A(G311), .ZN(G150) );
endmodule

