//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n800,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1020;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G22gat), .B(G78gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G228gat), .A2(G233gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT71), .ZN(new_n206));
  AND2_X1   g005(.A1(KEYINPUT70), .A2(G148gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(KEYINPUT70), .A2(G148gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n206), .B(G141gat), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210));
  INV_X1    g009(.A(G155gat), .ZN(new_n211));
  INV_X1    g010(.A(G162gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G141gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT70), .ZN(new_n217));
  INV_X1    g016(.A(G148gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(KEYINPUT70), .A2(G148gat), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n216), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n216), .A2(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT71), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n209), .B(new_n215), .C1(new_n221), .C2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n218), .A2(G141gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(new_n210), .ZN(new_n228));
  XOR2_X1   g027(.A(G155gat), .B(G162gat), .Z(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n224), .A2(new_n225), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT29), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(G197gat), .A2(G204gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(G197gat), .A2(G204gat), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT22), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G211gat), .ZN(new_n237));
  INV_X1    g036(.A(G218gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n238), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n236), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n237), .A2(new_n238), .A3(KEYINPUT22), .ZN(new_n245));
  OAI22_X1  g044(.A1(new_n245), .A2(new_n239), .B1(new_n235), .B2(new_n234), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n236), .A2(new_n240), .A3(KEYINPUT69), .A4(new_n241), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n244), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT78), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n251), .B1(new_n248), .B2(KEYINPUT29), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n244), .A2(new_n246), .A3(new_n247), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(KEYINPUT78), .A3(new_n232), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n252), .A2(new_n225), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n224), .A2(new_n230), .ZN(new_n256));
  AOI211_X1 g055(.A(new_n205), .B(new_n250), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT29), .B1(new_n242), .B2(new_n246), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n256), .B1(new_n258), .B2(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n249), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT77), .B1(new_n260), .B2(new_n205), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT77), .ZN(new_n262));
  INV_X1    g061(.A(new_n205), .ZN(new_n263));
  AOI211_X1 g062(.A(new_n262), .B(new_n263), .C1(new_n249), .C2(new_n259), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n204), .B1(new_n257), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n254), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT78), .B1(new_n253), .B2(new_n232), .ZN(new_n268));
  NOR3_X1   g067(.A1(new_n267), .A2(new_n268), .A3(KEYINPUT3), .ZN(new_n269));
  OAI21_X1  g068(.A(G141gat), .B1(new_n207), .B2(new_n208), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n206), .B1(new_n216), .B2(G148gat), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n270), .A2(new_n271), .B1(new_n214), .B2(new_n213), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n272), .A2(new_n209), .B1(new_n228), .B2(new_n229), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n263), .B(new_n249), .C1(new_n269), .C2(new_n273), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n275), .A2(new_n256), .B1(new_n233), .B2(new_n248), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n262), .B1(new_n276), .B2(new_n263), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n260), .A2(KEYINPUT77), .A3(new_n205), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n204), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n274), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n203), .B1(new_n266), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n203), .A3(new_n281), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G57gat), .B(G85gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(G1gat), .B(G29gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n288), .B(new_n289), .Z(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G225gat), .A2(G233gat), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G134gat), .ZN(new_n294));
  INV_X1    g093(.A(G127gat), .ZN(new_n295));
  INV_X1    g094(.A(G120gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G113gat), .ZN(new_n297));
  INV_X1    g096(.A(G113gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G120gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT1), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n295), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI211_X1 g101(.A(KEYINPUT1), .B(G127gat), .C1(new_n297), .C2(new_n299), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n294), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G113gat), .B(G120gat), .ZN(new_n305));
  OAI21_X1  g104(.A(G127gat), .B1(new_n305), .B2(KEYINPUT1), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n300), .A2(new_n301), .A3(new_n295), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n307), .A3(G134gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(new_n256), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n273), .B1(new_n308), .B2(new_n304), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n293), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT5), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(new_n309), .A3(new_n231), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT72), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT72), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n314), .A2(new_n309), .A3(new_n317), .A4(new_n231), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n293), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n304), .A2(new_n308), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .A4(new_n273), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n273), .A2(new_n304), .A3(new_n322), .A4(new_n308), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT73), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT4), .B1(new_n309), .B2(new_n256), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n313), .B1(new_n319), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n324), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n224), .A2(new_n225), .A3(new_n230), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n225), .B1(new_n224), .B2(new_n230), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n317), .B1(new_n332), .B2(new_n309), .ZN(new_n333));
  AND4_X1   g132(.A1(new_n317), .A2(new_n314), .A3(new_n309), .A4(new_n231), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n329), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n291), .B1(new_n328), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT5), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n309), .B(new_n256), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(new_n293), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n292), .B1(new_n333), .B2(new_n334), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n323), .A2(new_n326), .A3(new_n325), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n316), .A2(new_n318), .B1(new_n326), .B2(new_n324), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n336), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n290), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT75), .B(KEYINPUT6), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n339), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G8gat), .B(G36gat), .ZN(new_n351));
  INV_X1    g150(.A(G64gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G92gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G169gat), .ZN(new_n357));
  INV_X1    g156(.A(G176gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT66), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT26), .ZN(new_n360));
  AND2_X1   g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(G169gat), .A2(G176gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT26), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(KEYINPUT66), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT28), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT65), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT65), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT28), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT27), .B(G183gat), .ZN(new_n372));
  INV_X1    g171(.A(G190gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT65), .B(KEYINPUT28), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n366), .A2(new_n374), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT23), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(G169gat), .B2(G176gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT24), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n384), .A2(G183gat), .A3(G190gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n380), .A2(KEYINPUT24), .ZN(new_n386));
  NOR2_X1   g185(.A1(G183gat), .A2(G190gat), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n383), .B(new_n385), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n382), .A2(G169gat), .A3(G176gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT64), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n391), .A2(new_n357), .A3(new_n358), .A4(KEYINPUT23), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT25), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n394), .A2(new_n362), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n389), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n361), .B1(KEYINPUT23), .B2(new_n363), .ZN(new_n398));
  INV_X1    g197(.A(G183gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n373), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(KEYINPUT24), .A3(new_n380), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n398), .A2(new_n401), .A3(new_n383), .A4(new_n385), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT25), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n381), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G226gat), .A2(G233gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n232), .A3(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n388), .A2(new_n392), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n407), .A2(new_n396), .B1(new_n402), .B2(KEYINPUT25), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n408), .A2(G226gat), .A3(G233gat), .A4(new_n381), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n406), .A2(new_n253), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n253), .B1(new_n406), .B2(new_n409), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT37), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n406), .A2(new_n409), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n248), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT37), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n406), .A2(new_n409), .A3(new_n253), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n356), .B1(new_n412), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT38), .ZN(new_n419));
  OR2_X1    g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n414), .A2(new_n416), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n418), .A2(new_n419), .B1(new_n421), .B2(new_n356), .ZN(new_n422));
  INV_X1    g221(.A(new_n349), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n291), .B(new_n423), .C1(new_n328), .C2(new_n338), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n350), .A2(new_n420), .A3(new_n422), .A4(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n356), .B1(new_n410), .B2(new_n411), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n414), .A2(new_n416), .A3(new_n355), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n427), .A3(KEYINPUT30), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT30), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n421), .A2(new_n429), .A3(new_n356), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT39), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n341), .A2(new_n293), .ZN(new_n433));
  AOI211_X1 g232(.A(new_n432), .B(new_n433), .C1(new_n293), .C2(new_n335), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n346), .A2(KEYINPUT39), .A3(new_n292), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT79), .B1(new_n435), .B2(new_n291), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n335), .A2(new_n432), .A3(new_n293), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT79), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n438), .A3(new_n290), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n434), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n431), .B1(new_n440), .B2(KEYINPUT40), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n433), .B1(new_n335), .B2(new_n293), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT39), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n437), .A2(new_n438), .A3(new_n290), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n438), .B1(new_n437), .B2(new_n290), .ZN(new_n445));
  OAI211_X1 g244(.A(KEYINPUT40), .B(new_n443), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n339), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n285), .B(new_n425), .C1(new_n441), .C2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT80), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n285), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT76), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n350), .A2(new_n424), .ZN(new_n453));
  INV_X1    g252(.A(new_n431), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI211_X1 g254(.A(KEYINPUT76), .B(new_n431), .C1(new_n350), .C2(new_n424), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n451), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT40), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n460), .A2(new_n339), .A3(new_n431), .A4(new_n446), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n461), .A2(KEYINPUT80), .A3(new_n285), .A4(new_n425), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n408), .A2(new_n308), .A3(new_n304), .A4(new_n381), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n404), .A2(new_n309), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(G227gat), .ZN(new_n467));
  INV_X1    g266(.A(G233gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT68), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(KEYINPUT34), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n466), .A2(KEYINPUT68), .A3(new_n470), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT67), .B(G71gat), .ZN(new_n475));
  INV_X1    g274(.A(G99gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G15gat), .B(G43gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n470), .B1(new_n463), .B2(new_n464), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(KEYINPUT33), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT32), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  AOI221_X4 g283(.A(new_n482), .B1(new_n479), .B2(KEYINPUT33), .C1(new_n465), .C2(new_n469), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n474), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n404), .A2(new_n309), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n404), .A2(new_n309), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n469), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT32), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT33), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n492), .A3(new_n479), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n481), .A2(new_n483), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n473), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n472), .B1(new_n486), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n486), .A2(new_n495), .A3(new_n472), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT36), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n486), .A2(new_n495), .A3(new_n472), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n500), .A2(new_n496), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n450), .A2(new_n457), .A3(new_n462), .A4(new_n503), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n274), .A2(new_n279), .A3(new_n280), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n280), .B1(new_n274), .B2(new_n279), .ZN(new_n506));
  INV_X1    g305(.A(new_n203), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  OAI22_X1  g307(.A1(new_n500), .A2(new_n496), .B1(new_n508), .B2(new_n282), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT35), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n510), .A2(new_n511), .A3(new_n453), .A4(new_n454), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n455), .A2(new_n456), .A3(new_n509), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n512), .B1(new_n513), .B2(new_n511), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n504), .A2(new_n514), .A3(KEYINPUT81), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT81), .B1(new_n504), .B2(new_n514), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT83), .B(G36gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G29gat), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n520));
  NOR3_X1   g319(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT82), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT14), .ZN(new_n524));
  INV_X1    g323(.A(G29gat), .ZN(new_n525));
  INV_X1    g324(.A(G36gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(KEYINPUT82), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n519), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(G43gat), .B(G50gat), .Z(new_n530));
  INV_X1    g329(.A(KEYINPUT15), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT84), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT84), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n529), .A2(new_n535), .A3(new_n532), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n530), .A2(new_n531), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n530), .A2(new_n531), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n537), .A2(new_n519), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n527), .A2(new_n520), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n534), .A2(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT17), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n537), .A2(new_n540), .A3(new_n519), .A4(new_n538), .ZN(new_n543));
  INV_X1    g342(.A(new_n536), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n535), .B1(new_n529), .B2(new_n532), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT86), .ZN(new_n549));
  XNOR2_X1  g348(.A(G15gat), .B(G22gat), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n550), .A2(G1gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT16), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n552), .B2(G1gat), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n549), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n553), .A2(new_n549), .ZN(new_n555));
  NOR3_X1   g354(.A1(new_n554), .A2(new_n555), .A3(G8gat), .ZN(new_n556));
  INV_X1    g355(.A(G8gat), .ZN(new_n557));
  AOI211_X1 g356(.A(KEYINPUT85), .B(new_n557), .C1(new_n551), .C2(new_n553), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT85), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n551), .A2(new_n553), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n559), .B1(new_n560), .B2(G8gat), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n556), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n542), .A2(new_n548), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT87), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(new_n562), .B2(new_n541), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G229gat), .A2(G233gat), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n542), .A2(new_n548), .A3(new_n564), .A4(new_n562), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT18), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n562), .B(new_n541), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n567), .B(KEYINPUT13), .Z(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n566), .A2(KEYINPUT18), .A3(new_n567), .A4(new_n568), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n571), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G113gat), .B(G141gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G197gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT11), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(new_n357), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n580), .B(KEYINPUT12), .Z(new_n581));
  NAND2_X1  g380(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n581), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n583), .A2(new_n571), .A3(new_n574), .A4(new_n575), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(G230gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n587), .A2(new_n468), .ZN(new_n588));
  OR2_X1    g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT88), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(G57gat), .B(G64gat), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(G57gat), .ZN(new_n596));
  OR2_X1    g395(.A1(KEYINPUT89), .A2(G64gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(KEYINPUT89), .A2(G64gat), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT90), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n593), .B1(new_n589), .B2(new_n590), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT90), .B1(new_n352), .B2(G57gat), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n601), .B(new_n602), .C1(new_n599), .C2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n595), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G85gat), .A2(G92gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT7), .ZN(new_n608));
  NAND2_X1  g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  INV_X1    g408(.A(G85gat), .ZN(new_n610));
  AOI22_X1  g409(.A1(KEYINPUT8), .A2(new_n609), .B1(new_n610), .B2(new_n354), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G99gat), .B(G106gat), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n612), .B(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(KEYINPUT93), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n612), .B(new_n613), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT93), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g418(.A(KEYINPUT10), .B(new_n606), .C1(new_n616), .C2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n617), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n615), .A2(new_n604), .A3(new_n595), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT10), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n588), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n621), .A2(new_n622), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n588), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(new_n358), .ZN(new_n631));
  INV_X1    g430(.A(G204gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n633), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n626), .A2(new_n628), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n586), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT21), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n562), .B1(new_n639), .B2(new_n605), .ZN(new_n640));
  XOR2_X1   g439(.A(G127gat), .B(G155gat), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n606), .A2(KEYINPUT21), .ZN(new_n643));
  INV_X1    g442(.A(new_n641), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n562), .B(new_n644), .C1(new_n639), .C2(new_n605), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n643), .B1(new_n642), .B2(new_n645), .ZN(new_n648));
  OAI211_X1 g447(.A(G231gat), .B(G233gat), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n648), .ZN(new_n650));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n651), .A3(new_n646), .ZN(new_n652));
  XNOR2_X1  g451(.A(G183gat), .B(G211gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT20), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n649), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n656), .B1(new_n649), .B2(new_n652), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G232gat), .A2(G233gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT92), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n663), .A2(KEYINPUT41), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(new_n212), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n617), .B(KEYINPUT93), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n542), .A2(new_n667), .A3(new_n548), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n663), .A2(KEYINPUT41), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n546), .B1(new_n619), .B2(new_n616), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(G134gat), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n668), .A2(new_n294), .A3(new_n669), .A4(new_n670), .ZN(new_n673));
  XNOR2_X1  g472(.A(G190gat), .B(G218gat), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n675), .B1(new_n672), .B2(new_n673), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n666), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n678), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n665), .A3(new_n676), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n660), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n517), .A2(new_n638), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n453), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g487(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n552), .A2(new_n557), .ZN(new_n690));
  NOR4_X1   g489(.A1(new_n684), .A2(new_n454), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(KEYINPUT42), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT94), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G8gat), .B1(new_n684), .B2(new_n454), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(KEYINPUT42), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT95), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(G1325gat));
  XNOR2_X1  g497(.A(new_n503), .B(KEYINPUT96), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n685), .A2(G15gat), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n497), .A2(new_n498), .ZN(new_n702));
  AOI21_X1  g501(.A(G15gat), .B1(new_n685), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n701), .A2(new_n703), .ZN(G1326gat));
  OR3_X1    g503(.A1(new_n684), .A2(KEYINPUT97), .A3(new_n285), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT97), .B1(new_n684), .B2(new_n285), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT43), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n705), .A2(new_n709), .A3(new_n706), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(G22gat), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n708), .A2(G22gat), .A3(new_n710), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1327gat));
  INV_X1    g514(.A(new_n682), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n504), .B2(new_n514), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(KEYINPUT44), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n515), .A2(new_n516), .A3(new_n716), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(KEYINPUT44), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n638), .A2(new_n660), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G29gat), .B1(new_n723), .B2(new_n453), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n719), .A2(new_n525), .A3(new_n686), .A4(new_n722), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n725), .A2(KEYINPUT45), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(KEYINPUT45), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n724), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT98), .ZN(G1328gat));
  NAND2_X1  g528(.A1(new_n719), .A2(new_n722), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n730), .A2(new_n518), .A3(new_n454), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT46), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT99), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n518), .B1(new_n723), .B2(new_n454), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n734), .B(new_n735), .C1(new_n732), .C2(new_n731), .ZN(G1329gat));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT100), .ZN(new_n738));
  INV_X1    g537(.A(new_n503), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n720), .A2(new_n738), .A3(new_n739), .A4(new_n722), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n504), .A2(new_n514), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT81), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n504), .A2(new_n514), .A3(KEYINPUT81), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n743), .A2(KEYINPUT44), .A3(new_n744), .A4(new_n682), .ZN(new_n745));
  INV_X1    g544(.A(new_n718), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n745), .A2(new_n746), .A3(new_n739), .A4(new_n722), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT100), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n740), .A2(G43gat), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(G43gat), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n719), .A2(new_n750), .A3(new_n702), .A4(new_n722), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n737), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n751), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n720), .A2(new_n700), .A3(new_n722), .ZN(new_n754));
  AOI211_X1 g553(.A(KEYINPUT47), .B(new_n753), .C1(new_n754), .C2(G43gat), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT101), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(G43gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n757), .A2(new_n737), .A3(new_n751), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT101), .ZN(new_n759));
  AND4_X1   g558(.A1(new_n739), .A2(new_n745), .A3(new_n746), .A4(new_n722), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n750), .B1(new_n760), .B2(new_n738), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n753), .B1(new_n761), .B2(new_n748), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n758), .B(new_n759), .C1(new_n762), .C2(new_n737), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n756), .A2(new_n763), .ZN(G1330gat));
  NOR3_X1   g563(.A1(new_n730), .A2(G50gat), .A3(new_n285), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n720), .A2(new_n451), .A3(new_n722), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(G50gat), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT48), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT102), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n768), .A2(KEYINPUT102), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1331gat));
  NOR3_X1   g571(.A1(new_n660), .A2(new_n585), .A3(new_n682), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n741), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n637), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n453), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(new_n596), .ZN(G1332gat));
  INV_X1    g576(.A(new_n775), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT49), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n431), .B1(new_n779), .B2(new_n352), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT103), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n782), .A2(new_n779), .A3(new_n352), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n778), .B(new_n781), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT104), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT104), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n783), .A2(new_n787), .A3(new_n784), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n786), .A2(KEYINPUT105), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT105), .B1(new_n786), .B2(new_n788), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(G1333gat));
  NAND3_X1  g590(.A1(new_n778), .A2(G71gat), .A3(new_n700), .ZN(new_n792));
  INV_X1    g591(.A(G71gat), .ZN(new_n793));
  INV_X1    g592(.A(new_n702), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n775), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT106), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(G1334gat));
  NAND2_X1  g598(.A1(new_n778), .A2(new_n451), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g600(.A1(new_n659), .A2(new_n585), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n720), .A2(new_n637), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(G85gat), .B1(new_n803), .B2(new_n453), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n717), .A2(new_n802), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n637), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n686), .A2(new_n610), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n804), .B1(new_n808), .B2(new_n809), .ZN(G1336gat));
  INV_X1    g609(.A(new_n808), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n454), .A2(G92gat), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n811), .A2(new_n812), .B1(KEYINPUT108), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G92gat), .B1(new_n803), .B2(new_n454), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n814), .B(new_n815), .C1(KEYINPUT108), .C2(new_n813), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n805), .A2(KEYINPUT107), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n806), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n818), .B(new_n637), .C1(new_n807), .C2(new_n817), .ZN(new_n819));
  INV_X1    g618(.A(new_n812), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n815), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT52), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n816), .A2(new_n822), .ZN(G1337gat));
  OAI21_X1  g622(.A(G99gat), .B1(new_n803), .B2(new_n699), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n702), .A2(new_n476), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n808), .B2(new_n825), .ZN(G1338gat));
  OAI21_X1  g625(.A(G106gat), .B1(new_n803), .B2(new_n285), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n285), .A2(G106gat), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n827), .B1(new_n819), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT53), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n827), .B(new_n831), .C1(new_n808), .C2(new_n828), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1339gat));
  INV_X1    g632(.A(new_n637), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n773), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n567), .B1(new_n566), .B2(new_n568), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n572), .A2(new_n573), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n580), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n584), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(KEYINPUT109), .A3(new_n637), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n620), .A2(new_n588), .A3(new_n624), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT54), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n625), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n620), .A2(new_n624), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846));
  INV_X1    g645(.A(new_n588), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n633), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n841), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n635), .B1(new_n625), .B2(new_n846), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n851), .B(KEYINPUT55), .C1(new_n625), .C2(new_n843), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n852), .A3(new_n636), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n585), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n584), .A2(new_n637), .A3(new_n838), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT109), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n716), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n682), .A2(new_n839), .A3(new_n854), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(KEYINPUT110), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n660), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n861), .B1(new_n859), .B2(new_n716), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(KEYINPUT110), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n835), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n510), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n686), .A2(new_n454), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n298), .B1(new_n870), .B2(new_n585), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT111), .ZN(new_n872));
  INV_X1    g671(.A(new_n870), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n585), .A2(new_n298), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT112), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n872), .B1(new_n873), .B2(new_n875), .ZN(G1340gat));
  NAND2_X1  g675(.A1(new_n870), .A2(new_n637), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n296), .A2(KEYINPUT113), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n296), .A2(KEYINPUT113), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(new_n877), .B2(new_n878), .ZN(G1341gat));
  NAND2_X1  g680(.A1(new_n870), .A2(new_n659), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g682(.A1(new_n870), .A2(new_n682), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(G134gat), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT56), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(G134gat), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1343gat));
  AOI21_X1  g687(.A(KEYINPUT114), .B1(new_n867), .B2(new_n686), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n773), .A2(new_n834), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n659), .B1(new_n865), .B2(KEYINPUT110), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT110), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n856), .A2(new_n857), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n853), .B1(new_n582), .B2(new_n584), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n682), .B1(new_n895), .B2(new_n858), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n892), .B1(new_n896), .B2(new_n861), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n890), .B1(new_n891), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT114), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n898), .A2(new_n899), .A3(new_n453), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n699), .A2(new_n451), .A3(new_n454), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n889), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n216), .A3(new_n585), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n898), .A2(KEYINPUT57), .A3(new_n285), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n855), .A2(new_n856), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n716), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n659), .B1(new_n862), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n890), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT57), .B1(new_n908), .B2(new_n285), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n739), .A2(new_n869), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n904), .A2(new_n911), .A3(new_n586), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n903), .B1(new_n912), .B2(new_n216), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT58), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT58), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n903), .B(new_n915), .C1(new_n216), .C2(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1344gat));
  NAND2_X1  g716(.A1(new_n219), .A2(new_n220), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n918), .A3(new_n637), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT57), .B1(new_n898), .B2(new_n285), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT57), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n835), .A2(KEYINPUT115), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT115), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n773), .A2(new_n924), .A3(new_n834), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n922), .B(new_n451), .C1(new_n926), .C2(new_n907), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n921), .A2(new_n637), .A3(new_n910), .A4(new_n927), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n928), .A2(KEYINPUT116), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n218), .B1(new_n928), .B2(KEYINPUT116), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n920), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n904), .A2(new_n911), .ZN(new_n932));
  AOI211_X1 g731(.A(KEYINPUT59), .B(new_n918), .C1(new_n932), .C2(new_n637), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n919), .B1(new_n931), .B2(new_n933), .ZN(G1345gat));
  AOI21_X1  g733(.A(G155gat), .B1(new_n902), .B2(new_n659), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n660), .A2(new_n211), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n932), .B2(new_n936), .ZN(G1346gat));
  AOI21_X1  g736(.A(G162gat), .B1(new_n902), .B2(new_n682), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n716), .A2(new_n212), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n932), .B2(new_n939), .ZN(G1347gat));
  NOR2_X1   g739(.A1(new_n686), .A2(new_n454), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n867), .A2(new_n510), .A3(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(new_n357), .A3(new_n585), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT117), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n891), .A2(new_n897), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n509), .B1(new_n946), .B2(new_n835), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n945), .B1(new_n947), .B2(new_n941), .ZN(new_n948));
  INV_X1    g747(.A(new_n941), .ZN(new_n949));
  NOR4_X1   g748(.A1(new_n898), .A2(KEYINPUT117), .A3(new_n509), .A4(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n585), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT118), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n951), .A2(new_n952), .A3(G169gat), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n952), .B1(new_n951), .B2(G169gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n944), .B1(new_n953), .B2(new_n954), .ZN(G1348gat));
  AOI21_X1  g754(.A(G176gat), .B1(new_n943), .B2(new_n637), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n942), .A2(KEYINPUT117), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n947), .A2(new_n945), .A3(new_n941), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n834), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n956), .B1(new_n959), .B2(G176gat), .ZN(G1349gat));
  NAND3_X1  g759(.A1(new_n943), .A2(new_n372), .A3(new_n659), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n660), .B1(new_n957), .B2(new_n958), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(new_n399), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n716), .B1(new_n957), .B2(new_n958), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n966), .A2(KEYINPUT120), .A3(new_n373), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT120), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n682), .B1(new_n948), .B2(new_n950), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(G190gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n965), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(KEYINPUT120), .B1(new_n966), .B2(new_n373), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n969), .A2(new_n968), .A3(G190gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n972), .A2(new_n973), .A3(KEYINPUT61), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n943), .A2(new_n373), .A3(new_n682), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT119), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n971), .A2(new_n974), .A3(new_n976), .ZN(G1351gat));
  NAND2_X1  g776(.A1(new_n699), .A2(new_n941), .ZN(new_n978));
  XOR2_X1   g777(.A(new_n978), .B(KEYINPUT123), .Z(new_n979));
  INV_X1    g778(.A(KEYINPUT122), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n921), .A2(new_n980), .A3(new_n927), .ZN(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n980), .B1(new_n921), .B2(new_n927), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n585), .B(new_n979), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(KEYINPUT124), .ZN(new_n985));
  INV_X1    g784(.A(new_n927), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n922), .B1(new_n867), .B2(new_n451), .ZN(new_n987));
  OAI21_X1  g786(.A(KEYINPUT122), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(new_n981), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT124), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n989), .A2(new_n990), .A3(new_n585), .A4(new_n979), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n985), .A2(G197gat), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n699), .A2(new_n451), .A3(new_n431), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n993), .A2(KEYINPUT121), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n686), .B1(new_n993), .B2(KEYINPUT121), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n867), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  OR3_X1    g795(.A1(new_n996), .A2(G197gat), .A3(new_n586), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n992), .A2(new_n997), .ZN(G1352gat));
  INV_X1    g797(.A(new_n996), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n999), .A2(new_n632), .A3(new_n637), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT125), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g801(.A1(new_n999), .A2(KEYINPUT125), .A3(new_n632), .A4(new_n637), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n1004));
  OAI211_X1 g803(.A(new_n1002), .B(new_n1003), .C1(KEYINPUT126), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(KEYINPUT126), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n989), .A2(new_n637), .A3(new_n979), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(G204gat), .ZN(new_n1009));
  NAND4_X1  g808(.A1(new_n1002), .A2(KEYINPUT126), .A3(new_n1004), .A4(new_n1003), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(G1353gat));
  NAND3_X1  g810(.A1(new_n999), .A2(new_n237), .A3(new_n659), .ZN(new_n1012));
  OR4_X1    g811(.A1(new_n660), .A2(new_n986), .A3(new_n987), .A4(new_n978), .ZN(new_n1013));
  AND3_X1   g812(.A1(new_n1013), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1014));
  AOI21_X1  g813(.A(KEYINPUT63), .B1(new_n1013), .B2(G211gat), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(G1354gat));
  OAI21_X1  g815(.A(new_n238), .B1(new_n996), .B2(new_n716), .ZN(new_n1017));
  XOR2_X1   g816(.A(new_n1017), .B(KEYINPUT127), .Z(new_n1018));
  AND2_X1   g817(.A1(new_n989), .A2(new_n979), .ZN(new_n1019));
  NOR2_X1   g818(.A1(new_n716), .A2(new_n238), .ZN(new_n1020));
  AOI21_X1  g819(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(G1355gat));
endmodule


