//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1258, new_n1259, new_n1260,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT65), .Z(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  INV_X1    g0015(.A(G97), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  AND3_X1   g0026(.A1(KEYINPUT66), .A2(G1), .A3(G13), .ZN(new_n227));
  AOI21_X1  g0027(.A(KEYINPUT66), .B1(G1), .B2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n207), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n212), .A2(new_n226), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XOR2_X1   g0038(.A(G226), .B(G232), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n240), .B(new_n244), .Z(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT69), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  OAI21_X1  g0053(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT70), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G274), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  AOI21_X1  g0063(.A(G1), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT71), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n254), .A2(KEYINPUT71), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n258), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n261), .B1(G226), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G33), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G223), .A3(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G222), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n276), .B1(new_n222), .B2(new_n275), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G1), .A2(G13), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT66), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(KEYINPUT66), .A2(G1), .A3(G13), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n257), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n270), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G200), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n270), .A2(new_n288), .A3(G190), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT75), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT10), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n283), .A2(new_n284), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT72), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G58), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT8), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n271), .A2(G20), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n300), .A2(new_n301), .B1(G150), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n202), .A2(G20), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n297), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n220), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n296), .B1(new_n206), .B2(G20), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(new_n220), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n306), .A2(KEYINPUT9), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT9), .ZN(new_n312));
  INV_X1    g0112(.A(new_n310), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n305), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n292), .A2(new_n293), .A3(new_n294), .A4(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n290), .A2(new_n311), .A3(new_n291), .A4(new_n314), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT75), .B1(new_n317), .B2(KEYINPUT10), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(KEYINPUT10), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G179), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n289), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(G169), .B2(new_n289), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n306), .A2(new_n310), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n261), .B1(G244), .B2(new_n269), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n275), .A2(G232), .A3(new_n277), .ZN(new_n330));
  INV_X1    g0130(.A(G107), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(new_n275), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n272), .A2(new_n274), .ZN(new_n333));
  INV_X1    g0133(.A(G238), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n333), .A2(new_n334), .A3(new_n277), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n287), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G200), .ZN(new_n338));
  INV_X1    g0138(.A(G190), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT8), .B(G58), .ZN(new_n340));
  INV_X1    g0140(.A(new_n302), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n340), .A2(new_n341), .B1(new_n207), .B2(new_n222), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT15), .B(G87), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n342), .A2(KEYINPUT73), .B1(new_n301), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(KEYINPUT73), .B2(new_n342), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n296), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n307), .A2(new_n222), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n309), .B2(new_n222), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n338), .B1(new_n339), .B2(new_n337), .C1(new_n351), .C2(KEYINPUT74), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n351), .A2(KEYINPUT74), .ZN(new_n353));
  OR2_X1    g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n329), .A2(G179), .A3(new_n336), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n337), .A2(G169), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n351), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n321), .A2(new_n328), .A3(new_n354), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n301), .A2(G77), .ZN(new_n360));
  INV_X1    g0160(.A(G68), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G20), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n360), .B(new_n362), .C1(new_n220), .C2(new_n341), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n296), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT11), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n206), .A2(G13), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  XOR2_X1   g0167(.A(new_n367), .B(KEYINPUT12), .Z(new_n368));
  INV_X1    g0168(.A(new_n309), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n365), .B(new_n368), .C1(new_n361), .C2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n268), .A2(new_n334), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT76), .B1(new_n371), .B2(new_n261), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n256), .A2(new_n260), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT76), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n373), .B(new_n374), .C1(new_n334), .C2(new_n268), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n275), .A2(G232), .A3(G1698), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G97), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n376), .B(new_n377), .C1(new_n278), .C2(new_n221), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n287), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n372), .A2(new_n375), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT13), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT13), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n372), .A2(new_n382), .A3(new_n375), .A4(new_n379), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(G179), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G169), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(new_n381), .B2(new_n383), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT14), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n384), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI211_X1 g0188(.A(KEYINPUT14), .B(new_n385), .C1(new_n381), .C2(new_n383), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n370), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n381), .A2(G190), .A3(new_n383), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT77), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT77), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n381), .A2(new_n393), .A3(G190), .A4(new_n383), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n381), .A2(new_n383), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n370), .B1(new_n396), .B2(G200), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n390), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g0199(.A(G58), .B(G68), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n400), .A2(G20), .B1(G159), .B2(new_n302), .ZN(new_n401));
  INV_X1    g0201(.A(new_n272), .ZN(new_n402));
  XNOR2_X1  g0202(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n402), .B1(new_n403), .B2(G33), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n404), .A2(G20), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT7), .ZN(new_n406));
  OAI21_X1  g0206(.A(G68), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n273), .A2(KEYINPUT78), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT78), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT3), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n410), .A3(G33), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n272), .ZN(new_n412));
  XOR2_X1   g0212(.A(KEYINPUT79), .B(KEYINPUT7), .Z(new_n413));
  AND3_X1   g0213(.A1(new_n412), .A2(new_n207), .A3(new_n413), .ZN(new_n414));
  OAI211_X1 g0214(.A(KEYINPUT16), .B(new_n401), .C1(new_n407), .C2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT16), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n274), .B1(new_n403), .B2(G33), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n413), .B1(new_n275), .B2(G20), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n361), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n401), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n416), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n415), .A2(new_n296), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n300), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n307), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n309), .B2(new_n424), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g0227(.A(G232), .B(new_n258), .C1(new_n266), .C2(new_n267), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n373), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n277), .A2(G223), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n221), .B2(new_n277), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n411), .A2(new_n431), .A3(new_n272), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G33), .A2(G87), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n286), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT80), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n432), .A2(new_n433), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n287), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT80), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n437), .A2(new_n438), .A3(new_n373), .A4(new_n428), .ZN(new_n439));
  AOI21_X1  g0239(.A(G169), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n429), .A2(G179), .A3(new_n434), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n427), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT18), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n423), .A2(new_n426), .ZN(new_n445));
  AOI21_X1  g0245(.A(G200), .B1(new_n435), .B2(new_n439), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n429), .A2(G190), .A3(new_n434), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n445), .A2(new_n448), .A3(KEYINPUT17), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n423), .B(new_n426), .C1(new_n446), .C2(new_n447), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT18), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n427), .A2(new_n442), .A3(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n444), .A2(new_n449), .A3(new_n452), .A4(new_n454), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n359), .A2(new_n399), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n331), .B1(new_n418), .B2(new_n419), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT6), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n216), .A2(new_n331), .ZN(new_n459));
  NOR2_X1   g0259(.A1(G97), .A2(G107), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n331), .A2(KEYINPUT6), .A3(G97), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI22_X1  g0263(.A1(new_n463), .A2(new_n207), .B1(new_n222), .B2(new_n341), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n296), .B1(new_n457), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n307), .A2(new_n216), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n206), .A2(G33), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n307), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n296), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n466), .B1(new_n469), .B2(new_n216), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n223), .A2(G1698), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT4), .B1(new_n404), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n272), .A2(new_n274), .A3(G250), .A4(G1698), .ZN(new_n473));
  AND2_X1   g0273(.A1(KEYINPUT4), .A2(G244), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n272), .A2(new_n274), .A3(new_n474), .A4(new_n277), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n287), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n206), .B(G45), .C1(new_n262), .C2(KEYINPUT5), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT5), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G41), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n258), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT82), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n480), .B2(G41), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n262), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n263), .A2(G1), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n480), .A2(G41), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n482), .A2(new_n217), .B1(new_n488), .B2(new_n259), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n478), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n465), .B(new_n470), .C1(new_n491), .C2(new_n339), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n411), .A2(new_n272), .A3(new_n471), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n286), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n490), .B1(new_n497), .B2(KEYINPUT81), .ZN(new_n498));
  OAI211_X1 g0298(.A(KEYINPUT81), .B(new_n287), .C1(new_n472), .C2(new_n477), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(G200), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT83), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(KEYINPUT83), .B(G200), .C1(new_n498), .C2(new_n500), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n492), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(G264), .B(new_n258), .C1(new_n479), .C2(new_n481), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  MUX2_X1   g0307(.A(new_n215), .B(new_n217), .S(G1698), .Z(new_n508));
  INV_X1    g0308(.A(G294), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n412), .A2(new_n508), .B1(new_n271), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n507), .B1(new_n510), .B2(new_n287), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n488), .A2(new_n259), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(G200), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(G190), .B2(new_n513), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n366), .A2(new_n207), .A3(G107), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(KEYINPUT93), .A3(KEYINPUT25), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(KEYINPUT25), .B2(new_n517), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT93), .B1(new_n517), .B2(KEYINPUT25), .ZN(new_n520));
  OR2_X1    g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n469), .A2(G107), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n404), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT22), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n207), .A2(G87), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n333), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(G116), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT84), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT84), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G116), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n301), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT92), .B1(new_n331), .B2(G20), .ZN(new_n534));
  XOR2_X1   g0334(.A(new_n534), .B(KEYINPUT23), .Z(new_n535));
  NAND4_X1  g0335(.A1(new_n524), .A2(new_n527), .A3(new_n533), .A4(new_n535), .ZN(new_n536));
  XNOR2_X1  g0336(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n537));
  OR2_X1    g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n297), .B1(new_n536), .B2(new_n537), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n523), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n516), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n465), .A2(new_n470), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT81), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n477), .B1(new_n494), .B2(new_n493), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n543), .B1(new_n544), .B2(new_n286), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n545), .A2(new_n322), .A3(new_n490), .A4(new_n499), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n491), .A2(new_n385), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n542), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n505), .A2(new_n541), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n307), .A2(new_n467), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n551), .A2(G116), .A3(new_n229), .A4(new_n295), .ZN(new_n552));
  XNOR2_X1  g0352(.A(KEYINPUT84), .B(G116), .ZN(new_n553));
  INV_X1    g0353(.A(new_n307), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n207), .B1(new_n529), .B2(new_n531), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n271), .A2(G97), .ZN(new_n558));
  AOI21_X1  g0358(.A(G20), .B1(new_n558), .B2(new_n476), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n296), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT20), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(KEYINPUT20), .B(new_n296), .C1(new_n557), .C2(new_n559), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n556), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(G270), .ZN(new_n565));
  OAI22_X1  g0365(.A1(new_n482), .A2(new_n565), .B1(new_n488), .B2(new_n259), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G264), .A2(G1698), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n217), .B2(G1698), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n411), .A2(new_n272), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(G303), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT87), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT87), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G303), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n333), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n287), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n567), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(G190), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n286), .B1(new_n570), .B2(new_n576), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n581), .A2(new_n566), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n582), .A2(G200), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n564), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g0384(.A(new_n584), .B(KEYINPUT89), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(G179), .ZN(new_n586));
  OAI211_X1 g0386(.A(KEYINPUT21), .B(G169), .C1(new_n581), .C2(new_n566), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n564), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT88), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n469), .A2(G116), .B1(new_n554), .B2(new_n553), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n476), .B1(new_n216), .B2(G33), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n207), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n207), .B2(new_n553), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT20), .B1(new_n594), .B2(new_n296), .ZN(new_n595));
  INV_X1    g0395(.A(new_n563), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(G169), .A3(new_n579), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT21), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n590), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(G169), .B1(new_n581), .B2(new_n566), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n590), .B(new_n599), .C1(new_n564), .C2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n589), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT90), .B1(new_n585), .B2(new_n604), .ZN(new_n605));
  OR2_X1    g0405(.A1(new_n584), .A2(KEYINPUT89), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n599), .B1(new_n564), .B2(new_n601), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT88), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n588), .B1(new_n608), .B2(new_n602), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT90), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n584), .A2(KEYINPUT89), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n606), .A2(new_n609), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n513), .A2(G169), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n511), .A2(G179), .A3(new_n512), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n540), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT19), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n207), .B1(new_n377), .B2(new_n618), .ZN(new_n619));
  NOR4_X1   g0419(.A1(KEYINPUT85), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT85), .ZN(new_n621));
  NOR2_X1   g0421(.A1(G87), .A2(G97), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(new_n331), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n619), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n411), .A2(new_n207), .A3(G68), .A4(new_n272), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n618), .B1(new_n377), .B2(G20), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n296), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n469), .A2(new_n344), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT86), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n343), .A2(new_n554), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT86), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n469), .A2(new_n632), .A3(new_n344), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n628), .A2(new_n630), .A3(new_n631), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(G244), .A2(G1698), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n334), .B2(G1698), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n411), .A2(new_n272), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n532), .A2(G33), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n286), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n486), .A2(G274), .ZN(new_n640));
  OAI21_X1  g0440(.A(G250), .B1(new_n263), .B2(G1), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n258), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n385), .B1(new_n639), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n639), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n322), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n634), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(G190), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n627), .A2(new_n296), .B1(new_n554), .B2(new_n343), .ZN(new_n650));
  OAI21_X1  g0450(.A(G200), .B1(new_n639), .B2(new_n644), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n469), .A2(G87), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n649), .A2(new_n650), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n617), .A2(new_n654), .ZN(new_n655));
  AND4_X1   g0455(.A1(new_n456), .A2(new_n550), .A3(new_n613), .A4(new_n655), .ZN(G372));
  INV_X1    g0456(.A(new_n398), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n390), .B1(new_n657), .B2(new_n358), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n449), .A2(new_n452), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n454), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n453), .B1(new_n427), .B2(new_n442), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n327), .B1(new_n664), .B2(new_n321), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT98), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n546), .A2(new_n666), .A3(new_n547), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n666), .B1(new_n546), .B2(new_n547), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT94), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n643), .B1(new_n639), .B2(new_n670), .ZN(new_n671));
  AOI211_X1 g0471(.A(KEYINPUT94), .B(new_n286), .C1(new_n638), .C2(new_n637), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n385), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT95), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n630), .A2(new_n633), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n675), .A2(new_n650), .B1(new_n322), .B2(new_n646), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT95), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n677), .B(new_n385), .C1(new_n671), .C2(new_n672), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n674), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n650), .A2(new_n652), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n671), .A2(new_n672), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n680), .B(new_n649), .C1(new_n681), .C2(new_n514), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT26), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n669), .A2(new_n683), .A3(new_n684), .A4(new_n542), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT26), .B1(new_n548), .B2(new_n654), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT97), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n679), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n674), .A2(new_n676), .A3(KEYINPUT97), .A4(new_n678), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT96), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n604), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n609), .A2(KEYINPUT96), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n617), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n492), .ZN(new_n696));
  INV_X1    g0496(.A(new_n504), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n545), .A2(new_n490), .A3(new_n499), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT83), .B1(new_n698), .B2(G200), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n696), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n516), .A2(new_n540), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n683), .A2(new_n700), .A3(new_n701), .A4(new_n548), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n685), .B(new_n691), .C1(new_n695), .C2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n456), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n665), .A2(new_n704), .ZN(G369));
  OR3_X1    g0505(.A1(new_n366), .A2(KEYINPUT27), .A3(G20), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT27), .B1(new_n366), .B2(G20), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G213), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G343), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n605), .B(new_n612), .C1(new_n564), .C2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n608), .A2(new_n602), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT96), .B1(new_n713), .B2(new_n589), .ZN(new_n714));
  AOI211_X1 g0514(.A(new_n692), .B(new_n588), .C1(new_n608), .C2(new_n602), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n597), .B(new_n710), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n712), .A2(G330), .A3(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n701), .B1(new_n540), .B2(new_n711), .ZN(new_n719));
  INV_X1    g0519(.A(new_n617), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n617), .A2(new_n711), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n609), .A2(new_n710), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n721), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n722), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT99), .ZN(G399));
  INV_X1    g0530(.A(KEYINPUT100), .ZN(new_n731));
  INV_X1    g0531(.A(new_n210), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n731), .B1(new_n732), .B2(G41), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n210), .A2(KEYINPUT100), .A3(new_n262), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n206), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n620), .A2(new_n623), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n528), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n737), .A2(new_n740), .B1(new_n232), .B2(new_n736), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT28), .Z(new_n742));
  INV_X1    g0542(.A(G330), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT102), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  AOI21_X1  g0545(.A(KEYINPUT101), .B1(new_n582), .B2(G179), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT101), .ZN(new_n747));
  NOR4_X1   g0547(.A1(new_n581), .A2(new_n566), .A3(new_n747), .A4(new_n322), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n478), .A2(new_n511), .A3(new_n646), .A4(new_n490), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n745), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AND4_X1   g0551(.A1(new_n511), .A2(new_n478), .A3(new_n646), .A4(new_n490), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n752), .B(KEYINPUT30), .C1(new_n746), .C2(new_n748), .ZN(new_n753));
  INV_X1    g0553(.A(new_n681), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n582), .A2(G179), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n754), .A2(new_n698), .A3(new_n513), .A4(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n751), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n757), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n758));
  AOI21_X1  g0558(.A(KEYINPUT31), .B1(new_n757), .B2(new_n710), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n744), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n757), .A2(new_n710), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT31), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n757), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n763), .A2(KEYINPUT102), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n613), .A2(new_n550), .A3(new_n655), .A4(new_n711), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n743), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n703), .A2(new_n711), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT29), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n688), .A2(new_n689), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT103), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n542), .B1(new_n667), .B2(new_n668), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n679), .A2(new_n682), .ZN(new_n775));
  OAI21_X1  g0575(.A(KEYINPUT26), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n772), .A2(KEYINPUT103), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n549), .A2(new_n684), .A3(new_n648), .A4(new_n653), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n773), .A2(new_n776), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n702), .B1(new_n609), .B2(new_n720), .ZN(new_n780));
  OAI211_X1 g0580(.A(KEYINPUT29), .B(new_n711), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n768), .B1(new_n771), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n742), .B1(new_n782), .B2(G1), .ZN(G364));
  AOI21_X1  g0583(.A(new_n229), .B1(G20), .B2(new_n385), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n207), .A2(new_n339), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(G179), .A3(new_n514), .ZN(new_n786));
  INV_X1    g0586(.A(G58), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n339), .A2(G179), .A3(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n207), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n275), .B1(new_n786), .B2(new_n787), .C1(new_n216), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n322), .A2(new_n514), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n785), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n207), .A2(G190), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G50), .A2(new_n793), .B1(new_n796), .B2(G68), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n514), .A2(G179), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n794), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n800), .A2(new_n322), .A3(G200), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n797), .B1(new_n331), .B2(new_n799), .C1(new_n222), .C2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n785), .A2(new_n798), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n804), .A2(KEYINPUT105), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(KEYINPUT105), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n790), .B(new_n803), .C1(G87), .C2(new_n808), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n800), .A2(G179), .A3(G200), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n810), .A2(KEYINPUT104), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(KEYINPUT104), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(G159), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT32), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n809), .A2(new_n816), .A3(KEYINPUT106), .ZN(new_n817));
  INV_X1    g0617(.A(new_n813), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n818), .A2(G329), .B1(G303), .B2(new_n808), .ZN(new_n819));
  INV_X1    g0619(.A(G311), .ZN(new_n820));
  INV_X1    g0620(.A(G326), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n802), .A2(new_n820), .B1(new_n821), .B2(new_n792), .ZN(new_n822));
  INV_X1    g0622(.A(G322), .ZN(new_n823));
  XOR2_X1   g0623(.A(KEYINPUT33), .B(G317), .Z(new_n824));
  OAI22_X1  g0624(.A1(new_n823), .A2(new_n786), .B1(new_n824), .B2(new_n795), .ZN(new_n825));
  INV_X1    g0625(.A(G283), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n333), .B1(new_n799), .B2(new_n826), .C1(new_n789), .C2(new_n509), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n822), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n819), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n817), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(KEYINPUT106), .B1(new_n809), .B2(new_n816), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n784), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G13), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(G20), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(G45), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n737), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n732), .A2(new_n333), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n837), .A2(G355), .B1(new_n528), .B2(new_n732), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n232), .A2(G45), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n252), .B2(G45), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n732), .A2(new_n404), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n838), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(G13), .A2(G33), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(G20), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n784), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n836), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n832), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n712), .A2(new_n716), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n850), .B2(new_n846), .ZN(new_n851));
  INV_X1    g0651(.A(new_n836), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n718), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n850), .A2(new_n743), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G396));
  INV_X1    g0656(.A(new_n786), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n857), .A2(G143), .B1(new_n796), .B2(G150), .ZN(new_n858));
  INV_X1    g0658(.A(G137), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n858), .B1(new_n859), .B2(new_n792), .C1(new_n814), .C2(new_n802), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT34), .Z(new_n861));
  OAI221_X1 g0661(.A(new_n404), .B1(new_n361), .B2(new_n799), .C1(new_n787), .C2(new_n789), .ZN(new_n862));
  INV_X1    g0662(.A(G132), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n813), .A2(new_n863), .B1(new_n220), .B2(new_n807), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n813), .A2(new_n820), .B1(new_n331), .B2(new_n807), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n786), .A2(new_n509), .B1(new_n799), .B2(new_n214), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n802), .A2(new_n553), .B1(new_n571), .B2(new_n792), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n333), .B1(new_n795), .B2(new_n826), .C1(new_n789), .C2(new_n216), .ZN(new_n869));
  NOR4_X1   g0669(.A1(new_n866), .A2(new_n867), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n784), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n784), .A2(new_n844), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n836), .B1(new_n222), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n358), .A2(new_n710), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n352), .A2(new_n353), .B1(new_n351), .B2(new_n711), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n874), .B1(new_n875), .B2(new_n358), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n871), .B(new_n873), .C1(new_n876), .C2(new_n845), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n720), .B1(new_n714), .B2(new_n715), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n878), .A2(new_n550), .A3(new_n683), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n774), .A2(new_n775), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n690), .B1(new_n880), .B2(new_n684), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n710), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT107), .B1(new_n882), .B2(new_n876), .ZN(new_n883));
  AND4_X1   g0683(.A1(KEYINPUT107), .A2(new_n703), .A3(new_n711), .A4(new_n876), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n883), .A2(new_n884), .B1(new_n882), .B2(new_n876), .ZN(new_n885));
  INV_X1    g0685(.A(new_n768), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n836), .B1(new_n885), .B2(new_n886), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n877), .B1(new_n888), .B2(new_n889), .ZN(G384));
  INV_X1    g0690(.A(KEYINPUT35), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n463), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n463), .A2(new_n891), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n892), .A2(G116), .A3(new_n230), .A4(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n895), .A2(KEYINPUT36), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(KEYINPUT36), .ZN(new_n897));
  OAI21_X1  g0697(.A(G77), .B1(new_n787), .B2(new_n361), .ZN(new_n898));
  OAI22_X1  g0698(.A1(new_n898), .A2(new_n231), .B1(G50), .B2(new_n361), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(G1), .A3(new_n833), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n896), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT108), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n399), .A2(new_n370), .A3(new_n710), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n370), .A2(new_n710), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n390), .A2(new_n398), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n758), .A2(new_n759), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n767), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n906), .A2(new_n908), .A3(new_n876), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n415), .A2(new_n296), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n405), .A2(new_n413), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(G68), .C1(new_n406), .C2(new_n405), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT16), .B1(new_n912), .B2(new_n401), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n426), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n708), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n455), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n427), .A2(new_n915), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT37), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n443), .A2(new_n919), .A3(new_n920), .A4(new_n450), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n708), .B1(new_n440), .B2(new_n441), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n445), .A2(new_n448), .B1(new_n914), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n921), .B1(new_n923), .B2(new_n920), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n918), .A2(KEYINPUT38), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n919), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n443), .A2(new_n919), .A3(new_n450), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT37), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n455), .A2(new_n926), .B1(new_n928), .B2(new_n921), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n925), .B1(new_n929), .B2(KEYINPUT38), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT40), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n909), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n918), .A2(KEYINPUT38), .A3(new_n924), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT38), .B1(new_n918), .B2(new_n924), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n933), .B1(new_n909), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n456), .A2(new_n908), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n938), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(G330), .ZN(new_n941));
  INV_X1    g0741(.A(new_n874), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n883), .B2(new_n884), .ZN(new_n943));
  INV_X1    g0743(.A(new_n936), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(new_n906), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n663), .A2(new_n915), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT39), .B1(new_n934), .B2(new_n935), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT39), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n925), .B(new_n948), .C1(new_n929), .C2(KEYINPUT38), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n370), .B(new_n711), .C1(new_n388), .C2(new_n389), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT109), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n946), .B1(new_n950), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n945), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n771), .A2(new_n456), .A3(new_n781), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n665), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n956), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n941), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n206), .B2(new_n834), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n941), .A2(new_n959), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n902), .B1(new_n961), .B2(new_n962), .ZN(G367));
  NAND3_X1  g0763(.A1(new_n669), .A2(new_n542), .A3(new_n710), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n542), .A2(new_n710), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n700), .A2(new_n548), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NOR4_X1   g0767(.A1(new_n719), .A2(new_n609), .A3(new_n617), .A4(new_n710), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT42), .Z(new_n970));
  AOI21_X1  g0770(.A(new_n549), .B1(new_n967), .B2(new_n617), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n970), .B1(new_n710), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n772), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n680), .A2(new_n711), .ZN(new_n974));
  MUX2_X1   g0774(.A(new_n775), .B(new_n973), .S(new_n974), .Z(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT110), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT43), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n972), .B(new_n978), .C1(new_n977), .C2(new_n975), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n972), .B2(new_n978), .ZN(new_n980));
  INV_X1    g0780(.A(new_n967), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n724), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n980), .B(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n735), .B(KEYINPUT41), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n728), .A2(new_n967), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT45), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n985), .B(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n727), .A2(new_n981), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT44), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n988), .B(new_n989), .ZN(new_n990));
  AND3_X1   g0790(.A1(new_n987), .A2(new_n724), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n724), .B1(new_n987), .B2(new_n990), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT112), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n717), .A2(new_n726), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT111), .B1(new_n723), .B2(new_n725), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n712), .A2(G330), .A3(new_n716), .A4(new_n968), .ZN(new_n997));
  AND3_X1   g0797(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n996), .B1(new_n995), .B2(new_n997), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n782), .B(new_n994), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n998), .A2(new_n999), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n782), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT112), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n993), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n984), .B1(new_n1004), .B2(new_n782), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n835), .A2(G1), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n983), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n784), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n799), .A2(new_n216), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n575), .B2(new_n857), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n826), .B2(new_n802), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(new_n818), .B2(G317), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n792), .A2(new_n820), .B1(new_n795), .B2(new_n509), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n789), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n404), .B(new_n1013), .C1(G107), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT46), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n808), .B2(G116), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n807), .A2(KEYINPUT46), .A3(new_n553), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1012), .B(new_n1015), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n275), .B1(new_n799), .B2(new_n222), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT113), .Z(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n787), .B2(new_n807), .C1(new_n859), .C2(new_n813), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n857), .A2(G150), .B1(new_n793), .B2(G143), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n801), .A2(G50), .B1(new_n796), .B2(G159), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(new_n361), .C2(new_n789), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1019), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT114), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT47), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1008), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n975), .A2(new_n846), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n244), .A2(new_n841), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n846), .B(new_n784), .C1(new_n732), .C2(new_n344), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n836), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1030), .A2(new_n1031), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1007), .A2(new_n1035), .ZN(G387));
  NAND2_X1  g0836(.A1(new_n1003), .A2(new_n1000), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n735), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n837), .A2(new_n739), .B1(new_n331), .B2(new_n732), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n740), .B(new_n263), .C1(new_n361), .C2(new_n222), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT50), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n340), .A2(G50), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT115), .Z(new_n1044));
  AOI21_X1  g0844(.A(new_n1041), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n841), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n240), .A2(new_n263), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1040), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n836), .B1(new_n1049), .B2(new_n847), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n846), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1014), .A2(new_n344), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1052), .B(new_n404), .C1(new_n424), .C2(new_n795), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1009), .B1(G159), .B2(new_n793), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n801), .A2(G68), .B1(new_n857), .B2(G50), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n807), .C2(new_n222), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1053), .B(new_n1056), .C1(G150), .C2(new_n818), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n792), .A2(new_n823), .B1(new_n795), .B2(new_n820), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT116), .Z(new_n1059));
  INV_X1    g0859(.A(new_n575), .ZN(new_n1060));
  INV_X1    g0860(.A(G317), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n802), .A2(new_n1060), .B1(new_n1061), .B2(new_n786), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(KEYINPUT48), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n826), .B2(new_n789), .C1(new_n509), .C2(new_n807), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1063), .A2(KEYINPUT48), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(KEYINPUT49), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n412), .B1(new_n553), .B2(new_n799), .C1(new_n813), .C2(new_n821), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n1067), .B2(KEYINPUT49), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1057), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1050), .B1(new_n723), .B2(new_n1051), .C1(new_n1071), .C2(new_n1008), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1006), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1039), .B(new_n1072), .C1(new_n1001), .C2(new_n1073), .ZN(G393));
  NAND2_X1  g0874(.A1(new_n981), .A2(new_n846), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n249), .A2(new_n842), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n847), .B1(new_n216), .B2(new_n210), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n852), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n333), .B1(new_n799), .B2(new_n331), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n802), .A2(new_n509), .B1(new_n1060), .B2(new_n795), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(new_n532), .C2(new_n1014), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n818), .A2(G322), .B1(G283), .B2(new_n808), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n786), .A2(new_n820), .B1(new_n792), .B2(new_n1061), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT52), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n799), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n412), .B1(G87), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n807), .B2(new_n361), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G143), .B2(new_n818), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT117), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n857), .A2(G159), .B1(new_n793), .B2(G150), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n789), .A2(new_n222), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n802), .A2(new_n340), .B1(new_n220), .B2(new_n795), .ZN(new_n1094));
  OR3_X1    g0894(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1085), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1078), .B1(new_n1096), .B2(new_n784), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n993), .A2(new_n1006), .B1(new_n1075), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1004), .A2(new_n736), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n993), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(G390));
  NAND2_X1  g0901(.A1(new_n930), .A2(new_n953), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n875), .A2(new_n358), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n711), .B(new_n1103), .C1(new_n779), .C2(new_n780), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n942), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1102), .B1(new_n1105), .B2(new_n906), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n768), .A2(new_n876), .A3(new_n906), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n954), .B1(new_n943), .B2(new_n906), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1107), .B(new_n1108), .C1(new_n1109), .C2(new_n950), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n703), .A2(new_n711), .A3(new_n876), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT107), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n882), .A2(KEYINPUT107), .A3(new_n876), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n874), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n906), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n953), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n950), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1106), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n876), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(new_n743), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n908), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1122), .A2(new_n1116), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1110), .B(new_n1006), .C1(new_n1119), .C2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n872), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n852), .B1(new_n300), .B2(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n802), .A2(new_n216), .B1(new_n826), .B2(new_n792), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n786), .A2(new_n528), .B1(new_n795), .B2(new_n331), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n275), .B(new_n1093), .C1(G68), .C2(new_n1086), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1132), .B1(new_n214), .B2(new_n807), .C1(new_n509), .C2(new_n813), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT54), .B(G143), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n802), .A2(new_n1134), .B1(new_n859), .B2(new_n795), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT118), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n818), .A2(G125), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n275), .B1(new_n786), .B2(new_n863), .ZN(new_n1138));
  INV_X1    g0938(.A(G128), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n792), .A2(new_n1139), .B1(new_n799), .B2(new_n220), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1138), .B(new_n1140), .C1(G159), .C2(new_n1014), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1137), .B(new_n1141), .C1(new_n1136), .C2(new_n1135), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n808), .A2(G150), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT53), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1133), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1127), .B1(new_n1145), .B2(new_n784), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n950), .B2(new_n845), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1125), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(KEYINPUT119), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n456), .A2(G330), .A3(new_n908), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n665), .A2(new_n957), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n906), .B1(new_n768), .B2(new_n876), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n943), .B1(new_n1123), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1122), .A2(new_n1116), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1154), .A2(new_n1108), .A3(new_n942), .A4(new_n1104), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1151), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1124), .B1(new_n1158), .B2(new_n1107), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1108), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1106), .B(new_n1160), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1157), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1110), .B(new_n1156), .C1(new_n1119), .C2(new_n1124), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n736), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT119), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1125), .A2(new_n1165), .A3(new_n1147), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1149), .A2(new_n1164), .A3(new_n1166), .ZN(G378));
  INV_X1    g0967(.A(new_n1151), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1163), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n932), .A2(new_n937), .A3(G330), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n321), .A2(KEYINPUT120), .A3(new_n328), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT120), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n316), .A2(new_n318), .B1(KEYINPUT10), .B2(new_n317), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1174), .B1(new_n1175), .B2(new_n327), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n326), .A2(new_n708), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1173), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1177), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT121), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n1179), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1177), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1182), .B1(new_n1187), .B2(new_n1178), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1184), .A2(new_n1188), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n945), .A2(new_n955), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(new_n945), .B2(new_n955), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1172), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1189), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1115), .A2(new_n1116), .A3(new_n936), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n949), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n918), .A2(new_n924), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT38), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n948), .B1(new_n1198), .B2(new_n925), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n954), .B1(new_n1195), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n946), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1193), .B1(new_n1194), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n945), .A2(new_n1189), .A3(new_n955), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1203), .A2(new_n1171), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1192), .A2(new_n1205), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1169), .A2(new_n1170), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1170), .B1(new_n1169), .B2(new_n1206), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n736), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n404), .A2(G41), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n807), .B2(new_n222), .C1(new_n813), .C2(new_n826), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n789), .A2(new_n361), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G116), .A2(new_n793), .B1(new_n796), .B2(G97), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n331), .B2(new_n786), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1086), .A2(G58), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n802), .B2(new_n343), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1211), .A2(new_n1212), .A3(new_n1214), .A4(new_n1216), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G50), .B(new_n1210), .C1(new_n271), .C2(new_n262), .ZN(new_n1218));
  OAI21_X1  g1018(.A(KEYINPUT58), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(G125), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n786), .A2(new_n1139), .B1(new_n792), .B2(new_n1220), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n802), .A2(new_n859), .B1(new_n863), .B2(new_n795), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1221), .B(new_n1222), .C1(G150), .C2(new_n1014), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n807), .B2(new_n1134), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT59), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G33), .B(G41), .C1(new_n1086), .C2(G159), .ZN(new_n1226));
  INV_X1    g1026(.A(G124), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1226), .B1(new_n813), .B2(new_n1227), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1219), .B1(KEYINPUT58), .B2(new_n1217), .C1(new_n1225), .C2(new_n1228), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1229), .A2(new_n784), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n852), .B1(G50), .B2(new_n1126), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n1189), .C2(new_n844), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1206), .B2(new_n1006), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1209), .A2(new_n1233), .ZN(G375));
  OAI211_X1 g1034(.A(new_n1215), .B(new_n404), .C1(new_n795), .C2(new_n1134), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n801), .A2(G150), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n863), .B2(new_n792), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G137), .B2(new_n857), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n814), .B2(new_n807), .C1(new_n1139), .C2(new_n813), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1235), .B(new_n1239), .C1(G50), .C2(new_n1014), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n813), .A2(new_n571), .B1(new_n216), .B2(new_n807), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n857), .A2(G283), .B1(new_n796), .B2(new_n532), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1242), .B1(new_n509), .B2(new_n792), .C1(new_n331), .C2(new_n802), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1052), .B(new_n333), .C1(new_n222), .C2(new_n799), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1241), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n784), .B1(new_n1240), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n852), .B1(G68), .B2(new_n1126), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT122), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1116), .B2(new_n844), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1251), .B2(new_n1006), .ZN(new_n1252));
  XOR2_X1   g1052(.A(new_n1252), .B(KEYINPUT123), .Z(new_n1253));
  INV_X1    g1053(.A(new_n984), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1153), .A2(new_n1151), .A3(new_n1155), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1157), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(G381));
  NOR2_X1   g1057(.A1(G375), .A2(G378), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  OR4_X1    g1059(.A1(G396), .A2(G390), .A3(G393), .A4(G384), .ZN(new_n1260));
  OR4_X1    g1060(.A1(G387), .A2(new_n1259), .A3(G381), .A4(new_n1260), .ZN(G407));
  OAI211_X1 g1061(.A(G407), .B(G213), .C1(G343), .C2(new_n1259), .ZN(G409));
  XNOR2_X1  g1062(.A(G393), .B(new_n855), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1007), .A2(new_n1035), .A3(G390), .ZN(new_n1264));
  AOI21_X1  g1064(.A(G390), .B1(new_n1007), .B2(new_n1035), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT125), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1263), .B(new_n1264), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(G393), .B(G396), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT126), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n1007), .B2(new_n1035), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1269), .B1(new_n1271), .B2(G390), .ZN(new_n1272));
  AND3_X1   g1072(.A1(G387), .A2(KEYINPUT126), .A3(G390), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n1267), .A2(new_n1268), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1209), .A2(G378), .A3(new_n1233), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT124), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1169), .A2(new_n1254), .A3(new_n1206), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1277), .A2(new_n1233), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1278), .B2(G378), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1149), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1233), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(KEYINPUT124), .A3(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1275), .A2(new_n1279), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT62), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n709), .A2(G213), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1255), .B(KEYINPUT60), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(new_n736), .A3(new_n1157), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1253), .A2(G384), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G384), .B1(new_n1253), .B2(new_n1287), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .A4(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT61), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1285), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1278), .A2(new_n1276), .A3(G378), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT124), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1293), .B1(new_n1296), .B2(new_n1275), .ZN(new_n1297));
  OAI211_X1 g1097(.A(G2897), .B(new_n1293), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1253), .A2(new_n1287), .ZN(new_n1299));
  INV_X1    g1099(.A(G384), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1253), .A2(G384), .A3(new_n1287), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1293), .A2(G2897), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1298), .A2(new_n1304), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1291), .B(new_n1292), .C1(new_n1297), .C2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1283), .A2(new_n1285), .A3(new_n1290), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1307), .A2(KEYINPUT62), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1274), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1305), .B1(new_n1285), .B2(new_n1283), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT63), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1307), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1297), .A2(KEYINPUT63), .A3(new_n1290), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1274), .A2(KEYINPUT61), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1312), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1309), .A2(new_n1315), .ZN(G405));
  INV_X1    g1116(.A(KEYINPUT127), .ZN(new_n1317));
  AND2_X1   g1117(.A1(new_n1275), .A2(new_n1317), .ZN(new_n1318));
  OR2_X1    g1118(.A1(new_n1274), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(G375), .A2(new_n1280), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1290), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1320), .B(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1274), .A2(new_n1318), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1319), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1322), .B1(new_n1319), .B2(new_n1323), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1324), .A2(new_n1325), .ZN(G402));
endmodule


