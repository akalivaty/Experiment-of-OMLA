//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n612, new_n614, new_n615, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908;
  INV_X1    g000(.A(KEYINPUT34), .ZN(new_n202));
  XOR2_X1   g001(.A(G127gat), .B(G134gat), .Z(new_n203));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(KEYINPUT1), .B2(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G113gat), .B(G120gat), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207));
  XNOR2_X1  g006(.A(G127gat), .B(G134gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT24), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(KEYINPUT24), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n211), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT23), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n219), .B2(new_n216), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n212), .B(KEYINPUT24), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT64), .B(G183gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(G190gat), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n220), .A2(new_n222), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n221), .A2(new_n222), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT26), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n218), .A2(new_n228), .ZN(new_n229));
  MUX2_X1   g028(.A(new_n229), .B(new_n228), .S(new_n216), .Z(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n212), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT28), .ZN(new_n232));
  NOR2_X1   g031(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n233), .B1(new_n224), .B2(KEYINPUT27), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n232), .B1(new_n234), .B2(G190gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT27), .B(G183gat), .ZN(new_n236));
  INV_X1    g035(.A(G190gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(KEYINPUT28), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n231), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n210), .B1(new_n227), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n235), .A2(new_n238), .ZN(new_n241));
  INV_X1    g040(.A(new_n231), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n210), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n225), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n222), .B1(new_n215), .B2(new_n220), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n240), .A2(new_n248), .B1(G227gat), .B2(G233gat), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n202), .B1(new_n250), .B2(KEYINPUT66), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n252));
  NOR3_X1   g051(.A1(new_n249), .A2(new_n252), .A3(KEYINPUT34), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G15gat), .B(G43gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT65), .ZN(new_n256));
  XOR2_X1   g055(.A(G71gat), .B(G99gat), .Z(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n240), .A2(new_n248), .A3(G227gat), .A4(G233gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT33), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(KEYINPUT32), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n259), .B(KEYINPUT32), .C1(new_n260), .C2(new_n258), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n254), .B(new_n265), .Z(new_n266));
  OR2_X1    g065(.A1(new_n266), .A2(KEYINPUT36), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n268), .B1(new_n254), .B2(new_n265), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n254), .A2(new_n265), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n265), .A3(new_n268), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(KEYINPUT36), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G226gat), .ZN(new_n275));
  INV_X1    g074(.A(G233gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(new_n227), .B2(new_n239), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT29), .B1(new_n243), .B2(new_n247), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(new_n277), .ZN(new_n280));
  XNOR2_X1  g079(.A(G211gat), .B(G218gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT68), .ZN(new_n282));
  OR2_X1    g081(.A1(G211gat), .A2(G218gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n284));
  NAND2_X1  g083(.A1(G211gat), .A2(G218gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G204gat), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n288), .A2(G197gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT22), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n288), .A2(G197gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n282), .A2(new_n293), .A3(new_n286), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(KEYINPUT69), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n282), .A2(new_n298), .A3(new_n293), .A4(new_n286), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT70), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT70), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n297), .A2(new_n302), .A3(new_n299), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT71), .B1(new_n280), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n280), .A2(new_n304), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT29), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(new_n227), .B2(new_n239), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(new_n275), .B2(new_n276), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT71), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n301), .A2(new_n303), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n278), .A4(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G8gat), .B(G36gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(G64gat), .B(G92gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n307), .A2(new_n308), .A3(new_n314), .A4(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT30), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n305), .A2(new_n314), .A3(new_n306), .A4(new_n318), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT72), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n314), .A3(new_n306), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n324), .A2(new_n317), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n321), .A2(new_n320), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G1gat), .B(G29gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(KEYINPUT0), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT77), .ZN(new_n331));
  XNOR2_X1  g130(.A(G57gat), .B(G85gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT5), .ZN(new_n334));
  AND2_X1   g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(G141gat), .A2(G148gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(G155gat), .B(G162gat), .Z(new_n339));
  NAND2_X1  g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT2), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n338), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n340), .A2(new_n346), .A3(KEYINPUT2), .ZN(new_n347));
  INV_X1    g146(.A(new_n336), .ZN(new_n348));
  NAND2_X1  g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n346), .B1(new_n340), .B2(KEYINPUT2), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n345), .B(new_n339), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n341), .A2(KEYINPUT73), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(new_n337), .A3(new_n347), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n345), .B1(new_n355), .B2(new_n339), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n210), .B(new_n344), .C1(new_n353), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT76), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n339), .B1(new_n350), .B2(new_n351), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT74), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n352), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT76), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n361), .A2(new_n362), .A3(new_n344), .A4(new_n210), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n343), .B1(new_n360), .B2(new_n352), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n358), .B(new_n363), .C1(new_n364), .C2(new_n210), .ZN(new_n365));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n334), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n244), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n344), .B1(new_n353), .B2(new_n356), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n371), .A2(KEYINPUT3), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n210), .B1(new_n371), .B2(KEYINPUT3), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n364), .A2(new_n369), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT75), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n366), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT4), .B1(new_n358), .B2(new_n363), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n379), .B1(KEYINPUT4), .B2(new_n357), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n368), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n357), .A2(KEYINPUT76), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n362), .B1(new_n364), .B2(new_n210), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT4), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT78), .ZN(new_n385));
  INV_X1    g184(.A(new_n357), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(KEYINPUT4), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n384), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n358), .B2(new_n363), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT78), .B1(new_n391), .B2(new_n387), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n373), .B1(new_n370), .B2(new_n372), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n375), .A2(KEYINPUT75), .A3(new_n376), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n367), .A2(KEYINPUT5), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n389), .A2(new_n392), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n381), .B1(new_n397), .B2(KEYINPUT79), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n397), .A2(KEYINPUT79), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n333), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT6), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n392), .A2(new_n395), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT79), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n403), .A2(new_n404), .A3(new_n389), .A4(new_n396), .ZN(new_n405));
  INV_X1    g204(.A(new_n333), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n397), .A2(KEYINPUT79), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .A4(new_n381), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n400), .A2(new_n401), .A3(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(KEYINPUT6), .B(new_n333), .C1(new_n398), .C2(new_n399), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n328), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G228gat), .A2(G233gat), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n369), .B1(new_n300), .B2(KEYINPUT29), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n412), .B1(new_n413), .B2(new_n371), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n301), .B(new_n303), .C1(new_n372), .C2(KEYINPUT29), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  XOR2_X1   g216(.A(new_n412), .B(KEYINPUT80), .Z(new_n418));
  AOI21_X1  g217(.A(KEYINPUT29), .B1(new_n295), .B2(new_n296), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n371), .B1(new_n419), .B2(KEYINPUT3), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n418), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n417), .A2(new_n421), .A3(G22gat), .ZN(new_n422));
  INV_X1    g221(.A(G22gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n415), .A2(new_n420), .ZN(new_n424));
  INV_X1    g223(.A(new_n418), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n423), .B1(new_n426), .B2(new_n416), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT81), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G78gat), .B(G106gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT31), .B(G50gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n429), .B(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(G22gat), .B1(new_n417), .B2(new_n421), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT81), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n426), .A2(new_n423), .A3(new_n416), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n428), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n431), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n432), .A2(new_n434), .A3(new_n433), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n274), .B1(new_n411), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n409), .A2(KEYINPUT83), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n400), .A2(new_n443), .A3(new_n408), .A4(new_n401), .ZN(new_n444));
  INV_X1    g243(.A(new_n324), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT37), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n280), .B(new_n304), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT38), .B1(new_n448), .B2(KEYINPUT37), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n317), .A3(new_n449), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n450), .A2(new_n322), .A3(new_n319), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n442), .A2(new_n410), .A3(new_n444), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT84), .ZN(new_n453));
  INV_X1    g252(.A(new_n410), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n454), .B1(new_n409), .B2(KEYINPUT83), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n444), .A4(new_n451), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n447), .A2(new_n317), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n445), .A2(new_n446), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT38), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n453), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n389), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n367), .B1(new_n402), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n463), .B(KEYINPUT39), .C1(new_n367), .C2(new_n365), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT39), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n465), .B(new_n367), .C1(new_n402), .C2(new_n462), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT82), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n466), .A2(new_n467), .A3(new_n406), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n467), .B1(new_n466), .B2(new_n406), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n464), .B(KEYINPUT40), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n470), .A2(new_n400), .A3(new_n328), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n439), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n441), .B1(new_n461), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT35), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n323), .A2(new_n327), .A3(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n478), .A2(new_n438), .A3(new_n436), .A4(new_n266), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n444), .B2(new_n455), .ZN(new_n480));
  AND4_X1   g279(.A1(new_n272), .A2(new_n436), .A3(new_n271), .A4(new_n438), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n477), .B1(new_n411), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G15gat), .B(G22gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT16), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n485), .B1(new_n486), .B2(G1gat), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n487), .B(KEYINPUT89), .C1(G1gat), .C2(new_n485), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n488), .B(G8gat), .Z(new_n489));
  OR3_X1    g288(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G29gat), .A2(G36gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(G43gat), .B(G50gat), .Z(new_n495));
  INV_X1    g294(.A(KEYINPUT15), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT86), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT15), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT87), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n491), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n490), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(KEYINPUT87), .B2(new_n490), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n495), .A2(new_n499), .A3(new_n496), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n501), .A2(new_n505), .A3(new_n493), .A4(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n489), .B1(new_n498), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n498), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT88), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n508), .B1(new_n512), .B2(new_n489), .ZN(new_n513));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n515), .A2(KEYINPUT18), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n489), .B(new_n509), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n514), .B(KEYINPUT13), .Z(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n520), .B1(new_n515), .B2(KEYINPUT18), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G113gat), .B(G141gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(G169gat), .B(G197gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(KEYINPUT12), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT90), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT90), .ZN(new_n530));
  INV_X1    g329(.A(new_n528), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n516), .A2(new_n521), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n522), .A2(new_n528), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n484), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G57gat), .B(G64gat), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G71gat), .B(G78gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT21), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G127gat), .B(G155gat), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT20), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n547), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G183gat), .B(G211gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n489), .B1(new_n542), .B2(new_n541), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT92), .Z(new_n554));
  XNOR2_X1  g353(.A(new_n552), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556));
  INV_X1    g355(.A(G85gat), .ZN(new_n557));
  INV_X1    g356(.A(G92gat), .ZN(new_n558));
  AOI22_X1  g357(.A1(KEYINPUT8), .A2(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT94), .ZN(new_n560));
  NAND2_X1  g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT7), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G99gat), .B(G106gat), .Z(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n512), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n565), .ZN(new_n567));
  AND2_X1   g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n567), .A2(new_n509), .B1(KEYINPUT41), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G190gat), .B(G218gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT93), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n568), .A2(KEYINPUT41), .ZN(new_n575));
  XNOR2_X1  g374(.A(G134gat), .B(G162gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n575), .B(new_n576), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT95), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n574), .B(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(G230gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n580), .A2(new_n276), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n565), .B(new_n541), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n582), .A2(KEYINPUT10), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n565), .A2(new_n541), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT10), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n581), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n582), .A2(new_n581), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT96), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G120gat), .B(G148gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(G176gat), .B(G204gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n587), .A2(new_n595), .A3(new_n589), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n555), .A2(new_n579), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n536), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n409), .A2(new_n410), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n601), .B(G1gat), .Z(G1324gat));
  INV_X1    g401(.A(new_n328), .ZN(new_n603));
  OAI21_X1  g402(.A(G8gat), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT42), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT16), .B(G8gat), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n599), .A2(new_n603), .A3(new_n606), .ZN(new_n607));
  MUX2_X1   g406(.A(new_n605), .B(KEYINPUT42), .S(new_n607), .Z(G1325gat));
  OAI21_X1  g407(.A(G15gat), .B1(new_n599), .B2(new_n274), .ZN(new_n609));
  INV_X1    g408(.A(G15gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n266), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n609), .B1(new_n599), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT97), .ZN(G1326gat));
  NOR2_X1   g412(.A1(new_n599), .A2(new_n440), .ZN(new_n614));
  XOR2_X1   g413(.A(KEYINPUT43), .B(G22gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(G1327gat));
  INV_X1    g415(.A(G29gat), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT44), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n452), .A2(KEYINPUT84), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n460), .B1(new_n452), .B2(KEYINPUT84), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n475), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n441), .ZN(new_n622));
  OAI21_X1  g421(.A(KEYINPUT101), .B1(new_n480), .B2(new_n482), .ZN(new_n623));
  INV_X1    g422(.A(new_n479), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n455), .A2(new_n444), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n411), .A2(new_n481), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT35), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n626), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n621), .A2(new_n622), .B1(new_n623), .B2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n574), .B(new_n578), .Z(new_n632));
  OAI21_X1  g431(.A(new_n618), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI211_X1 g432(.A(KEYINPUT44), .B(new_n579), .C1(new_n476), .C2(new_n483), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n600), .ZN(new_n636));
  INV_X1    g435(.A(new_n597), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n535), .A2(new_n555), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT100), .Z(new_n639));
  NAND3_X1  g438(.A1(new_n635), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n617), .B1(new_n640), .B2(KEYINPUT102), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n641), .B1(KEYINPUT102), .B2(new_n640), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n555), .A2(new_n579), .A3(new_n637), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT98), .Z(new_n644));
  NAND3_X1  g443(.A1(new_n484), .A2(new_n535), .A3(new_n644), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n645), .A2(G29gat), .A3(new_n600), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT99), .B(KEYINPUT45), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n642), .A2(new_n648), .ZN(G1328gat));
  NOR3_X1   g448(.A1(new_n645), .A2(G36gat), .A3(new_n603), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT46), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n639), .ZN(new_n652));
  OAI21_X1  g451(.A(G36gat), .B1(new_n652), .B2(new_n603), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT103), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n651), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(G1329gat));
  INV_X1    g457(.A(G43gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n266), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(KEYINPUT104), .Z(new_n662));
  OAI21_X1  g461(.A(G43gat), .B1(new_n652), .B2(new_n274), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT47), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n662), .A2(KEYINPUT47), .A3(new_n663), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(G1330gat));
  NOR3_X1   g467(.A1(new_n645), .A2(G50gat), .A3(new_n440), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n633), .A2(new_n439), .A3(new_n634), .A4(new_n639), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(G50gat), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n670), .A2(KEYINPUT48), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n669), .B1(new_n672), .B2(KEYINPUT105), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n671), .A2(new_n676), .A3(G50gat), .ZN(new_n677));
  AOI211_X1 g476(.A(new_n674), .B(KEYINPUT48), .C1(new_n675), .C2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n672), .A2(KEYINPUT105), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n677), .A3(new_n670), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT48), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT106), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n673), .B1(new_n678), .B2(new_n682), .ZN(G1331gat));
  NOR3_X1   g482(.A1(new_n535), .A2(new_n555), .A3(new_n579), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n631), .A2(new_n637), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n636), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g487(.A(new_n603), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT107), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n691), .B(new_n692), .Z(G1333gat));
  INV_X1    g492(.A(G71gat), .ZN(new_n694));
  INV_X1    g493(.A(new_n274), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n686), .B2(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n266), .A2(new_n694), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(new_n686), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g498(.A1(new_n686), .A2(new_n439), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g500(.A1(new_n621), .A2(new_n622), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n623), .A2(new_n630), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n632), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n555), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n535), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT51), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT51), .ZN(new_n708));
  INV_X1    g507(.A(new_n706), .ZN(new_n709));
  NOR4_X1   g508(.A1(new_n631), .A2(new_n708), .A3(new_n632), .A4(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n597), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(new_n557), .A3(new_n636), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n705), .A2(new_n535), .A3(new_n637), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n635), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n716), .B2(new_n600), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G85gat), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n716), .A2(new_n714), .A3(new_n600), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n713), .B1(new_n718), .B2(new_n719), .ZN(G1336gat));
  NAND4_X1  g519(.A1(new_n635), .A2(G92gat), .A3(new_n328), .A4(new_n715), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n711), .A2(new_n603), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(G92gat), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI211_X1 g524(.A(KEYINPUT52), .B(new_n721), .C1(new_n722), .C2(G92gat), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(G1337gat));
  AOI21_X1  g526(.A(G99gat), .B1(new_n712), .B2(new_n266), .ZN(new_n728));
  INV_X1    g527(.A(G99gat), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n716), .A2(new_n729), .A3(new_n274), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n728), .A2(new_n730), .ZN(G1338gat));
  NOR2_X1   g530(.A1(new_n440), .A2(G106gat), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n597), .B(new_n732), .C1(new_n707), .C2(new_n710), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n633), .A2(new_n439), .A3(new_n634), .A4(new_n715), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G106gat), .ZN(new_n735));
  NAND2_X1  g534(.A1(KEYINPUT109), .A2(KEYINPUT53), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n733), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT110), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT109), .A2(KEYINPUT53), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n734), .A2(G106gat), .B1(KEYINPUT109), .B2(KEYINPUT53), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n740), .A2(new_n741), .A3(new_n733), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n738), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n739), .B1(new_n738), .B2(new_n742), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(G1339gat));
  NAND2_X1  g544(.A1(new_n684), .A2(new_n637), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n583), .A2(new_n585), .A3(new_n581), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n587), .A2(KEYINPUT54), .A3(new_n747), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n749));
  AOI21_X1  g548(.A(new_n595), .B1(new_n586), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n748), .A2(KEYINPUT55), .A3(new_n750), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(new_n596), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n513), .A2(new_n514), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n517), .A2(new_n519), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n527), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n529), .B2(new_n532), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n756), .A2(new_n760), .A3(new_n579), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n755), .A2(new_n632), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n764), .A2(KEYINPUT112), .A3(new_n760), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n760), .A2(new_n597), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n533), .A2(new_n534), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(new_n755), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n763), .A2(new_n765), .B1(new_n768), .B2(new_n632), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n746), .B1(new_n769), .B2(new_n705), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n600), .A2(new_n328), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n266), .A2(new_n436), .A3(new_n438), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(G113gat), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n774), .A2(new_n775), .A3(new_n767), .ZN(new_n776));
  INV_X1    g575(.A(new_n772), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(new_n481), .A3(new_n535), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n776), .B1(new_n775), .B2(new_n778), .ZN(G1340gat));
  OAI21_X1  g578(.A(G120gat), .B1(new_n774), .B2(new_n637), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n481), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n637), .A2(G120gat), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT113), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n780), .B1(new_n781), .B2(new_n783), .ZN(G1341gat));
  INV_X1    g583(.A(G127gat), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n774), .A2(new_n785), .A3(new_n555), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n781), .A2(KEYINPUT114), .A3(new_n555), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(G127gat), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT114), .B1(new_n781), .B2(new_n555), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n786), .B1(new_n788), .B2(new_n789), .ZN(G1342gat));
  INV_X1    g589(.A(new_n481), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(G134gat), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n770), .A2(new_n579), .A3(new_n771), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT56), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT116), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n793), .A2(KEYINPUT56), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT115), .ZN(new_n798));
  OAI21_X1  g597(.A(G134gat), .B1(new_n774), .B2(new_n632), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n796), .A2(new_n798), .A3(KEYINPUT117), .A4(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n797), .A2(KEYINPUT115), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n797), .A2(KEYINPUT115), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n801), .B1(new_n804), .B2(new_n795), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n800), .A2(new_n805), .ZN(G1343gat));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807));
  INV_X1    g606(.A(new_n746), .ZN(new_n808));
  AND4_X1   g607(.A1(KEYINPUT112), .A2(new_n756), .A3(new_n579), .A4(new_n760), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT112), .B1(new_n764), .B2(new_n760), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n756), .A2(new_n535), .B1(new_n597), .B2(new_n760), .ZN(new_n811));
  OAI22_X1  g610(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(new_n579), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n808), .B1(new_n812), .B2(new_n555), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n807), .B1(new_n813), .B2(new_n440), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n770), .A2(KEYINPUT57), .A3(new_n439), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n771), .A2(new_n274), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT118), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  AND4_X1   g618(.A1(KEYINPUT120), .A2(new_n816), .A3(new_n535), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n818), .B1(new_n814), .B2(new_n815), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT120), .B1(new_n821), .B2(new_n535), .ZN(new_n822));
  OAI21_X1  g621(.A(G141gat), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n695), .A2(new_n440), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n772), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(G141gat), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n827), .A3(new_n535), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n823), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n535), .A3(new_n819), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(G141gat), .ZN(new_n833));
  AOI211_X1 g632(.A(KEYINPUT119), .B(new_n829), .C1(new_n833), .C2(new_n828), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n835));
  AOI211_X1 g634(.A(new_n767), .B(new_n818), .C1(new_n814), .C2(new_n815), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n828), .B1(new_n836), .B2(new_n827), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n837), .B2(KEYINPUT58), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n831), .B1(new_n834), .B2(new_n838), .ZN(G1344gat));
  INV_X1    g638(.A(G148gat), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n777), .A2(new_n840), .A3(new_n597), .A4(new_n824), .ZN(new_n841));
  AOI211_X1 g640(.A(KEYINPUT59), .B(new_n840), .C1(new_n821), .C2(new_n597), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n761), .B1(new_n811), .B2(new_n579), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n808), .B1(new_n844), .B2(new_n555), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n807), .B1(new_n845), .B2(new_n440), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n637), .B1(new_n815), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n840), .B1(new_n847), .B2(new_n819), .ZN(new_n848));
  OAI22_X1  g647(.A1(new_n842), .A2(KEYINPUT121), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n821), .A2(new_n597), .ZN(new_n850));
  AND4_X1   g649(.A1(KEYINPUT121), .A2(new_n850), .A3(new_n843), .A4(G148gat), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n841), .B1(new_n849), .B2(new_n851), .ZN(G1345gat));
  INV_X1    g651(.A(G155gat), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n826), .A2(new_n853), .A3(new_n705), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n821), .A2(new_n705), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(new_n853), .ZN(G1346gat));
  OR4_X1    g655(.A1(G162gat), .A2(new_n772), .A3(new_n632), .A4(new_n825), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n821), .A2(new_n579), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n858), .A2(KEYINPUT122), .ZN(new_n859));
  OAI21_X1  g658(.A(G162gat), .B1(new_n858), .B2(KEYINPUT122), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(G1347gat));
  NOR2_X1   g660(.A1(new_n813), .A2(new_n636), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n328), .A3(new_n481), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(G169gat), .B1(new_n864), .B2(new_n535), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n636), .A2(new_n603), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n813), .A2(new_n773), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n535), .A2(G169gat), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(G1348gat));
  NAND3_X1  g669(.A1(new_n868), .A2(G176gat), .A3(new_n597), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT123), .ZN(new_n872));
  AOI21_X1  g671(.A(G176gat), .B1(new_n864), .B2(new_n597), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(G1349gat));
  AND2_X1   g673(.A1(new_n705), .A2(new_n236), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n868), .A2(new_n705), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n864), .A2(new_n875), .B1(new_n876), .B2(new_n224), .ZN(new_n877));
  XOR2_X1   g676(.A(new_n877), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g677(.A1(new_n864), .A2(new_n237), .A3(new_n579), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n237), .B1(new_n868), .B2(new_n579), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n882), .A2(KEYINPUT124), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n881), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(new_n882), .B2(KEYINPUT124), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n879), .B1(new_n883), .B2(new_n885), .ZN(G1351gat));
  NAND3_X1  g685(.A1(new_n862), .A2(new_n328), .A3(new_n824), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(G197gat), .A3(new_n767), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT125), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n815), .A2(new_n846), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n867), .A2(new_n695), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n767), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n893), .A2(KEYINPUT126), .ZN(new_n894));
  OAI21_X1  g693(.A(G197gat), .B1(new_n893), .B2(KEYINPUT126), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n889), .B1(new_n894), .B2(new_n895), .ZN(G1352gat));
  NOR3_X1   g695(.A1(new_n887), .A2(G204gat), .A3(new_n637), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT62), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n847), .A2(new_n891), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n288), .B2(new_n899), .ZN(G1353gat));
  OR3_X1    g699(.A1(new_n887), .A2(G211gat), .A3(new_n555), .ZN(new_n901));
  OAI21_X1  g700(.A(G211gat), .B1(new_n892), .B2(new_n555), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT63), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n902), .A2(new_n903), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(G1354gat));
  OAI21_X1  g705(.A(G218gat), .B1(new_n892), .B2(new_n632), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n632), .A2(G218gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n887), .B2(new_n908), .ZN(G1355gat));
endmodule


