//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT27), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT26), .B(G101), .Z(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT28), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n196));
  INV_X1    g010(.A(G113), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT2), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G113), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G116), .B(G119), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n203));
  NOR3_X1   g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT2), .B(G113), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G116), .ZN(new_n207));
  INV_X1    g021(.A(G116), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G119), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n205), .B1(KEYINPUT66), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n196), .B1(new_n204), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n201), .B1(new_n202), .B2(new_n203), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n205), .A3(KEYINPUT66), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT67), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT64), .B(G143), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n219), .B1(new_n220), .B2(G146), .ZN(new_n221));
  AND2_X1   g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  OR2_X1    g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n217), .A2(G143), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(new_n220), .B2(G146), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n221), .A2(new_n225), .B1(new_n228), .B2(new_n222), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n230));
  INV_X1    g044(.A(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G137), .ZN(new_n232));
  INV_X1    g046(.A(G137), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT11), .A3(G134), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(G137), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G131), .ZN(new_n237));
  INV_X1    g051(.A(G131), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n232), .A2(new_n234), .A3(new_n238), .A4(new_n235), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G143), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT64), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT64), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G143), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n244), .A3(G146), .ZN(new_n245));
  INV_X1    g059(.A(G128), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(KEYINPUT1), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n226), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n242), .A2(new_n244), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n218), .B1(new_n249), .B2(new_n217), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n246), .B1(new_n226), .B2(KEYINPUT1), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n233), .A2(KEYINPUT65), .A3(G134), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n231), .B2(G137), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n233), .A2(G134), .ZN(new_n256));
  OAI211_X1 g070(.A(G131), .B(new_n253), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n239), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n229), .A2(new_n240), .B1(new_n252), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n216), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n252), .A2(new_n259), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n221), .A2(new_n225), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n245), .A2(new_n226), .A3(new_n222), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n240), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(KEYINPUT69), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n195), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT67), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT67), .B1(new_n213), .B2(new_n214), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n263), .A2(new_n266), .B1(new_n213), .B2(new_n214), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT28), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n194), .B1(new_n269), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n237), .A2(new_n239), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n265), .B1(new_n250), .B2(new_n224), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n251), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n221), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n258), .B1(new_n282), .B2(new_n248), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT30), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT30), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n263), .A2(new_n266), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n213), .A2(new_n214), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n193), .B1(new_n260), .B2(new_n216), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n287), .A2(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n194), .B1(new_n267), .B2(new_n272), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT68), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT31), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n263), .A2(new_n266), .A3(new_n285), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n285), .B1(new_n263), .B2(new_n266), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n288), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n216), .A2(new_n263), .A3(new_n266), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(new_n290), .A3(new_n194), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n293), .A2(new_n297), .A3(KEYINPUT31), .A4(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n277), .B1(new_n294), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(G472), .A2(G902), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n187), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n293), .A2(new_n297), .A3(new_n299), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT31), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n276), .B1(new_n307), .B2(new_n300), .ZN(new_n308));
  INV_X1    g122(.A(new_n303), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n308), .A2(KEYINPUT32), .A3(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G472), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT70), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n297), .A2(new_n298), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT29), .B1(new_n314), .B2(new_n193), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n269), .A2(new_n275), .A3(new_n194), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n193), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n272), .B1(new_n280), .B2(new_n283), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n298), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n320), .B1(new_n322), .B2(KEYINPUT28), .ZN(new_n323));
  AOI211_X1 g137(.A(KEYINPUT71), .B(new_n195), .C1(new_n321), .C2(new_n298), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n269), .B(new_n319), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G902), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n317), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n315), .A2(new_n313), .A3(new_n316), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n312), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT72), .B1(new_n311), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT76), .B(KEYINPUT25), .Z(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n206), .A2(G128), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT23), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT73), .B1(new_n246), .B2(G119), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n206), .A2(G128), .ZN(new_n339));
  OAI211_X1 g153(.A(KEYINPUT23), .B(new_n335), .C1(new_n339), .C2(KEYINPUT73), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n339), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n342), .A2(new_n335), .ZN(new_n343));
  XOR2_X1   g157(.A(KEYINPUT24), .B(G110), .Z(new_n344));
  AOI22_X1  g158(.A1(new_n341), .A2(G110), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(G125), .B(G140), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(KEYINPUT74), .A3(KEYINPUT16), .ZN(new_n347));
  INV_X1    g161(.A(G140), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G125), .ZN(new_n349));
  INV_X1    g163(.A(G125), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G140), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n351), .A3(KEYINPUT16), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n349), .B2(KEYINPUT16), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n347), .B(new_n217), .C1(new_n353), .C2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n352), .B(new_n354), .C1(KEYINPUT16), .C2(new_n349), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n217), .B1(new_n358), .B2(new_n347), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n345), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  OAI22_X1  g174(.A1(new_n341), .A2(G110), .B1(new_n343), .B2(new_n344), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n347), .B1(new_n353), .B2(new_n355), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G146), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n346), .A2(new_n217), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n366), .B(KEYINPUT75), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT22), .B(G137), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n360), .A2(new_n365), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n369), .B1(new_n360), .B2(new_n365), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n334), .B1(new_n373), .B2(new_n326), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n360), .A2(new_n365), .ZN(new_n375));
  INV_X1    g189(.A(new_n369), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n377), .A2(new_n378), .A3(new_n326), .A4(new_n370), .ZN(new_n379));
  INV_X1    g193(.A(G217), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(G234), .B2(new_n326), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n332), .B1(new_n374), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n377), .A2(new_n370), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n333), .B1(new_n384), .B2(G902), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n385), .A2(KEYINPUT77), .A3(new_n379), .A4(new_n381), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n381), .A2(G902), .ZN(new_n387));
  XOR2_X1   g201(.A(new_n387), .B(KEYINPUT78), .Z(new_n388));
  NAND2_X1  g202(.A1(new_n373), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n383), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n302), .A2(new_n187), .A3(new_n303), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT32), .B1(new_n308), .B2(new_n309), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n273), .B1(new_n287), .B2(new_n288), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n318), .B1(new_n395), .B2(new_n194), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n272), .B1(new_n267), .B2(KEYINPUT69), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n260), .A2(new_n261), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT28), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n267), .A2(new_n288), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n195), .B1(new_n400), .B2(new_n298), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n399), .A2(new_n401), .A3(new_n193), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT70), .B1(new_n396), .B2(new_n402), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n403), .A2(new_n326), .A3(new_n329), .A4(new_n325), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G472), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT72), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n394), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n331), .A2(new_n391), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT20), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n188), .A2(new_n189), .A3(G143), .A4(G214), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n410), .B1(new_n249), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G131), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n220), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n238), .A3(new_n410), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT92), .B1(new_n417), .B2(KEYINPUT17), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n357), .A2(new_n359), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n412), .A2(KEYINPUT17), .A3(G131), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT91), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n238), .B1(new_n415), .B2(new_n410), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT91), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT17), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT92), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT17), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n413), .A2(new_n426), .A3(new_n427), .A4(new_n416), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n418), .A2(new_n419), .A3(new_n425), .A4(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(G113), .B(G122), .ZN(new_n430));
  INV_X1    g244(.A(G104), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(KEYINPUT18), .A2(G131), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n415), .A2(new_n410), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n349), .A2(new_n351), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G146), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n364), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n422), .A2(KEYINPUT18), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n429), .A2(new_n432), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT90), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT19), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n435), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n346), .A2(KEYINPUT19), .ZN(new_n445));
  AOI21_X1  g259(.A(G146), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n417), .A2(new_n363), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n440), .ZN(new_n449));
  INV_X1    g263(.A(new_n432), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n442), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI211_X1 g265(.A(KEYINPUT90), .B(new_n432), .C1(new_n448), .C2(new_n440), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n441), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(G475), .A2(G902), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT93), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n409), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n453), .A2(new_n409), .A3(new_n456), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n429), .A2(new_n432), .A3(new_n440), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n432), .B1(new_n429), .B2(new_n440), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n326), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n458), .A2(new_n459), .B1(G475), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(G234), .A2(G237), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n464), .A2(G952), .A3(new_n189), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n464), .A2(G902), .A3(G953), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(G898), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G478), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(KEYINPUT15), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n220), .A2(G128), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n246), .A2(G143), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n231), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(G116), .B(G122), .ZN(new_n475));
  INV_X1    g289(.A(G107), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n472), .A2(KEYINPUT13), .A3(new_n473), .ZN(new_n478));
  OAI21_X1  g292(.A(G134), .B1(new_n472), .B2(KEYINPUT13), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n474), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G122), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G116), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n476), .B1(new_n482), .B2(KEYINPUT14), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(new_n475), .ZN(new_n484));
  INV_X1    g298(.A(new_n474), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n231), .B1(new_n472), .B2(new_n473), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT9), .B(G234), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT79), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n489), .A2(G217), .A3(new_n189), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n480), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n490), .B1(new_n480), .B2(new_n487), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n326), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n471), .B1(new_n493), .B2(KEYINPUT94), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(KEYINPUT94), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT94), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n496), .B(new_n326), .C1(new_n491), .C2(new_n492), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n494), .B1(new_n498), .B2(new_n471), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n463), .A2(KEYINPUT95), .A3(new_n469), .A4(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT95), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n462), .A2(G475), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n446), .B1(G146), .B2(new_n362), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n503), .A2(new_n417), .B1(new_n439), .B2(new_n438), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT90), .B1(new_n504), .B2(new_n432), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n449), .A2(new_n442), .A3(new_n450), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI211_X1 g321(.A(KEYINPUT20), .B(new_n455), .C1(new_n507), .C2(new_n441), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n499), .B(new_n502), .C1(new_n457), .C2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n501), .B1(new_n509), .B2(new_n468), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n500), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(G214), .B1(G237), .B2(G902), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  XOR2_X1   g327(.A(G110), .B(G122), .Z(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT84), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT8), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT3), .B1(new_n431), .B2(G107), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT3), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n476), .A3(G104), .ZN(new_n519));
  INV_X1    g333(.A(G101), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n431), .A2(G107), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n517), .A2(new_n519), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n476), .A2(G104), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n431), .A2(G107), .ZN(new_n524));
  OAI21_X1  g338(.A(G101), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT5), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT5), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n206), .A3(G116), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n527), .A2(KEYINPUT83), .A3(G113), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n201), .A2(new_n202), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n529), .A2(G113), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT83), .B1(new_n533), .B2(new_n527), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n526), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n526), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n527), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n531), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n282), .A2(new_n350), .A3(new_n248), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n229), .B2(new_n350), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n189), .A2(G224), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT88), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT7), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n544), .B2(new_n545), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n516), .A2(new_n539), .B1(new_n541), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT80), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n517), .A2(new_n519), .A3(new_n521), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n550), .A2(G101), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n522), .A2(KEYINPUT4), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n549), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(G101), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n554), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n522), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT4), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n550), .A2(new_n557), .A3(G101), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n288), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n532), .A2(new_n534), .A3(new_n526), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(new_n563), .A3(new_n515), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT86), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n243), .A2(G143), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n241), .A2(KEYINPUT64), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n217), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n224), .B1(new_n568), .B2(new_n219), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n245), .A2(new_n226), .A3(new_n222), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n565), .B(G125), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n540), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n565), .B1(new_n279), .B2(G125), .ZN(new_n573));
  NOR4_X1   g387(.A1(new_n572), .A2(new_n573), .A3(new_n545), .A4(new_n543), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT89), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n548), .B(new_n564), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n574), .A2(new_n575), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(G902), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT85), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n515), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n559), .B1(new_n553), .B2(new_n555), .ZN(new_n583));
  OAI211_X1 g397(.A(KEYINPUT6), .B(new_n582), .C1(new_n583), .C2(new_n562), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT6), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n562), .B1(new_n556), .B2(new_n560), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n585), .B1(new_n586), .B2(new_n515), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n582), .B1(new_n583), .B2(new_n562), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n584), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT87), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n572), .A2(new_n573), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(new_n542), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n591), .B1(new_n590), .B2(new_n593), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n580), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(G210), .B1(G237), .B2(G902), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n584), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n564), .A2(KEYINPUT6), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n600), .B1(new_n601), .B2(new_n588), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n592), .B(new_n543), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT87), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n597), .A3(new_n580), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n513), .B1(new_n599), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n489), .A2(new_n326), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n609), .A2(G221), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT81), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n522), .A2(new_n525), .A3(KEYINPUT10), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n252), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n611), .B1(new_n252), .B2(new_n612), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n279), .B1(new_n557), .B2(new_n551), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n556), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n618));
  INV_X1    g432(.A(new_n248), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n245), .A2(new_n226), .ZN(new_n620));
  AOI21_X1  g434(.A(G146), .B1(new_n242), .B2(new_n244), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT1), .ZN(new_n622));
  OAI21_X1  g436(.A(G128), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n619), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n618), .B1(new_n624), .B2(new_n526), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n615), .A2(new_n617), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n240), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n615), .A2(new_n617), .A3(new_n278), .A4(new_n625), .ZN(new_n628));
  XNOR2_X1  g442(.A(G110), .B(G140), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n189), .A2(G227), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n623), .A2(new_n620), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n526), .B1(new_n634), .B2(new_n248), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n252), .A2(new_n536), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n240), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT82), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT12), .B1(new_n240), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  OAI221_X1 g454(.A(new_n240), .B1(new_n638), .B2(KEYINPUT12), .C1(new_n635), .C2(new_n636), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n628), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n627), .A2(new_n633), .B1(new_n643), .B2(new_n631), .ZN(new_n644));
  OAI21_X1  g458(.A(G469), .B1(new_n644), .B2(G902), .ZN(new_n645));
  INV_X1    g459(.A(G469), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n642), .A2(new_n628), .A3(new_n632), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n632), .B1(new_n627), .B2(new_n628), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n646), .B(new_n326), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n610), .B1(new_n645), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n511), .A2(new_n608), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n408), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n520), .ZN(G3));
  NAND2_X1  g467(.A1(new_n599), .A2(new_n607), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n502), .B1(new_n508), .B2(new_n457), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n493), .A2(KEYINPUT97), .A3(new_n470), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT97), .B1(new_n493), .B2(new_n470), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n480), .A2(new_n487), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT96), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(KEYINPUT33), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n661), .B1(new_n491), .B2(new_n492), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n491), .A2(new_n492), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(KEYINPUT33), .A3(new_n660), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n326), .A2(G478), .ZN(new_n666));
  OAI22_X1  g480(.A1(new_n656), .A2(new_n657), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n655), .A2(new_n667), .A3(new_n469), .ZN(new_n668));
  AND4_X1   g482(.A1(KEYINPUT98), .A2(new_n654), .A3(new_n512), .A4(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT98), .B1(new_n608), .B2(new_n668), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n650), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n390), .ZN(new_n673));
  OAI21_X1  g487(.A(G472), .B1(new_n308), .B2(G902), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n302), .A2(new_n303), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G104), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT99), .B(KEYINPUT34), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G6));
  NAND2_X1  g496(.A1(new_n498), .A2(new_n471), .ZN(new_n683));
  INV_X1    g497(.A(new_n494), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n685), .B(new_n502), .C1(new_n457), .C2(new_n508), .ZN(new_n686));
  OAI21_X1  g500(.A(KEYINPUT100), .B1(new_n686), .B2(new_n468), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT100), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n463), .A2(new_n688), .A3(new_n469), .A4(new_n685), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n608), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n608), .A2(new_n687), .A3(new_n689), .A4(KEYINPUT101), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n678), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT102), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT35), .B(G107), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G9));
  NOR2_X1   g511(.A1(new_n376), .A2(KEYINPUT36), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(new_n375), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n388), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n383), .A2(new_n386), .A3(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n610), .ZN(new_n702));
  INV_X1    g516(.A(new_n649), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n643), .A2(new_n631), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n627), .A2(new_n628), .A3(new_n632), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n704), .A2(G469), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(G469), .A2(G902), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n701), .B(new_n702), .C1(new_n703), .C2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n676), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n511), .A2(new_n710), .A3(new_n608), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT37), .B(G110), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G12));
  INV_X1    g527(.A(new_n465), .ZN(new_n714));
  INV_X1    g528(.A(new_n466), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n714), .B1(new_n715), .B2(G900), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n463), .A2(new_n685), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n709), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n331), .A2(new_n718), .A3(new_n407), .A4(new_n608), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G128), .ZN(G30));
  NOR4_X1   g534(.A1(new_n463), .A2(new_n701), .A3(new_n513), .A4(new_n499), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n291), .A2(new_n293), .B1(new_n193), .B2(new_n322), .ZN(new_n722));
  OAI21_X1  g536(.A(G472), .B1(new_n722), .B2(G902), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n394), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n716), .B(KEYINPUT39), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n650), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n725), .B1(KEYINPUT40), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n654), .B(KEYINPUT38), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n728), .B(new_n729), .C1(KEYINPUT40), .C2(new_n727), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n249), .ZN(G45));
  NAND3_X1  g545(.A1(new_n655), .A2(new_n667), .A3(new_n716), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n709), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n331), .A2(new_n407), .A3(new_n608), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G146), .ZN(G48));
  NOR2_X1   g549(.A1(new_n647), .A2(new_n648), .ZN(new_n736));
  OAI21_X1  g550(.A(G469), .B1(new_n736), .B2(G902), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n649), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n610), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n331), .A2(new_n391), .A3(new_n407), .A4(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n670), .B2(new_n669), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT41), .B(G113), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G15));
  AOI21_X1  g558(.A(new_n740), .B1(new_n692), .B2(new_n693), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT103), .B(G116), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G18));
  AND2_X1   g561(.A1(new_n608), .A2(new_n739), .ZN(new_n748));
  INV_X1    g562(.A(new_n701), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n749), .B1(new_n500), .B2(new_n510), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n748), .A2(new_n331), .A3(new_n407), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G119), .ZN(G21));
  NOR2_X1   g566(.A1(new_n463), .A2(new_n499), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n608), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n323), .A2(new_n324), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n193), .B1(new_n755), .B2(new_n399), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n756), .B1(new_n294), .B2(new_n301), .ZN(new_n757));
  XOR2_X1   g571(.A(new_n303), .B(KEYINPUT104), .Z(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n674), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n390), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n754), .A2(new_n469), .A3(new_n739), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  NOR2_X1   g577(.A1(new_n760), .A2(new_n749), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n655), .A2(new_n667), .A3(new_n716), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n764), .A2(new_n608), .A3(new_n765), .A4(new_n739), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G125), .ZN(G27));
  NAND3_X1  g581(.A1(new_n599), .A2(new_n607), .A3(new_n512), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n768), .A2(new_n672), .A3(new_n732), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT105), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n394), .A2(new_n405), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n770), .B1(new_n771), .B2(new_n391), .ZN(new_n772));
  AOI211_X1 g586(.A(KEYINPUT105), .B(new_n390), .C1(new_n394), .C2(new_n405), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n769), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT42), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n394), .A2(new_n405), .A3(new_n406), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n406), .B1(new_n394), .B2(new_n405), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT42), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n778), .A2(new_n769), .A3(new_n779), .A4(new_n391), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  INV_X1    g596(.A(KEYINPUT106), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n717), .B(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n768), .A2(new_n672), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n778), .A2(new_n784), .A3(new_n391), .A4(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  NAND2_X1  g601(.A1(new_n463), .A2(new_n667), .ZN(new_n788));
  NAND2_X1  g602(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n791));
  OAI21_X1  g605(.A(new_n790), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n677), .A2(new_n749), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n768), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n792), .A2(KEYINPUT44), .A3(new_n793), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n644), .A2(KEYINPUT45), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n644), .A2(KEYINPUT45), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(G469), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT46), .B1(new_n802), .B2(new_n707), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n703), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(KEYINPUT46), .A3(new_n707), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n610), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n726), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n799), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(new_n233), .ZN(G39));
  NOR3_X1   g623(.A1(new_n768), .A2(new_n391), .A3(new_n732), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n806), .A2(KEYINPUT47), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n806), .A2(KEYINPUT47), .ZN(new_n812));
  OAI221_X1 g626(.A(new_n810), .B1(new_n777), .B2(new_n776), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G140), .ZN(G42));
  XNOR2_X1  g628(.A(new_n738), .B(KEYINPUT108), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(KEYINPUT49), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT109), .ZN(new_n817));
  INV_X1    g631(.A(new_n729), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n815), .A2(KEYINPUT49), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n391), .A2(new_n512), .A3(new_n702), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n724), .A2(new_n820), .A3(new_n788), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n817), .A2(new_n818), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n792), .A2(new_n465), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT114), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n761), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n739), .A2(new_n513), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT115), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n818), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT50), .ZN(new_n831));
  INV_X1    g645(.A(new_n826), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n811), .A2(new_n812), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n815), .A2(new_n702), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n832), .B(new_n797), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n797), .A2(new_n739), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n824), .A2(new_n836), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n836), .A2(new_n390), .A3(new_n714), .A4(new_n724), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n655), .A2(new_n667), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n837), .A2(new_n764), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n831), .A2(KEYINPUT51), .A3(new_n835), .A4(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n830), .A2(KEYINPUT50), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT50), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n826), .A2(new_n843), .A3(new_n829), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n835), .B(new_n840), .C1(new_n842), .C2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT51), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n772), .A2(new_n773), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n837), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n832), .A2(new_n748), .ZN(new_n853));
  INV_X1    g667(.A(G952), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n655), .A2(new_n667), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  AOI211_X1 g670(.A(new_n854), .B(G953), .C1(new_n838), .C2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n852), .A2(new_n853), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n849), .A2(new_n851), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n841), .A2(new_n847), .A3(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n751), .B(new_n762), .C1(new_n671), .C2(new_n740), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n468), .B1(new_n686), .B2(new_n855), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n673), .A2(new_n608), .A3(new_n863), .A4(new_n677), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n864), .B(new_n711), .C1(new_n408), .C2(new_n651), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n862), .A2(new_n745), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n645), .A2(new_n649), .ZN(new_n867));
  AND4_X1   g681(.A1(new_n702), .A2(new_n867), .A3(new_n749), .A4(new_n716), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(new_n608), .A3(new_n724), .A4(new_n753), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n719), .A2(new_n734), .A3(new_n766), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT110), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n597), .B1(new_n606), .B2(new_n580), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n326), .B1(new_n576), .B2(new_n578), .ZN(new_n873));
  AOI211_X1 g687(.A(new_n598), .B(new_n873), .C1(new_n604), .C2(new_n605), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n512), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n875), .A2(new_n709), .A3(new_n717), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n765), .A2(new_n650), .A3(new_n701), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n875), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n778), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT110), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(new_n880), .A3(new_n766), .A4(new_n869), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n871), .A2(new_n881), .A3(KEYINPUT52), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n768), .A2(new_n672), .A3(new_n749), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n463), .A2(new_n499), .A3(new_n716), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n776), .A2(new_n777), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n760), .A2(new_n732), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AND4_X1   g701(.A1(new_n775), .A2(new_n887), .A3(new_n780), .A4(new_n786), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n866), .A2(new_n882), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT52), .B1(new_n871), .B2(new_n881), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n865), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n751), .A2(new_n762), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n692), .A2(new_n693), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n741), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n893), .A2(new_n894), .A3(new_n742), .A4(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n775), .A2(new_n887), .A3(new_n780), .A4(new_n786), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n870), .A2(KEYINPUT52), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n871), .A2(new_n881), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT52), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT53), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT54), .B1(new_n892), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT113), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n890), .B1(new_n889), .B2(new_n891), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT112), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n862), .B2(new_n745), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n894), .A2(new_n742), .A3(new_n896), .A4(KEYINPUT112), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n893), .A2(KEYINPUT53), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n903), .A2(new_n911), .A3(new_n888), .A4(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n907), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n905), .A2(new_n906), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n906), .B1(new_n905), .B2(new_n915), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n861), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(G952), .A2(G953), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n822), .B1(new_n918), .B2(new_n919), .ZN(G75));
  NOR2_X1   g734(.A1(new_n189), .A2(G952), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n326), .B1(new_n907), .B2(new_n913), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(G210), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n590), .B(KEYINPUT117), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT55), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n603), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n928), .A2(KEYINPUT56), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n922), .B1(new_n925), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT56), .B1(new_n924), .B2(KEYINPUT118), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(KEYINPUT118), .B2(new_n924), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n930), .B1(new_n932), .B2(new_n928), .ZN(G51));
  AOI211_X1 g747(.A(new_n326), .B(new_n802), .C1(new_n907), .C2(new_n913), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n907), .A2(new_n913), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT54), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n915), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n707), .B(KEYINPUT57), .Z(new_n938));
  AOI21_X1  g752(.A(new_n736), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n934), .B1(new_n939), .B2(KEYINPUT119), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT119), .ZN(new_n941));
  INV_X1    g755(.A(new_n938), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n936), .B2(new_n915), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n941), .B1(new_n943), .B2(new_n736), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n921), .B1(new_n940), .B2(new_n944), .ZN(G54));
  NAND3_X1  g759(.A1(new_n923), .A2(KEYINPUT58), .A3(G475), .ZN(new_n946));
  INV_X1    g760(.A(new_n453), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n948), .A2(new_n949), .A3(new_n921), .ZN(G60));
  INV_X1    g764(.A(new_n937), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n665), .B(KEYINPUT120), .ZN(new_n952));
  NAND2_X1  g766(.A1(G478), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT59), .Z(new_n954));
  OR2_X1    g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n922), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n954), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n916), .B2(new_n917), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n956), .B1(new_n958), .B2(new_n952), .ZN(G63));
  NAND2_X1  g773(.A1(G217), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT60), .Z(new_n961));
  NAND3_X1  g775(.A1(new_n935), .A2(new_n699), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n962), .A2(KEYINPUT121), .A3(new_n922), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT61), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n935), .A2(new_n961), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n922), .B(new_n962), .C1(new_n965), .C2(new_n373), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n964), .B(new_n966), .ZN(G66));
  INV_X1    g781(.A(new_n467), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n189), .B1(new_n968), .B2(G224), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n897), .B2(new_n189), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n926), .B1(G898), .B2(new_n189), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n970), .B(new_n971), .Z(G69));
  NOR2_X1   g786(.A1(new_n189), .A2(G900), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n781), .A2(new_n786), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n974), .A2(KEYINPUT125), .ZN(new_n975));
  INV_X1    g789(.A(new_n808), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n879), .A2(new_n766), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n848), .A2(new_n806), .A3(new_n726), .A4(new_n754), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n974), .A2(KEYINPUT125), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n975), .A2(new_n979), .A3(new_n813), .A4(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n973), .B1(new_n981), .B2(new_n189), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n444), .A2(new_n445), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n287), .B(new_n983), .Z(new_n984));
  OR2_X1    g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT124), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT126), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n977), .A2(new_n730), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT123), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n727), .B1(new_n855), .B2(new_n686), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n778), .A2(new_n994), .A3(new_n391), .A4(new_n797), .ZN(new_n995));
  AND4_X1   g809(.A1(new_n976), .A2(new_n993), .A3(new_n813), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n189), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n984), .B(KEYINPUT122), .Z(new_n999));
  AOI21_X1  g813(.A(new_n989), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n987), .A2(new_n988), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n985), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1001), .B1(new_n985), .B2(new_n1000), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n1002), .A2(new_n1003), .ZN(G72));
  NAND2_X1  g818(.A1(G472), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT63), .Z(new_n1006));
  OAI21_X1  g820(.A(new_n1006), .B1(new_n997), .B2(new_n897), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1007), .A2(new_n194), .A3(new_n314), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n305), .B1(new_n395), .B2(new_n194), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n1006), .B(new_n1009), .C1(new_n892), .C2(new_n904), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1006), .B1(new_n981), .B2(new_n897), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n314), .A2(new_n194), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n921), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n1008), .A2(new_n1010), .A3(new_n1013), .ZN(G57));
endmodule


