

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779;

  INV_X1 U374 ( .A(n655), .ZN(n453) );
  NOR2_X1 U375 ( .A1(G953), .A2(G237), .ZN(n514) );
  XNOR2_X1 U376 ( .A(n411), .B(G119), .ZN(n416) );
  XNOR2_X1 U377 ( .A(n372), .B(n450), .ZN(n682) );
  XNOR2_X1 U378 ( .A(n374), .B(n584), .ZN(n598) );
  INV_X2 U379 ( .A(G953), .ZN(n757) );
  XNOR2_X2 U380 ( .A(n369), .B(n596), .ZN(n389) );
  XNOR2_X1 U381 ( .A(n377), .B(n376), .ZN(n375) );
  XNOR2_X2 U382 ( .A(n554), .B(n513), .ZN(n391) );
  NOR2_X2 U383 ( .A1(n738), .A2(n741), .ZN(n409) );
  XNOR2_X1 U384 ( .A(n378), .B(KEYINPUT4), .ZN(n377) );
  XNOR2_X2 U385 ( .A(n502), .B(n713), .ZN(n530) );
  INV_X2 U386 ( .A(G137), .ZN(n378) );
  AND2_X1 U387 ( .A1(n379), .A2(n652), .ZN(n407) );
  AND2_X1 U388 ( .A1(n384), .A2(n383), .ZN(n382) );
  XNOR2_X1 U389 ( .A(n619), .B(n618), .ZN(n717) );
  XNOR2_X1 U390 ( .A(n455), .B(KEYINPUT110), .ZN(n738) );
  NOR2_X1 U391 ( .A1(n432), .A2(n431), .ZN(n430) );
  NAND2_X1 U392 ( .A1(n722), .A2(n604), .ZN(n727) );
  XNOR2_X1 U393 ( .A(n725), .B(KEYINPUT105), .ZN(n559) );
  XNOR2_X1 U394 ( .A(G131), .B(KEYINPUT68), .ZN(n376) );
  OR2_X1 U395 ( .A1(n435), .A2(n436), .ZN(n511) );
  XNOR2_X2 U396 ( .A(n650), .B(n649), .ZN(n655) );
  NAND2_X1 U397 ( .A1(n475), .A2(G953), .ZN(n600) );
  INV_X1 U398 ( .A(G237), .ZN(n506) );
  XNOR2_X1 U399 ( .A(n599), .B(KEYINPUT82), .ZN(n769) );
  OR2_X1 U400 ( .A1(n673), .A2(G902), .ZN(n447) );
  AND2_X1 U401 ( .A1(n739), .A2(KEYINPUT88), .ZN(n434) );
  XNOR2_X1 U402 ( .A(n600), .B(KEYINPUT107), .ZN(n443) );
  NAND2_X1 U403 ( .A1(n438), .A2(n437), .ZN(n436) );
  NAND2_X1 U404 ( .A1(n676), .A2(n454), .ZN(n438) );
  INV_X1 U405 ( .A(n553), .ZN(n448) );
  NAND2_X1 U406 ( .A1(n740), .A2(n739), .ZN(n455) );
  NOR2_X1 U407 ( .A1(n676), .A2(n362), .ZN(n435) );
  AND2_X1 U408 ( .A1(n435), .A2(n434), .ZN(n431) );
  NAND2_X1 U409 ( .A1(n354), .A2(n424), .ZN(n432) );
  AND2_X1 U410 ( .A1(n425), .A2(n433), .ZN(n424) );
  OR2_X1 U411 ( .A1(n739), .A2(KEYINPUT88), .ZN(n433) );
  NOR2_X1 U412 ( .A1(n436), .A2(KEYINPUT88), .ZN(n428) );
  AND2_X1 U413 ( .A1(n385), .A2(n623), .ZN(n384) );
  XNOR2_X1 U414 ( .A(n493), .B(n492), .ZN(n557) );
  XNOR2_X1 U415 ( .A(n406), .B(n603), .ZN(n620) );
  NAND2_X1 U416 ( .A1(n391), .A2(n353), .ZN(n406) );
  XNOR2_X1 U417 ( .A(n463), .B(n462), .ZN(n402) );
  XNOR2_X1 U418 ( .A(G107), .B(KEYINPUT103), .ZN(n533) );
  XOR2_X1 U419 ( .A(KEYINPUT104), .B(KEYINPUT9), .Z(n534) );
  XNOR2_X1 U420 ( .A(G116), .B(G122), .ZN(n536) );
  INV_X1 U421 ( .A(G146), .ZN(n451) );
  XOR2_X1 U422 ( .A(G101), .B(G140), .Z(n489) );
  XNOR2_X1 U423 ( .A(n405), .B(KEYINPUT73), .ZN(n719) );
  NAND2_X1 U424 ( .A1(n583), .A2(n582), .ZN(n374) );
  BUF_X1 U425 ( .A(n722), .Z(n403) );
  NAND2_X1 U426 ( .A1(n664), .A2(n631), .ZN(n546) );
  INV_X1 U427 ( .A(n434), .ZN(n426) );
  NAND2_X1 U428 ( .A1(n454), .A2(n652), .ZN(n437) );
  XNOR2_X1 U429 ( .A(KEYINPUT15), .B(G902), .ZN(n651) );
  NOR2_X1 U430 ( .A1(n426), .A2(n509), .ZN(n423) );
  OR2_X1 U431 ( .A1(n437), .A2(n426), .ZN(n425) );
  XOR2_X1 U432 ( .A(G110), .B(G137), .Z(n459) );
  XNOR2_X1 U433 ( .A(G119), .B(G128), .ZN(n458) );
  XNOR2_X1 U434 ( .A(KEYINPUT94), .B(KEYINPUT24), .ZN(n460) );
  XOR2_X1 U435 ( .A(KEYINPUT23), .B(KEYINPUT81), .Z(n461) );
  XOR2_X1 U436 ( .A(G131), .B(KEYINPUT12), .Z(n516) );
  XNOR2_X1 U437 ( .A(G113), .B(G143), .ZN(n521) );
  XOR2_X1 U438 ( .A(G104), .B(G122), .Z(n522) );
  XNOR2_X1 U439 ( .A(KEYINPUT101), .B(KEYINPUT100), .ZN(n517) );
  XOR2_X1 U440 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n518) );
  NAND2_X1 U441 ( .A1(n655), .A2(n422), .ZN(n379) );
  INV_X1 U442 ( .A(n651), .ZN(n652) );
  XNOR2_X1 U443 ( .A(KEYINPUT76), .B(KEYINPUT4), .ZN(n501) );
  XNOR2_X1 U444 ( .A(n371), .B(n588), .ZN(n370) );
  XNOR2_X1 U445 ( .A(n439), .B(n361), .ZN(n476) );
  XNOR2_X1 U446 ( .A(KEYINPUT71), .B(KEYINPUT14), .ZN(n439) );
  INV_X1 U447 ( .A(KEYINPUT38), .ZN(n446) );
  XNOR2_X1 U448 ( .A(n401), .B(KEYINPUT72), .ZN(n625) );
  NOR2_X1 U449 ( .A1(n726), .A2(n727), .ZN(n401) );
  XNOR2_X1 U450 ( .A(n441), .B(n440), .ZN(n478) );
  INV_X1 U451 ( .A(KEYINPUT108), .ZN(n440) );
  XOR2_X1 U452 ( .A(KEYINPUT5), .B(KEYINPUT98), .Z(n484) );
  XNOR2_X1 U453 ( .A(n496), .B(n495), .ZN(n414) );
  XNOR2_X1 U454 ( .A(KEYINPUT16), .B(G122), .ZN(n495) );
  AND2_X1 U455 ( .A1(n444), .A2(n494), .ZN(n579) );
  XNOR2_X1 U456 ( .A(n487), .B(KEYINPUT28), .ZN(n444) );
  AND2_X1 U457 ( .A1(n559), .A2(n448), .ZN(n487) );
  INV_X1 U458 ( .A(KEYINPUT41), .ZN(n408) );
  NAND2_X1 U459 ( .A1(n430), .A2(n427), .ZN(n554) );
  NAND2_X1 U460 ( .A1(n429), .A2(n428), .ZN(n427) );
  INV_X1 U461 ( .A(n435), .ZN(n429) );
  XNOR2_X1 U462 ( .A(n387), .B(KEYINPUT35), .ZN(n642) );
  NAND2_X1 U463 ( .A1(n382), .A2(n380), .ZN(n387) );
  NAND2_X1 U464 ( .A1(n381), .A2(KEYINPUT34), .ZN(n380) );
  XNOR2_X1 U465 ( .A(n410), .B(n560), .ZN(n583) );
  BUF_X1 U466 ( .A(n557), .Z(n627) );
  BUF_X1 U467 ( .A(n725), .Z(n404) );
  XNOR2_X1 U468 ( .A(n539), .B(n538), .ZN(n658) );
  XNOR2_X1 U469 ( .A(n496), .B(n490), .ZN(n491) );
  NAND2_X1 U470 ( .A1(n453), .A2(n420), .ZN(n419) );
  INV_X1 U471 ( .A(G134), .ZN(n713) );
  XNOR2_X1 U472 ( .A(n373), .B(KEYINPUT40), .ZN(n388) );
  BUF_X1 U473 ( .A(n642), .Z(n693) );
  AND2_X1 U474 ( .A1(n612), .A2(n611), .ZN(n445) );
  INV_X1 U475 ( .A(n572), .ZN(n664) );
  INV_X1 U476 ( .A(KEYINPUT122), .ZN(n399) );
  INV_X1 U477 ( .A(KEYINPUT60), .ZN(n397) );
  INV_X1 U478 ( .A(KEYINPUT56), .ZN(n394) );
  OR2_X1 U479 ( .A1(n602), .A2(n601), .ZN(n353) );
  NAND2_X1 U480 ( .A1(n676), .A2(n423), .ZN(n354) );
  XOR2_X1 U481 ( .A(n484), .B(n483), .Z(n355) );
  INV_X1 U482 ( .A(n509), .ZN(n454) );
  AND2_X1 U483 ( .A1(n609), .A2(n449), .ZN(n356) );
  AND2_X1 U484 ( .A1(n630), .A2(n621), .ZN(n357) );
  AND2_X1 U485 ( .A1(n638), .A2(n637), .ZN(n358) );
  AND2_X1 U486 ( .A1(n419), .A2(n422), .ZN(n359) );
  XOR2_X1 U487 ( .A(n473), .B(n472), .Z(n360) );
  AND2_X1 U488 ( .A1(G234), .A2(G237), .ZN(n361) );
  OR2_X1 U489 ( .A1(n454), .A2(n652), .ZN(n362) );
  AND2_X1 U490 ( .A1(n714), .A2(KEYINPUT2), .ZN(n363) );
  XOR2_X1 U491 ( .A(n689), .B(n688), .Z(n364) );
  XOR2_X1 U492 ( .A(n676), .B(n678), .Z(n365) );
  XOR2_X1 U493 ( .A(n682), .B(n681), .Z(n366) );
  XNOR2_X1 U494 ( .A(KEYINPUT121), .B(n673), .ZN(n367) );
  XNOR2_X1 U495 ( .A(KEYINPUT112), .B(KEYINPUT63), .ZN(n368) );
  NAND2_X1 U496 ( .A1(n370), .A2(n666), .ZN(n369) );
  NAND2_X1 U497 ( .A1(n587), .A2(n457), .ZN(n371) );
  XNOR2_X1 U498 ( .A(n372), .B(n491), .ZN(n696) );
  XNOR2_X2 U499 ( .A(n772), .B(n451), .ZN(n372) );
  NAND2_X1 U500 ( .A1(n598), .A2(n701), .ZN(n373) );
  XNOR2_X2 U501 ( .A(n530), .B(n375), .ZN(n772) );
  XNOR2_X2 U502 ( .A(G143), .B(G128), .ZN(n502) );
  INV_X1 U503 ( .A(n717), .ZN(n381) );
  NAND2_X1 U504 ( .A1(n717), .A2(n357), .ZN(n383) );
  NAND2_X1 U505 ( .A1(n386), .A2(KEYINPUT34), .ZN(n385) );
  INV_X1 U506 ( .A(n630), .ZN(n386) );
  NAND2_X1 U507 ( .A1(n388), .A2(n671), .ZN(n586) );
  XNOR2_X1 U508 ( .A(n388), .B(G131), .ZN(G33) );
  NAND2_X1 U509 ( .A1(n389), .A2(n714), .ZN(n599) );
  NAND2_X1 U510 ( .A1(n389), .A2(n363), .ZN(n654) );
  XNOR2_X2 U511 ( .A(n414), .B(n390), .ZN(n764) );
  XNOR2_X1 U512 ( .A(n390), .B(n355), .ZN(n450) );
  XNOR2_X2 U513 ( .A(n417), .B(n416), .ZN(n390) );
  NAND2_X1 U514 ( .A1(n579), .A2(n391), .ZN(n572) );
  NAND2_X1 U515 ( .A1(n392), .A2(n445), .ZN(n613) );
  NAND2_X1 U516 ( .A1(n392), .A2(n356), .ZN(n610) );
  NAND2_X1 U517 ( .A1(n392), .A2(n611), .ZN(n633) );
  XNOR2_X2 U518 ( .A(n418), .B(n607), .ZN(n392) );
  XNOR2_X1 U519 ( .A(n393), .B(n640), .ZN(n648) );
  NAND2_X1 U520 ( .A1(n639), .A2(n358), .ZN(n393) );
  XNOR2_X1 U521 ( .A(n395), .B(n394), .ZN(G51) );
  NAND2_X1 U522 ( .A1(n680), .A2(n684), .ZN(n395) );
  XNOR2_X1 U523 ( .A(n396), .B(n368), .ZN(G57) );
  NAND2_X1 U524 ( .A1(n685), .A2(n684), .ZN(n396) );
  XNOR2_X1 U525 ( .A(n398), .B(n397), .ZN(G60) );
  NAND2_X1 U526 ( .A1(n691), .A2(n684), .ZN(n398) );
  XNOR2_X1 U527 ( .A(n400), .B(n399), .ZN(G66) );
  NAND2_X1 U528 ( .A1(n675), .A2(n684), .ZN(n400) );
  XNOR2_X1 U529 ( .A(n409), .B(n408), .ZN(n716) );
  INV_X1 U530 ( .A(KEYINPUT2), .ZN(n422) );
  XNOR2_X1 U531 ( .A(n467), .B(n402), .ZN(n673) );
  NAND2_X1 U532 ( .A1(n656), .A2(n453), .ZN(n405) );
  NAND2_X1 U533 ( .A1(n407), .A2(n421), .ZN(n653) );
  NAND2_X1 U534 ( .A1(n559), .A2(n739), .ZN(n410) );
  XNOR2_X2 U535 ( .A(n557), .B(n556), .ZN(n726) );
  XNOR2_X2 U536 ( .A(G116), .B(KEYINPUT3), .ZN(n411) );
  XNOR2_X2 U537 ( .A(n413), .B(n412), .ZN(n417) );
  XNOR2_X2 U538 ( .A(G101), .B(KEYINPUT69), .ZN(n412) );
  XNOR2_X2 U539 ( .A(KEYINPUT91), .B(G113), .ZN(n413) );
  XNOR2_X2 U540 ( .A(n415), .B(G104), .ZN(n496) );
  XNOR2_X2 U541 ( .A(G110), .B(G107), .ZN(n415) );
  NAND2_X1 U542 ( .A1(n620), .A2(n606), .ZN(n418) );
  NAND2_X1 U543 ( .A1(n769), .A2(n422), .ZN(n421) );
  INV_X1 U544 ( .A(n770), .ZN(n420) );
  NAND2_X1 U545 ( .A1(n443), .A2(n442), .ZN(n441) );
  INV_X1 U546 ( .A(G900), .ZN(n442) );
  INV_X1 U547 ( .A(n511), .ZN(n594) );
  XNOR2_X2 U548 ( .A(n511), .B(n446), .ZN(n740) );
  XNOR2_X2 U549 ( .A(G146), .B(G125), .ZN(n499) );
  XNOR2_X2 U550 ( .A(n447), .B(n360), .ZN(n722) );
  INV_X1 U551 ( .A(n559), .ZN(n449) );
  NAND2_X1 U552 ( .A1(n452), .A2(n672), .ZN(n641) );
  XNOR2_X1 U553 ( .A(n452), .B(G110), .ZN(G12) );
  XNOR2_X2 U554 ( .A(n610), .B(KEYINPUT106), .ZN(n452) );
  NAND2_X1 U555 ( .A1(n453), .A2(n757), .ZN(n763) );
  XNOR2_X2 U556 ( .A(n764), .B(n505), .ZN(n676) );
  XNOR2_X1 U557 ( .A(n659), .B(n658), .ZN(n661) );
  XNOR2_X2 U558 ( .A(n580), .B(KEYINPUT42), .ZN(n671) );
  AND2_X1 U559 ( .A1(n661), .A2(n684), .ZN(G63) );
  AND2_X1 U560 ( .A1(n576), .A2(n575), .ZN(n457) );
  XNOR2_X1 U561 ( .A(n660), .B(KEYINPUT90), .ZN(n699) );
  INV_X1 U562 ( .A(KEYINPUT46), .ZN(n585) );
  INV_X1 U563 ( .A(KEYINPUT65), .ZN(n614) );
  NAND2_X1 U564 ( .A1(n625), .A2(n616), .ZN(n619) );
  INV_X1 U565 ( .A(KEYINPUT75), .ZN(n470) );
  XNOR2_X1 U566 ( .A(n471), .B(n470), .ZN(n472) );
  BUF_X1 U567 ( .A(n686), .Z(n694) );
  INV_X1 U568 ( .A(n699), .ZN(n684) );
  XNOR2_X1 U569 ( .A(n459), .B(n458), .ZN(n463) );
  XNOR2_X1 U570 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U571 ( .A(KEYINPUT10), .B(G140), .ZN(n464) );
  XOR2_X2 U572 ( .A(n499), .B(n464), .Z(n771) );
  NAND2_X1 U573 ( .A1(G234), .A2(n757), .ZN(n465) );
  XOR2_X1 U574 ( .A(KEYINPUT8), .B(n465), .Z(n529) );
  NAND2_X1 U575 ( .A1(G221), .A2(n529), .ZN(n466) );
  XNOR2_X1 U576 ( .A(n771), .B(n466), .ZN(n467) );
  XOR2_X1 U577 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n469) );
  NAND2_X1 U578 ( .A1(G234), .A2(n651), .ZN(n468) );
  XNOR2_X1 U579 ( .A(n469), .B(n468), .ZN(n479) );
  NAND2_X1 U580 ( .A1(n479), .A2(G217), .ZN(n473) );
  XNOR2_X1 U581 ( .A(KEYINPUT25), .B(KEYINPUT96), .ZN(n471) );
  NAND2_X1 U582 ( .A1(G902), .A2(n476), .ZN(n474) );
  XNOR2_X1 U583 ( .A(KEYINPUT93), .B(n474), .ZN(n475) );
  NAND2_X1 U584 ( .A1(G952), .A2(n476), .ZN(n750) );
  NOR2_X1 U585 ( .A1(G953), .A2(n750), .ZN(n477) );
  XNOR2_X1 U586 ( .A(n477), .B(KEYINPUT92), .ZN(n601) );
  NOR2_X1 U587 ( .A1(n478), .A2(n601), .ZN(n562) );
  NOR2_X1 U588 ( .A1(n722), .A2(n562), .ZN(n482) );
  NAND2_X1 U589 ( .A1(n479), .A2(G221), .ZN(n481) );
  INV_X1 U590 ( .A(KEYINPUT21), .ZN(n480) );
  XNOR2_X1 U591 ( .A(n481), .B(n480), .ZN(n721) );
  NAND2_X1 U592 ( .A1(n482), .A2(n721), .ZN(n553) );
  NAND2_X1 U593 ( .A1(n514), .A2(G210), .ZN(n483) );
  INV_X1 U594 ( .A(G902), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n682), .A2(n540), .ZN(n486) );
  INV_X1 U596 ( .A(G472), .ZN(n485) );
  XNOR2_X2 U597 ( .A(n486), .B(n485), .ZN(n725) );
  NAND2_X1 U598 ( .A1(G227), .A2(n757), .ZN(n488) );
  XNOR2_X1 U599 ( .A(n489), .B(n488), .ZN(n490) );
  NAND2_X1 U600 ( .A1(n696), .A2(n540), .ZN(n493) );
  INV_X1 U601 ( .A(G469), .ZN(n492) );
  INV_X1 U602 ( .A(n627), .ZN(n494) );
  XNOR2_X1 U603 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n498) );
  NAND2_X1 U604 ( .A1(n757), .A2(G224), .ZN(n497) );
  XNOR2_X1 U605 ( .A(n498), .B(n497), .ZN(n500) );
  XNOR2_X1 U606 ( .A(n500), .B(n499), .ZN(n504) );
  XNOR2_X1 U607 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U608 ( .A(n504), .B(n503), .ZN(n505) );
  NAND2_X1 U609 ( .A1(n540), .A2(n506), .ZN(n510) );
  NAND2_X1 U610 ( .A1(n510), .A2(G210), .ZN(n508) );
  INV_X1 U611 ( .A(KEYINPUT77), .ZN(n507) );
  XNOR2_X1 U612 ( .A(n508), .B(n507), .ZN(n509) );
  NAND2_X1 U613 ( .A1(n510), .A2(G214), .ZN(n739) );
  XNOR2_X1 U614 ( .A(KEYINPUT74), .B(KEYINPUT19), .ZN(n512) );
  XNOR2_X1 U615 ( .A(n512), .B(KEYINPUT67), .ZN(n513) );
  XNOR2_X1 U616 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n527) );
  NAND2_X1 U617 ( .A1(G214), .A2(n514), .ZN(n515) );
  XNOR2_X1 U618 ( .A(n516), .B(n515), .ZN(n520) );
  XNOR2_X1 U619 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U620 ( .A(n520), .B(n519), .Z(n525) );
  XNOR2_X1 U621 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U622 ( .A(n771), .B(n523), .ZN(n524) );
  XNOR2_X1 U623 ( .A(n525), .B(n524), .ZN(n689) );
  NOR2_X1 U624 ( .A1(G902), .A2(n689), .ZN(n526) );
  XNOR2_X1 U625 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U626 ( .A(n528), .B(G475), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n529), .A2(G217), .ZN(n532) );
  INV_X1 U628 ( .A(n530), .ZN(n531) );
  XNOR2_X1 U629 ( .A(n532), .B(n531), .ZN(n539) );
  XNOR2_X1 U630 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U631 ( .A(n535), .B(KEYINPUT7), .Z(n537) );
  XNOR2_X1 U632 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U633 ( .A1(n658), .A2(n540), .ZN(n542) );
  INV_X1 U634 ( .A(G478), .ZN(n541) );
  XNOR2_X1 U635 ( .A(n542), .B(n541), .ZN(n577) );
  AND2_X1 U636 ( .A1(n564), .A2(n577), .ZN(n701) );
  INV_X1 U637 ( .A(n701), .ZN(n543) );
  INV_X1 U638 ( .A(n564), .ZN(n578) );
  INV_X1 U639 ( .A(n577), .ZN(n565) );
  NAND2_X1 U640 ( .A1(n578), .A2(n565), .ZN(n597) );
  NAND2_X1 U641 ( .A1(n543), .A2(n597), .ZN(n631) );
  NOR2_X1 U642 ( .A1(KEYINPUT79), .A2(KEYINPUT47), .ZN(n544) );
  AND2_X1 U643 ( .A1(n544), .A2(KEYINPUT80), .ZN(n545) );
  NAND2_X1 U644 ( .A1(n546), .A2(n545), .ZN(n551) );
  INV_X1 U645 ( .A(KEYINPUT79), .ZN(n571) );
  NAND2_X1 U646 ( .A1(n572), .A2(n571), .ZN(n549) );
  INV_X1 U647 ( .A(n631), .ZN(n737) );
  NAND2_X1 U648 ( .A1(n737), .A2(KEYINPUT80), .ZN(n547) );
  AND2_X1 U649 ( .A1(n547), .A2(KEYINPUT47), .ZN(n548) );
  NAND2_X1 U650 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U651 ( .A1(n551), .A2(n550), .ZN(n576) );
  XNOR2_X1 U652 ( .A(n725), .B(KEYINPUT6), .ZN(n616) );
  NAND2_X1 U653 ( .A1(n616), .A2(n701), .ZN(n552) );
  NOR2_X1 U654 ( .A1(n553), .A2(n552), .ZN(n589) );
  AND2_X1 U655 ( .A1(n554), .A2(n589), .ZN(n555) );
  XNOR2_X1 U656 ( .A(n555), .B(KEYINPUT36), .ZN(n558) );
  XNOR2_X1 U657 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n556) );
  INV_X1 U658 ( .A(n726), .ZN(n608) );
  NAND2_X1 U659 ( .A1(n558), .A2(n608), .ZN(n711) );
  INV_X1 U660 ( .A(KEYINPUT30), .ZN(n560) );
  INV_X1 U661 ( .A(KEYINPUT97), .ZN(n561) );
  XNOR2_X1 U662 ( .A(n721), .B(n561), .ZN(n604) );
  OR2_X2 U663 ( .A1(n562), .A2(n727), .ZN(n563) );
  NOR2_X2 U664 ( .A1(n563), .A2(n627), .ZN(n581) );
  AND2_X1 U665 ( .A1(n583), .A2(n581), .ZN(n567) );
  NAND2_X1 U666 ( .A1(n565), .A2(n564), .ZN(n622) );
  NOR2_X1 U667 ( .A1(n622), .A2(n594), .ZN(n566) );
  NAND2_X1 U668 ( .A1(n567), .A2(n566), .ZN(n709) );
  INV_X1 U669 ( .A(KEYINPUT80), .ZN(n568) );
  NAND2_X1 U670 ( .A1(n631), .A2(n568), .ZN(n569) );
  AND2_X1 U671 ( .A1(n709), .A2(n569), .ZN(n570) );
  NAND2_X1 U672 ( .A1(n711), .A2(n570), .ZN(n574) );
  NOR2_X1 U673 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U674 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U675 ( .A1(n578), .A2(n577), .ZN(n741) );
  NAND2_X1 U676 ( .A1(n579), .A2(n716), .ZN(n580) );
  AND2_X1 U677 ( .A1(n581), .A2(n740), .ZN(n582) );
  XNOR2_X1 U678 ( .A(KEYINPUT70), .B(KEYINPUT39), .ZN(n584) );
  XNOR2_X1 U679 ( .A(n586), .B(n585), .ZN(n587) );
  INV_X1 U680 ( .A(KEYINPUT48), .ZN(n588) );
  NAND2_X1 U681 ( .A1(n589), .A2(n739), .ZN(n590) );
  XOR2_X1 U682 ( .A(KEYINPUT109), .B(n590), .Z(n591) );
  NOR2_X1 U683 ( .A1(n591), .A2(n608), .ZN(n593) );
  INV_X1 U684 ( .A(KEYINPUT43), .ZN(n592) );
  XNOR2_X1 U685 ( .A(n593), .B(n592), .ZN(n595) );
  NAND2_X1 U686 ( .A1(n595), .A2(n594), .ZN(n666) );
  INV_X1 U687 ( .A(KEYINPUT84), .ZN(n596) );
  INV_X1 U688 ( .A(n597), .ZN(n703) );
  NAND2_X1 U689 ( .A1(n598), .A2(n703), .ZN(n714) );
  NOR2_X1 U690 ( .A1(n600), .A2(G898), .ZN(n602) );
  INV_X1 U691 ( .A(KEYINPUT0), .ZN(n603) );
  INV_X1 U692 ( .A(n604), .ZN(n605) );
  NOR2_X1 U693 ( .A1(n741), .A2(n605), .ZN(n606) );
  INV_X1 U694 ( .A(KEYINPUT22), .ZN(n607) );
  NOR2_X1 U695 ( .A1(n403), .A2(n608), .ZN(n609) );
  INV_X1 U696 ( .A(n616), .ZN(n611) );
  NOR2_X1 U697 ( .A1(n403), .A2(n726), .ZN(n612) );
  XNOR2_X2 U698 ( .A(n613), .B(KEYINPUT32), .ZN(n672) );
  NAND2_X1 U699 ( .A1(n641), .A2(KEYINPUT44), .ZN(n615) );
  XNOR2_X1 U700 ( .A(n615), .B(n614), .ZN(n639) );
  INV_X1 U701 ( .A(KEYINPUT89), .ZN(n617) );
  XNOR2_X1 U702 ( .A(n617), .B(KEYINPUT33), .ZN(n618) );
  BUF_X2 U703 ( .A(n620), .Z(n630) );
  INV_X1 U704 ( .A(KEYINPUT34), .ZN(n621) );
  INV_X1 U705 ( .A(n622), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n642), .A2(KEYINPUT44), .ZN(n638) );
  INV_X1 U707 ( .A(n404), .ZN(n624) );
  AND2_X1 U708 ( .A1(n625), .A2(n624), .ZN(n732) );
  NAND2_X1 U709 ( .A1(n630), .A2(n732), .ZN(n626) );
  XNOR2_X1 U710 ( .A(n626), .B(KEYINPUT31), .ZN(n668) );
  NOR2_X1 U711 ( .A1(n627), .A2(n727), .ZN(n628) );
  AND2_X1 U712 ( .A1(n404), .A2(n628), .ZN(n629) );
  AND2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n704) );
  OR2_X1 U714 ( .A1(n668), .A2(n704), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n636) );
  XNOR2_X1 U716 ( .A(n633), .B(KEYINPUT85), .ZN(n635) );
  AND2_X1 U717 ( .A1(n403), .A2(n726), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n635), .A2(n634), .ZN(n670) );
  AND2_X1 U719 ( .A1(n636), .A2(n670), .ZN(n637) );
  INV_X1 U720 ( .A(KEYINPUT86), .ZN(n640) );
  XNOR2_X1 U721 ( .A(n641), .B(KEYINPUT87), .ZN(n646) );
  INV_X1 U722 ( .A(n693), .ZN(n644) );
  INV_X1 U723 ( .A(KEYINPUT44), .ZN(n643) );
  AND2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n648), .A2(n647), .ZN(n650) );
  INV_X1 U727 ( .A(KEYINPUT45), .ZN(n649) );
  XNOR2_X1 U728 ( .A(n653), .B(KEYINPUT64), .ZN(n657) );
  XNOR2_X1 U729 ( .A(n654), .B(KEYINPUT83), .ZN(n656) );
  NOR2_X2 U730 ( .A1(n657), .A2(n719), .ZN(n686) );
  NAND2_X1 U731 ( .A1(n694), .A2(G478), .ZN(n659) );
  NOR2_X1 U732 ( .A1(n757), .A2(G952), .ZN(n660) );
  NAND2_X1 U733 ( .A1(n664), .A2(n703), .ZN(n663) );
  XOR2_X1 U734 ( .A(G128), .B(KEYINPUT29), .Z(n662) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(G30) );
  NAND2_X1 U736 ( .A1(n664), .A2(n701), .ZN(n665) );
  XNOR2_X1 U737 ( .A(n665), .B(G146), .ZN(G48) );
  XNOR2_X1 U738 ( .A(n666), .B(G140), .ZN(G42) );
  NAND2_X1 U739 ( .A1(n668), .A2(n701), .ZN(n667) );
  XNOR2_X1 U740 ( .A(n667), .B(G113), .ZN(G15) );
  NAND2_X1 U741 ( .A1(n668), .A2(n703), .ZN(n669) );
  XNOR2_X1 U742 ( .A(n669), .B(G116), .ZN(G18) );
  XNOR2_X1 U743 ( .A(n670), .B(G101), .ZN(G3) );
  XNOR2_X1 U744 ( .A(n671), .B(G137), .ZN(G39) );
  XNOR2_X1 U745 ( .A(n672), .B(G119), .ZN(G21) );
  NAND2_X1 U746 ( .A1(n686), .A2(G217), .ZN(n674) );
  XNOR2_X1 U747 ( .A(n674), .B(n367), .ZN(n675) );
  NAND2_X1 U748 ( .A1(n686), .A2(G210), .ZN(n679) );
  XNOR2_X1 U749 ( .A(KEYINPUT78), .B(KEYINPUT54), .ZN(n677) );
  XOR2_X1 U750 ( .A(n677), .B(KEYINPUT55), .Z(n678) );
  XNOR2_X1 U751 ( .A(n679), .B(n365), .ZN(n680) );
  NAND2_X1 U752 ( .A1(n686), .A2(G472), .ZN(n683) );
  XNOR2_X1 U753 ( .A(KEYINPUT111), .B(KEYINPUT62), .ZN(n681) );
  XNOR2_X1 U754 ( .A(n683), .B(n366), .ZN(n685) );
  NAND2_X1 U755 ( .A1(n686), .A2(G475), .ZN(n690) );
  XNOR2_X1 U756 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n687) );
  XNOR2_X1 U757 ( .A(n687), .B(KEYINPUT59), .ZN(n688) );
  XNOR2_X1 U758 ( .A(n690), .B(n364), .ZN(n691) );
  XNOR2_X1 U759 ( .A(G122), .B(KEYINPUT127), .ZN(n692) );
  XNOR2_X1 U760 ( .A(n693), .B(n692), .ZN(G24) );
  NAND2_X1 U761 ( .A1(n694), .A2(G469), .ZN(n698) );
  XNOR2_X1 U762 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n695) );
  XNOR2_X1 U763 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U764 ( .A(n698), .B(n697), .ZN(n700) );
  NOR2_X1 U765 ( .A1(n700), .A2(n699), .ZN(G54) );
  NAND2_X1 U766 ( .A1(n704), .A2(n701), .ZN(n702) );
  XNOR2_X1 U767 ( .A(n702), .B(G104), .ZN(G6) );
  XOR2_X1 U768 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n706) );
  NAND2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U770 ( .A(n706), .B(n705), .ZN(n708) );
  XOR2_X1 U771 ( .A(G107), .B(KEYINPUT113), .Z(n707) );
  XNOR2_X1 U772 ( .A(n708), .B(n707), .ZN(G9) );
  XNOR2_X1 U773 ( .A(G143), .B(n709), .ZN(G45) );
  XOR2_X1 U774 ( .A(KEYINPUT114), .B(KEYINPUT37), .Z(n710) );
  XNOR2_X1 U775 ( .A(n711), .B(n710), .ZN(n712) );
  XNOR2_X1 U776 ( .A(G125), .B(n712), .ZN(G27) );
  XNOR2_X1 U777 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U778 ( .A(n715), .B(KEYINPUT115), .ZN(G36) );
  INV_X1 U779 ( .A(n716), .ZN(n735) );
  NOR2_X1 U780 ( .A1(n735), .A2(n381), .ZN(n718) );
  NOR2_X1 U781 ( .A1(n718), .A2(G953), .ZN(n755) );
  NOR2_X1 U782 ( .A1(n719), .A2(n359), .ZN(n753) );
  XOR2_X1 U783 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n720) );
  XNOR2_X1 U784 ( .A(KEYINPUT116), .B(n720), .ZN(n734) );
  NOR2_X1 U785 ( .A1(n403), .A2(n721), .ZN(n723) );
  XNOR2_X1 U786 ( .A(n723), .B(KEYINPUT49), .ZN(n724) );
  NAND2_X1 U787 ( .A1(n404), .A2(n724), .ZN(n730) );
  NAND2_X1 U788 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U789 ( .A(KEYINPUT50), .B(n728), .Z(n729) );
  NOR2_X1 U790 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U791 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U792 ( .A(n734), .B(n733), .Z(n736) );
  NOR2_X1 U793 ( .A1(n736), .A2(n735), .ZN(n747) );
  NOR2_X1 U794 ( .A1(n738), .A2(n737), .ZN(n744) );
  NOR2_X1 U795 ( .A1(n740), .A2(n739), .ZN(n742) );
  NOR2_X1 U796 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U797 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U798 ( .A1(n745), .A2(n381), .ZN(n746) );
  NOR2_X1 U799 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U800 ( .A(n748), .B(KEYINPUT52), .ZN(n749) );
  NOR2_X1 U801 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U802 ( .A(n751), .B(KEYINPUT118), .ZN(n752) );
  NOR2_X1 U803 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U804 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U805 ( .A(KEYINPUT53), .B(n756), .Z(G75) );
  XOR2_X1 U806 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n759) );
  NAND2_X1 U807 ( .A1(G224), .A2(G953), .ZN(n758) );
  XNOR2_X1 U808 ( .A(n759), .B(n758), .ZN(n760) );
  XNOR2_X1 U809 ( .A(KEYINPUT123), .B(n760), .ZN(n761) );
  NAND2_X1 U810 ( .A1(n761), .A2(G898), .ZN(n762) );
  NAND2_X1 U811 ( .A1(n763), .A2(n762), .ZN(n768) );
  XOR2_X1 U812 ( .A(KEYINPUT125), .B(n764), .Z(n766) );
  NOR2_X1 U813 ( .A1(n757), .A2(G898), .ZN(n765) );
  NOR2_X1 U814 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U815 ( .A(n768), .B(n767), .ZN(G69) );
  BUF_X1 U816 ( .A(n769), .Z(n770) );
  XNOR2_X1 U817 ( .A(n772), .B(n771), .ZN(n774) );
  XNOR2_X1 U818 ( .A(n770), .B(n774), .ZN(n773) );
  NAND2_X1 U819 ( .A1(n773), .A2(n757), .ZN(n779) );
  XNOR2_X1 U820 ( .A(G227), .B(n774), .ZN(n775) );
  NAND2_X1 U821 ( .A1(n775), .A2(G900), .ZN(n776) );
  XNOR2_X1 U822 ( .A(KEYINPUT126), .B(n776), .ZN(n777) );
  NAND2_X1 U823 ( .A1(n777), .A2(G953), .ZN(n778) );
  NAND2_X1 U824 ( .A1(n779), .A2(n778), .ZN(G72) );
endmodule

