

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755;

  OR2_X1 U375 ( .A1(n653), .A2(n618), .ZN(n371) );
  NAND2_X1 U376 ( .A1(n352), .A2(n584), .ZN(n614) );
  NAND2_X1 U377 ( .A1(n581), .A2(n582), .ZN(n352) );
  INV_X1 U378 ( .A(KEYINPUT66), .ZN(n411) );
  XNOR2_X1 U379 ( .A(n411), .B(G101), .ZN(n473) );
  XNOR2_X1 U380 ( .A(G119), .B(G116), .ZN(n449) );
  XNOR2_X1 U381 ( .A(n393), .B(n392), .ZN(n515) );
  INV_X2 U382 ( .A(G953), .ZN(n406) );
  AND2_X4 U383 ( .A1(n619), .A2(n663), .ZN(n652) );
  NOR2_X2 U384 ( .A1(n403), .A2(n516), .ZN(n720) );
  XNOR2_X1 U385 ( .A(n353), .B(KEYINPUT13), .ZN(n516) );
  XNOR2_X1 U386 ( .A(n377), .B(KEYINPUT67), .ZN(n379) );
  XNOR2_X2 U387 ( .A(n533), .B(n494), .ZN(n555) );
  INV_X1 U388 ( .A(n628), .ZN(n567) );
  XNOR2_X1 U389 ( .A(n427), .B(n426), .ZN(n527) );
  INV_X1 U390 ( .A(G131), .ZN(n377) );
  AND2_X1 U391 ( .A1(n365), .A2(KEYINPUT44), .ZN(n581) );
  XNOR2_X1 U392 ( .A(n473), .B(n475), .ZN(n361) );
  XNOR2_X1 U393 ( .A(n478), .B(KEYINPUT77), .ZN(n359) );
  XNOR2_X1 U394 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n472) );
  XNOR2_X1 U395 ( .A(KEYINPUT18), .B(KEYINPUT83), .ZN(n471) );
  NAND2_X1 U396 ( .A1(n372), .A2(n666), .ZN(n586) );
  INV_X1 U397 ( .A(n572), .ZN(n372) );
  XNOR2_X1 U398 ( .A(n356), .B(KEYINPUT0), .ZN(n587) );
  INV_X1 U399 ( .A(KEYINPUT48), .ZN(n540) );
  XNOR2_X1 U400 ( .A(n481), .B(n482), .ZN(n731) );
  XNOR2_X1 U401 ( .A(n476), .B(n394), .ZN(n745) );
  XNOR2_X1 U402 ( .A(KEYINPUT108), .B(KEYINPUT28), .ZN(n490) );
  INV_X1 U403 ( .A(n514), .ZN(n683) );
  XNOR2_X1 U404 ( .A(n455), .B(n416), .ZN(n744) );
  INV_X1 U405 ( .A(KEYINPUT92), .ZN(n416) );
  XNOR2_X1 U406 ( .A(n527), .B(n526), .ZN(n572) );
  AND2_X1 U407 ( .A1(n431), .A2(G221), .ZN(n432) );
  XNOR2_X1 U408 ( .A(n745), .B(n354), .ZN(n401) );
  XNOR2_X1 U409 ( .A(n474), .B(n359), .ZN(n358) );
  XNOR2_X1 U410 ( .A(n511), .B(KEYINPUT39), .ZN(n542) );
  OR2_X2 U411 ( .A1(n587), .A2(n557), .ZN(n560) );
  BUF_X1 U412 ( .A(n572), .Z(n600) );
  XNOR2_X1 U413 ( .A(n580), .B(n366), .ZN(n365) );
  INV_X1 U414 ( .A(KEYINPUT35), .ZN(n366) );
  NOR2_X1 U415 ( .A1(n520), .A2(n495), .ZN(n718) );
  XNOR2_X1 U416 ( .A(n365), .B(G122), .ZN(G24) );
  XOR2_X1 U417 ( .A(G475), .B(n402), .Z(n353) );
  OR2_X2 U418 ( .A1(n507), .A2(n493), .ZN(n533) );
  AND2_X1 U419 ( .A1(n456), .A2(G214), .ZN(n354) );
  NOR2_X1 U420 ( .A1(n514), .A2(n508), .ZN(n355) );
  INV_X1 U421 ( .A(n666), .ZN(n373) );
  NAND2_X1 U422 ( .A1(n555), .A2(n554), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n731), .B(n357), .ZN(n653) );
  XNOR2_X1 U424 ( .A(n360), .B(n358), .ZN(n357) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n477), .B(n476), .ZN(n362) );
  AND2_X2 U427 ( .A1(n363), .A2(n617), .ZN(n662) );
  NAND2_X1 U428 ( .A1(n737), .A2(n616), .ZN(n363) );
  XNOR2_X2 U429 ( .A(n364), .B(KEYINPUT45), .ZN(n737) );
  NAND2_X1 U430 ( .A1(n614), .A2(n613), .ZN(n364) );
  NAND2_X1 U431 ( .A1(n365), .A2(n583), .ZN(n607) );
  OR2_X1 U432 ( .A1(n370), .A2(n367), .ZN(n368) );
  INV_X1 U433 ( .A(n454), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n482), .B(n453), .ZN(n370) );
  NAND2_X1 U435 ( .A1(n369), .A2(n368), .ZN(n460) );
  NAND2_X1 U436 ( .A1(n370), .A2(n367), .ZN(n369) );
  XNOR2_X2 U437 ( .A(n371), .B(n486), .ZN(n507) );
  AND2_X1 U438 ( .A1(n572), .A2(n373), .ZN(n668) );
  NAND2_X1 U439 ( .A1(n647), .A2(n465), .ZN(n427) );
  XNOR2_X2 U440 ( .A(n374), .B(n423), .ZN(n647) );
  NAND2_X1 U441 ( .A1(n376), .A2(n375), .ZN(n374) );
  NAND2_X1 U442 ( .A1(n744), .A2(n454), .ZN(n375) );
  NAND2_X1 U443 ( .A1(n417), .A2(n367), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n564), .B(n563), .ZN(n630) );
  BUF_X1 U445 ( .A(n630), .Z(n631) );
  XNOR2_X1 U446 ( .A(n415), .B(n414), .ZN(n455) );
  XNOR2_X1 U447 ( .A(n414), .B(n384), .ZN(n385) );
  XNOR2_X1 U448 ( .A(n422), .B(n480), .ZN(n423) );
  XOR2_X1 U449 ( .A(G122), .B(G116), .Z(n378) );
  AND2_X1 U450 ( .A1(n509), .A2(n355), .ZN(n380) );
  OR2_X1 U451 ( .A1(n508), .A2(n470), .ZN(n381) );
  NOR2_X1 U452 ( .A1(n755), .A2(n754), .ZN(n525) );
  INV_X1 U453 ( .A(n726), .ZN(n536) );
  XNOR2_X1 U454 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U455 ( .A(n460), .B(n459), .ZN(n637) );
  XNOR2_X1 U456 ( .A(KEYINPUT102), .B(KEYINPUT7), .ZN(n384) );
  XNOR2_X1 U457 ( .A(n541), .B(n540), .ZN(n548) );
  NOR2_X2 U458 ( .A1(n662), .A2(n483), .ZN(n619) );
  XNOR2_X1 U459 ( .A(n447), .B(n446), .ZN(n671) );
  AND2_X1 U460 ( .A1(n542), .A2(n720), .ZN(n513) );
  INV_X1 U461 ( .A(KEYINPUT42), .ZN(n523) );
  INV_X1 U462 ( .A(KEYINPUT60), .ZN(n626) );
  XNOR2_X1 U463 ( .A(n524), .B(n523), .ZN(n754) );
  XOR2_X1 U464 ( .A(KEYINPUT101), .B(KEYINPUT9), .Z(n383) );
  XNOR2_X1 U465 ( .A(G107), .B(KEYINPUT103), .ZN(n382) );
  XNOR2_X1 U466 ( .A(n383), .B(n382), .ZN(n386) );
  XNOR2_X2 U467 ( .A(G143), .B(G128), .ZN(n478) );
  XNOR2_X1 U468 ( .A(n478), .B(G134), .ZN(n414) );
  XOR2_X1 U469 ( .A(n386), .B(n385), .Z(n391) );
  NAND2_X1 U470 ( .A1(G234), .A2(n406), .ZN(n387) );
  XOR2_X1 U471 ( .A(KEYINPUT8), .B(n387), .Z(n431) );
  NAND2_X1 U472 ( .A1(G217), .A2(n431), .ZN(n389) );
  XNOR2_X1 U473 ( .A(KEYINPUT100), .B(n378), .ZN(n388) );
  XNOR2_X1 U474 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U475 ( .A(n391), .B(n390), .ZN(n643) );
  INV_X1 U476 ( .A(G902), .ZN(n465) );
  NAND2_X1 U477 ( .A1(n643), .A2(n465), .ZN(n393) );
  XOR2_X1 U478 ( .A(KEYINPUT104), .B(G478), .Z(n392) );
  INV_X1 U479 ( .A(n515), .ZN(n403) );
  XNOR2_X1 U480 ( .A(G146), .B(G125), .ZN(n476) );
  XNOR2_X1 U481 ( .A(G140), .B(KEYINPUT10), .ZN(n394) );
  NOR2_X1 U482 ( .A1(G953), .A2(G237), .ZN(n456) );
  XNOR2_X1 U483 ( .A(G113), .B(G122), .ZN(n395) );
  XNOR2_X1 U484 ( .A(n379), .B(n395), .ZN(n399) );
  XOR2_X1 U485 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n397) );
  XNOR2_X1 U486 ( .A(G104), .B(G143), .ZN(n396) );
  XNOR2_X1 U487 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U488 ( .A(n399), .B(n398), .Z(n400) );
  XNOR2_X1 U489 ( .A(n401), .B(n400), .ZN(n621) );
  NOR2_X1 U490 ( .A1(n621), .A2(G902), .ZN(n402) );
  INV_X1 U491 ( .A(n516), .ZN(n404) );
  NOR2_X2 U492 ( .A1(n404), .A2(n515), .ZN(n723) );
  OR2_X1 U493 ( .A1(n720), .A2(n723), .ZN(n405) );
  XNOR2_X1 U494 ( .A(KEYINPUT105), .B(n405), .ZN(n687) );
  NAND2_X1 U495 ( .A1(KEYINPUT47), .A2(n687), .ZN(n504) );
  NOR2_X1 U496 ( .A1(G900), .A2(n406), .ZN(n407) );
  NAND2_X1 U497 ( .A1(G902), .A2(n407), .ZN(n408) );
  NAND2_X1 U498 ( .A1(n406), .A2(G952), .ZN(n551) );
  NAND2_X1 U499 ( .A1(n408), .A2(n551), .ZN(n410) );
  NAND2_X1 U500 ( .A1(G237), .A2(G234), .ZN(n409) );
  XNOR2_X1 U501 ( .A(n409), .B(KEYINPUT14), .ZN(n697) );
  NAND2_X1 U502 ( .A1(n410), .A2(n697), .ZN(n508) );
  INV_X1 U503 ( .A(n473), .ZN(n412) );
  XNOR2_X1 U504 ( .A(G146), .B(n412), .ZN(n454) );
  XOR2_X1 U505 ( .A(G137), .B(KEYINPUT4), .Z(n413) );
  XNOR2_X1 U506 ( .A(n379), .B(n413), .ZN(n415) );
  INV_X1 U507 ( .A(n744), .ZN(n417) );
  XOR2_X1 U508 ( .A(G140), .B(KEYINPUT76), .Z(n419) );
  NAND2_X1 U509 ( .A1(G227), .A2(n406), .ZN(n418) );
  XNOR2_X1 U510 ( .A(n419), .B(n418), .ZN(n422) );
  XNOR2_X1 U511 ( .A(G110), .B(G107), .ZN(n421) );
  INV_X1 U512 ( .A(G104), .ZN(n420) );
  XNOR2_X1 U513 ( .A(n421), .B(n420), .ZN(n480) );
  XNOR2_X1 U514 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n425) );
  INV_X1 U515 ( .A(G469), .ZN(n424) );
  XNOR2_X1 U516 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U517 ( .A(KEYINPUT15), .B(G902), .ZN(n483) );
  NAND2_X1 U518 ( .A1(G234), .A2(n483), .ZN(n428) );
  XNOR2_X1 U519 ( .A(KEYINPUT20), .B(n428), .ZN(n441) );
  AND2_X1 U520 ( .A1(n441), .A2(G221), .ZN(n430) );
  INV_X1 U521 ( .A(KEYINPUT21), .ZN(n429) );
  XNOR2_X1 U522 ( .A(n430), .B(n429), .ZN(n672) );
  XNOR2_X1 U523 ( .A(n745), .B(n432), .ZN(n440) );
  XOR2_X1 U524 ( .A(G137), .B(G110), .Z(n434) );
  XNOR2_X1 U525 ( .A(G128), .B(G119), .ZN(n433) );
  XNOR2_X1 U526 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U527 ( .A(KEYINPUT93), .B(KEYINPUT23), .Z(n436) );
  XNOR2_X1 U528 ( .A(KEYINPUT24), .B(KEYINPUT94), .ZN(n435) );
  XNOR2_X1 U529 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U530 ( .A(n438), .B(n437), .Z(n439) );
  XNOR2_X1 U531 ( .A(n440), .B(n439), .ZN(n632) );
  NAND2_X1 U532 ( .A1(n632), .A2(n465), .ZN(n447) );
  XOR2_X1 U533 ( .A(KEYINPUT25), .B(KEYINPUT75), .Z(n443) );
  NAND2_X1 U534 ( .A1(n441), .A2(G217), .ZN(n442) );
  XNOR2_X1 U535 ( .A(n443), .B(n442), .ZN(n445) );
  INV_X1 U536 ( .A(KEYINPUT95), .ZN(n444) );
  XNOR2_X1 U537 ( .A(n445), .B(n444), .ZN(n446) );
  NOR2_X1 U538 ( .A1(n672), .A2(n671), .ZN(n666) );
  NAND2_X1 U539 ( .A1(n527), .A2(n666), .ZN(n448) );
  XNOR2_X1 U540 ( .A(n448), .B(KEYINPUT96), .ZN(n591) );
  XNOR2_X1 U541 ( .A(KEYINPUT107), .B(KEYINPUT30), .ZN(n469) );
  XNOR2_X1 U542 ( .A(n449), .B(KEYINPUT3), .ZN(n451) );
  XNOR2_X1 U543 ( .A(G113), .B(KEYINPUT85), .ZN(n450) );
  XNOR2_X1 U544 ( .A(n451), .B(n450), .ZN(n482) );
  XOR2_X1 U545 ( .A(KEYINPUT73), .B(KEYINPUT5), .Z(n452) );
  XNOR2_X1 U546 ( .A(n452), .B(KEYINPUT97), .ZN(n453) );
  INV_X1 U547 ( .A(n455), .ZN(n458) );
  NAND2_X1 U548 ( .A1(G210), .A2(n456), .ZN(n457) );
  NAND2_X1 U549 ( .A1(n637), .A2(n465), .ZN(n463) );
  INV_X1 U550 ( .A(KEYINPUT98), .ZN(n461) );
  XNOR2_X1 U551 ( .A(n461), .B(G472), .ZN(n462) );
  XNOR2_X1 U552 ( .A(n463), .B(n462), .ZN(n528) );
  INV_X1 U553 ( .A(G237), .ZN(n464) );
  NAND2_X1 U554 ( .A1(n465), .A2(n464), .ZN(n484) );
  NAND2_X1 U555 ( .A1(n484), .A2(G214), .ZN(n467) );
  INV_X1 U556 ( .A(KEYINPUT89), .ZN(n466) );
  XNOR2_X1 U557 ( .A(n467), .B(n466), .ZN(n682) );
  INV_X1 U558 ( .A(n682), .ZN(n493) );
  NOR2_X1 U559 ( .A1(n528), .A2(n493), .ZN(n468) );
  XOR2_X1 U560 ( .A(n469), .B(n468), .Z(n509) );
  NAND2_X1 U561 ( .A1(n510), .A2(n509), .ZN(n470) );
  NOR2_X1 U562 ( .A1(n516), .A2(n515), .ZN(n578) );
  XNOR2_X1 U563 ( .A(n472), .B(n471), .ZN(n474) );
  XNOR2_X1 U564 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n475) );
  NAND2_X1 U565 ( .A1(n406), .A2(G224), .ZN(n477) );
  XNOR2_X1 U566 ( .A(KEYINPUT16), .B(G122), .ZN(n479) );
  XNOR2_X1 U567 ( .A(n480), .B(n479), .ZN(n481) );
  INV_X1 U568 ( .A(n483), .ZN(n618) );
  NAND2_X1 U569 ( .A1(n484), .A2(G210), .ZN(n485) );
  XNOR2_X1 U570 ( .A(n485), .B(KEYINPUT88), .ZN(n486) );
  INV_X1 U571 ( .A(n507), .ZN(n487) );
  NAND2_X1 U572 ( .A1(n578), .A2(n487), .ZN(n488) );
  NOR2_X1 U573 ( .A1(n381), .A2(n488), .ZN(n717) );
  NOR2_X1 U574 ( .A1(n672), .A2(n508), .ZN(n489) );
  NAND2_X1 U575 ( .A1(n671), .A2(n489), .ZN(n530) );
  NOR2_X1 U576 ( .A1(n528), .A2(n530), .ZN(n491) );
  XNOR2_X1 U577 ( .A(n491), .B(n490), .ZN(n492) );
  NAND2_X1 U578 ( .A1(n492), .A2(n527), .ZN(n520) );
  XNOR2_X1 U579 ( .A(KEYINPUT74), .B(KEYINPUT19), .ZN(n494) );
  INV_X1 U580 ( .A(n555), .ZN(n495) );
  INV_X1 U581 ( .A(KEYINPUT47), .ZN(n496) );
  NOR2_X1 U582 ( .A1(n718), .A2(n496), .ZN(n497) );
  XNOR2_X1 U583 ( .A(n497), .B(KEYINPUT79), .ZN(n501) );
  NOR2_X1 U584 ( .A1(n687), .A2(KEYINPUT47), .ZN(n498) );
  XNOR2_X1 U585 ( .A(n498), .B(KEYINPUT72), .ZN(n499) );
  NAND2_X1 U586 ( .A1(n499), .A2(n718), .ZN(n500) );
  NAND2_X1 U587 ( .A1(n501), .A2(n500), .ZN(n502) );
  NOR2_X1 U588 ( .A1(n717), .A2(n502), .ZN(n503) );
  NAND2_X1 U589 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U590 ( .A(n505), .B(KEYINPUT71), .ZN(n539) );
  INV_X1 U591 ( .A(n591), .ZN(n510) );
  INV_X1 U592 ( .A(KEYINPUT38), .ZN(n506) );
  XNOR2_X1 U593 ( .A(n507), .B(n506), .ZN(n514) );
  NAND2_X1 U594 ( .A1(n510), .A2(n380), .ZN(n511) );
  XOR2_X1 U595 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n512) );
  XNOR2_X1 U596 ( .A(n513), .B(n512), .ZN(n755) );
  XOR2_X1 U597 ( .A(KEYINPUT41), .B(KEYINPUT110), .Z(n519) );
  NAND2_X1 U598 ( .A1(n683), .A2(n682), .ZN(n686) );
  INV_X1 U599 ( .A(n686), .ZN(n517) );
  AND2_X1 U600 ( .A1(n516), .A2(n515), .ZN(n681) );
  NAND2_X1 U601 ( .A1(n517), .A2(n681), .ZN(n518) );
  XNOR2_X1 U602 ( .A(n519), .B(n518), .ZN(n699) );
  NOR2_X1 U603 ( .A1(n699), .A2(n520), .ZN(n522) );
  XNOR2_X1 U604 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n521) );
  XNOR2_X1 U605 ( .A(n522), .B(n521), .ZN(n524) );
  XNOR2_X1 U606 ( .A(n525), .B(KEYINPUT46), .ZN(n537) );
  INV_X1 U607 ( .A(KEYINPUT1), .ZN(n526) );
  BUF_X1 U608 ( .A(n528), .Z(n669) );
  INV_X1 U609 ( .A(KEYINPUT6), .ZN(n529) );
  XNOR2_X1 U610 ( .A(n669), .B(n529), .ZN(n598) );
  INV_X1 U611 ( .A(n720), .ZN(n531) );
  NOR2_X1 U612 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U613 ( .A1(n574), .A2(n532), .ZN(n544) );
  NOR2_X1 U614 ( .A1(n544), .A2(n533), .ZN(n534) );
  XOR2_X1 U615 ( .A(KEYINPUT36), .B(n534), .Z(n535) );
  NOR2_X1 U616 ( .A1(n600), .A2(n535), .ZN(n726) );
  AND2_X1 U617 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U618 ( .A1(n539), .A2(n538), .ZN(n541) );
  NAND2_X1 U619 ( .A1(n723), .A2(n542), .ZN(n728) );
  NAND2_X1 U620 ( .A1(n682), .A2(n600), .ZN(n543) );
  NOR2_X1 U621 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U622 ( .A(n545), .B(KEYINPUT43), .Z(n546) );
  NAND2_X1 U623 ( .A1(n546), .A2(n507), .ZN(n729) );
  AND2_X1 U624 ( .A1(n728), .A2(n729), .ZN(n547) );
  NAND2_X1 U625 ( .A1(n548), .A2(n547), .ZN(n747) );
  INV_X1 U626 ( .A(n747), .ZN(n616) );
  NAND2_X1 U627 ( .A1(n616), .A2(KEYINPUT2), .ZN(n549) );
  XNOR2_X1 U628 ( .A(n549), .B(KEYINPUT81), .ZN(n615) );
  XOR2_X1 U629 ( .A(G898), .B(KEYINPUT90), .Z(n736) );
  NAND2_X1 U630 ( .A1(n736), .A2(G953), .ZN(n550) );
  XNOR2_X1 U631 ( .A(n550), .B(KEYINPUT91), .ZN(n732) );
  NAND2_X1 U632 ( .A1(n732), .A2(G902), .ZN(n552) );
  NAND2_X1 U633 ( .A1(n552), .A2(n551), .ZN(n553) );
  AND2_X1 U634 ( .A1(n553), .A2(n697), .ZN(n554) );
  INV_X1 U635 ( .A(n672), .ZN(n556) );
  NAND2_X1 U636 ( .A1(n681), .A2(n556), .ZN(n557) );
  XNOR2_X1 U637 ( .A(KEYINPUT70), .B(KEYINPUT22), .ZN(n558) );
  XNOR2_X1 U638 ( .A(n558), .B(KEYINPUT65), .ZN(n559) );
  XNOR2_X2 U639 ( .A(n560), .B(n559), .ZN(n596) );
  NAND2_X1 U640 ( .A1(n598), .A2(n671), .ZN(n561) );
  NOR2_X1 U641 ( .A1(n600), .A2(n561), .ZN(n562) );
  NAND2_X1 U642 ( .A1(n596), .A2(n562), .ZN(n564) );
  INV_X1 U643 ( .A(KEYINPUT32), .ZN(n563) );
  INV_X1 U644 ( .A(n630), .ZN(n568) );
  AND2_X1 U645 ( .A1(n669), .A2(n671), .ZN(n565) );
  AND2_X1 U646 ( .A1(n600), .A2(n565), .ZN(n566) );
  AND2_X1 U647 ( .A1(n596), .A2(n566), .ZN(n628) );
  NAND2_X1 U648 ( .A1(n568), .A2(n567), .ZN(n570) );
  INV_X1 U649 ( .A(KEYINPUT82), .ZN(n569) );
  XNOR2_X1 U650 ( .A(n570), .B(n569), .ZN(n609) );
  INV_X1 U651 ( .A(n609), .ZN(n571) );
  NAND2_X1 U652 ( .A1(n571), .A2(KEYINPUT64), .ZN(n582) );
  INV_X1 U653 ( .A(n598), .ZN(n574) );
  INV_X1 U654 ( .A(n586), .ZN(n573) );
  NAND2_X1 U655 ( .A1(n574), .A2(n573), .ZN(n576) );
  INV_X1 U656 ( .A(KEYINPUT33), .ZN(n575) );
  XNOR2_X1 U657 ( .A(n576), .B(n575), .ZN(n700) );
  NOR2_X1 U658 ( .A1(n700), .A2(n587), .ZN(n577) );
  XNOR2_X1 U659 ( .A(n577), .B(KEYINPUT34), .ZN(n579) );
  NAND2_X1 U660 ( .A1(n579), .A2(n578), .ZN(n580) );
  INV_X1 U661 ( .A(KEYINPUT44), .ZN(n583) );
  NAND2_X1 U662 ( .A1(n583), .A2(KEYINPUT64), .ZN(n584) );
  NOR2_X1 U663 ( .A1(n586), .A2(n669), .ZN(n677) );
  INV_X1 U664 ( .A(n587), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n677), .A2(n592), .ZN(n589) );
  XOR2_X1 U666 ( .A(KEYINPUT31), .B(KEYINPUT99), .Z(n588) );
  XNOR2_X1 U667 ( .A(n589), .B(n588), .ZN(n724) );
  INV_X1 U668 ( .A(n669), .ZN(n590) );
  NOR2_X1 U669 ( .A1(n591), .A2(n590), .ZN(n593) );
  AND2_X1 U670 ( .A1(n593), .A2(n592), .ZN(n710) );
  OR2_X1 U671 ( .A1(n724), .A2(n710), .ZN(n595) );
  INV_X1 U672 ( .A(n687), .ZN(n594) );
  NAND2_X1 U673 ( .A1(n595), .A2(n594), .ZN(n603) );
  INV_X1 U674 ( .A(n596), .ZN(n602) );
  INV_X1 U675 ( .A(n671), .ZN(n597) );
  AND2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n601) );
  OR2_X1 U678 ( .A1(n602), .A2(n601), .ZN(n629) );
  NAND2_X1 U679 ( .A1(n603), .A2(n629), .ZN(n608) );
  INV_X1 U680 ( .A(KEYINPUT106), .ZN(n604) );
  XNOR2_X1 U681 ( .A(n608), .B(n604), .ZN(n605) );
  AND2_X1 U682 ( .A1(KEYINPUT64), .A2(n605), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n612) );
  XNOR2_X1 U684 ( .A(n608), .B(KEYINPUT106), .ZN(n610) );
  OR2_X2 U685 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n615), .A2(n737), .ZN(n663) );
  INV_X1 U688 ( .A(KEYINPUT2), .ZN(n617) );
  NAND2_X1 U689 ( .A1(n652), .A2(G475), .ZN(n623) );
  XNOR2_X1 U690 ( .A(KEYINPUT84), .B(KEYINPUT59), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U692 ( .A(n623), .B(n622), .ZN(n625) );
  INV_X1 U693 ( .A(G952), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n624), .A2(G953), .ZN(n658) );
  NAND2_X1 U695 ( .A1(n625), .A2(n658), .ZN(n627) );
  XNOR2_X1 U696 ( .A(n627), .B(n626), .ZN(G60) );
  XOR2_X1 U697 ( .A(G110), .B(n628), .Z(G12) );
  XNOR2_X1 U698 ( .A(n629), .B(G101), .ZN(G3) );
  XOR2_X1 U699 ( .A(n631), .B(G119), .Z(G21) );
  INV_X1 U700 ( .A(KEYINPUT124), .ZN(n636) );
  NAND2_X1 U701 ( .A1(n652), .A2(G217), .ZN(n633) );
  XNOR2_X1 U702 ( .A(n633), .B(n632), .ZN(n634) );
  NAND2_X1 U703 ( .A1(n634), .A2(n658), .ZN(n635) );
  XNOR2_X1 U704 ( .A(n636), .B(n635), .ZN(G66) );
  NAND2_X1 U705 ( .A1(n652), .A2(G472), .ZN(n639) );
  XNOR2_X1 U706 ( .A(n637), .B(KEYINPUT62), .ZN(n638) );
  XNOR2_X1 U707 ( .A(n639), .B(n638), .ZN(n640) );
  NAND2_X1 U708 ( .A1(n640), .A2(n658), .ZN(n641) );
  XNOR2_X1 U709 ( .A(n641), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U710 ( .A1(n652), .A2(G478), .ZN(n642) );
  XOR2_X1 U711 ( .A(n643), .B(n642), .Z(n644) );
  INV_X1 U712 ( .A(n658), .ZN(n650) );
  NOR2_X1 U713 ( .A1(n644), .A2(n650), .ZN(G63) );
  NAND2_X1 U714 ( .A1(n652), .A2(G469), .ZN(n649) );
  XOR2_X1 U715 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n645) );
  XNOR2_X1 U716 ( .A(n645), .B(KEYINPUT58), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n649), .B(n648), .ZN(n651) );
  NOR2_X1 U719 ( .A1(n651), .A2(n650), .ZN(G54) );
  NAND2_X1 U720 ( .A1(n652), .A2(G210), .ZN(n657) );
  XNOR2_X1 U721 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n654) );
  XOR2_X1 U722 ( .A(n654), .B(KEYINPUT55), .Z(n655) );
  XNOR2_X1 U723 ( .A(n653), .B(n655), .ZN(n656) );
  XNOR2_X1 U724 ( .A(n657), .B(n656), .ZN(n659) );
  NAND2_X1 U725 ( .A1(n659), .A2(n658), .ZN(n661) );
  XOR2_X1 U726 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n660) );
  XNOR2_X1 U727 ( .A(n661), .B(n660), .ZN(G51) );
  XOR2_X1 U728 ( .A(n662), .B(KEYINPUT78), .Z(n664) );
  NAND2_X1 U729 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U730 ( .A(n665), .B(KEYINPUT80), .ZN(n706) );
  INV_X1 U731 ( .A(KEYINPUT50), .ZN(n667) );
  XNOR2_X1 U732 ( .A(n668), .B(n667), .ZN(n670) );
  NAND2_X1 U733 ( .A1(n670), .A2(n669), .ZN(n675) );
  NAND2_X1 U734 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U735 ( .A(KEYINPUT49), .B(n673), .ZN(n674) );
  NOR2_X1 U736 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U737 ( .A(n676), .B(KEYINPUT116), .ZN(n678) );
  NOR2_X1 U738 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U739 ( .A(KEYINPUT51), .B(n679), .Z(n680) );
  NOR2_X1 U740 ( .A1(n699), .A2(n680), .ZN(n693) );
  INV_X1 U741 ( .A(n681), .ZN(n685) );
  NOR2_X1 U742 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U743 ( .A1(n685), .A2(n684), .ZN(n689) );
  NOR2_X1 U744 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U745 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U746 ( .A1(n700), .A2(n690), .ZN(n691) );
  XOR2_X1 U747 ( .A(KEYINPUT117), .B(n691), .Z(n692) );
  NOR2_X1 U748 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U749 ( .A(KEYINPUT52), .B(n694), .Z(n695) );
  XNOR2_X1 U750 ( .A(KEYINPUT118), .B(n695), .ZN(n696) );
  AND2_X1 U751 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U752 ( .A1(G952), .A2(n698), .ZN(n702) );
  OR2_X1 U753 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U754 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U755 ( .A(KEYINPUT119), .B(n703), .ZN(n704) );
  AND2_X1 U756 ( .A1(n704), .A2(n406), .ZN(n705) );
  NAND2_X1 U757 ( .A1(n706), .A2(n705), .ZN(n708) );
  XOR2_X1 U758 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n707) );
  XNOR2_X1 U759 ( .A(n708), .B(n707), .ZN(G75) );
  NAND2_X1 U760 ( .A1(n710), .A2(n720), .ZN(n709) );
  XNOR2_X1 U761 ( .A(n709), .B(G104), .ZN(G6) );
  XOR2_X1 U762 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n712) );
  NAND2_X1 U763 ( .A1(n710), .A2(n723), .ZN(n711) );
  XNOR2_X1 U764 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U765 ( .A(G107), .B(n713), .ZN(G9) );
  XOR2_X1 U766 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n715) );
  NAND2_X1 U767 ( .A1(n718), .A2(n723), .ZN(n714) );
  XNOR2_X1 U768 ( .A(n715), .B(n714), .ZN(n716) );
  XOR2_X1 U769 ( .A(G128), .B(n716), .Z(G30) );
  XOR2_X1 U770 ( .A(G143), .B(n717), .Z(G45) );
  NAND2_X1 U771 ( .A1(n718), .A2(n720), .ZN(n719) );
  XNOR2_X1 U772 ( .A(n719), .B(G146), .ZN(G48) );
  NAND2_X1 U773 ( .A1(n724), .A2(n720), .ZN(n721) );
  XNOR2_X1 U774 ( .A(n721), .B(KEYINPUT114), .ZN(n722) );
  XNOR2_X1 U775 ( .A(G113), .B(n722), .ZN(G15) );
  NAND2_X1 U776 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U777 ( .A(n725), .B(G116), .ZN(G18) );
  XNOR2_X1 U778 ( .A(G125), .B(n726), .ZN(n727) );
  XNOR2_X1 U779 ( .A(n727), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U780 ( .A(G134), .B(n728), .ZN(G36) );
  XOR2_X1 U781 ( .A(G140), .B(n729), .Z(n730) );
  XNOR2_X1 U782 ( .A(n730), .B(KEYINPUT115), .ZN(G42) );
  XNOR2_X1 U783 ( .A(n731), .B(G101), .ZN(n733) );
  NOR2_X1 U784 ( .A1(n733), .A2(n732), .ZN(n742) );
  NAND2_X1 U785 ( .A1(G953), .A2(G224), .ZN(n734) );
  XOR2_X1 U786 ( .A(KEYINPUT61), .B(n734), .Z(n735) );
  NOR2_X1 U787 ( .A1(n736), .A2(n735), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n737), .A2(n406), .ZN(n738) );
  XNOR2_X1 U789 ( .A(n738), .B(KEYINPUT125), .ZN(n739) );
  NOR2_X1 U790 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U791 ( .A(n742), .B(n741), .Z(n743) );
  XNOR2_X1 U792 ( .A(KEYINPUT126), .B(n743), .ZN(G69) );
  XNOR2_X1 U793 ( .A(n744), .B(KEYINPUT127), .ZN(n746) );
  XNOR2_X1 U794 ( .A(n746), .B(n745), .ZN(n749) );
  XNOR2_X1 U795 ( .A(n749), .B(n747), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n748), .A2(n406), .ZN(n753) );
  XNOR2_X1 U797 ( .A(G227), .B(n749), .ZN(n750) );
  NAND2_X1 U798 ( .A1(n750), .A2(G900), .ZN(n751) );
  NAND2_X1 U799 ( .A1(G953), .A2(n751), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n753), .A2(n752), .ZN(G72) );
  XOR2_X1 U801 ( .A(G137), .B(n754), .Z(G39) );
  XOR2_X1 U802 ( .A(G131), .B(n755), .Z(G33) );
endmodule

