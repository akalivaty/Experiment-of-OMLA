//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G8gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G43gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(KEYINPUT86), .A3(G50gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT15), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT86), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n214), .B1(new_n208), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT14), .ZN(new_n217));
  INV_X1    g016(.A(G36gat), .ZN(new_n218));
  NOR3_X1   g017(.A1(new_n217), .A2(new_n218), .A3(G29gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT14), .B(G29gat), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n219), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n210), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(new_n210), .B2(new_n221), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(new_n223), .B(KEYINPUT17), .Z(new_n225));
  AOI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(new_n207), .ZN(new_n226));
  NAND2_X1  g025(.A1(G229gat), .A2(G233gat), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n228), .A2(KEYINPUT18), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(KEYINPUT18), .A3(new_n227), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n206), .B(new_n223), .Z(new_n231));
  XOR2_X1   g030(.A(new_n227), .B(KEYINPUT13), .Z(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n229), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G113gat), .B(G141gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(G197gat), .ZN(new_n236));
  XOR2_X1   g035(.A(KEYINPUT11), .B(G169gat), .Z(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n238), .B(KEYINPUT12), .Z(new_n239));
  NAND2_X1  g038(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n239), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n229), .A2(new_n241), .A3(new_n230), .A4(new_n233), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT30), .ZN(new_n245));
  XNOR2_X1  g044(.A(G8gat), .B(G36gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(G64gat), .B(G92gat), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g047(.A(new_n248), .B(KEYINPUT70), .Z(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n251));
  INV_X1    g050(.A(G226gat), .ZN(new_n252));
  INV_X1    g051(.A(G233gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(KEYINPUT29), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT27), .B(G183gat), .ZN(new_n258));
  INV_X1    g057(.A(G190gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT28), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT66), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT66), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT28), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n258), .A2(new_n259), .A3(new_n261), .A4(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G183gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT27), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT27), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G183gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n268), .A3(new_n259), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n261), .A2(new_n263), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT26), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n264), .A2(new_n271), .A3(new_n272), .A4(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n272), .A2(KEYINPUT24), .ZN(new_n279));
  OR2_X1    g078(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n280));
  NAND2_X1  g079(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n273), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT24), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n265), .A2(G190gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n259), .A2(G183gat), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT25), .B1(new_n284), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT25), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293));
  OAI221_X1 g092(.A(new_n291), .B1(KEYINPUT65), .B2(new_n292), .C1(new_n283), .C2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n278), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n273), .B1(new_n280), .B2(new_n281), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n296), .A2(new_n288), .A3(new_n279), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n291), .B1(new_n283), .B2(new_n293), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT65), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n292), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n257), .B1(new_n295), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n300), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n284), .A2(new_n289), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT25), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n294), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(new_n297), .B2(KEYINPUT25), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT68), .A4(new_n278), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n256), .B1(new_n302), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n305), .A2(new_n307), .A3(new_n278), .ZN(new_n310));
  INV_X1    g109(.A(new_n254), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  OR2_X1    g112(.A1(G197gat), .A2(G204gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(G197gat), .A2(G204gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT22), .ZN(new_n316));
  NAND2_X1  g115(.A1(G211gat), .A2(G218gat), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n314), .A2(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G211gat), .ZN(new_n319));
  INV_X1    g118(.A(G218gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(KEYINPUT67), .A3(new_n317), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n318), .B(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n251), .B1(new_n313), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  OAI211_X1 g125(.A(KEYINPUT69), .B(new_n323), .C1(new_n309), .C2(new_n312), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n255), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n302), .A2(new_n308), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n324), .B(new_n328), .C1(new_n329), .C2(new_n311), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n250), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n327), .A2(new_n330), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n333), .A2(new_n248), .A3(new_n325), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n245), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G134gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G127gat), .ZN(new_n337));
  INV_X1    g136(.A(G127gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G134gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G113gat), .B(G120gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(KEYINPUT1), .ZN(new_n342));
  INV_X1    g141(.A(G120gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G113gat), .ZN(new_n344));
  INV_X1    g143(.A(G113gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G120gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G127gat), .B(G134gat), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT1), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n342), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(new_n295), .B2(new_n301), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n342), .A2(new_n350), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n305), .A2(new_n307), .A3(new_n353), .A4(new_n278), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT34), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT34), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n352), .A2(new_n354), .A3(new_n359), .A4(new_n356), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(G15gat), .B(G43gat), .Z(new_n362));
  XNOR2_X1  g161(.A(G71gat), .B(G99gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n355), .A2(new_n357), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT33), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n361), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n361), .A2(new_n368), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n369), .A2(KEYINPUT32), .A3(new_n366), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n366), .A2(KEYINPUT32), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n361), .A2(new_n368), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n361), .A2(new_n368), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n334), .A2(new_n245), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n335), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT35), .ZN(new_n379));
  NAND2_X1  g178(.A1(G228gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n324), .B2(KEYINPUT29), .ZN(new_n382));
  AND2_X1   g181(.A1(G141gat), .A2(G148gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(G141gat), .A2(G148gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT2), .ZN(new_n387));
  AND2_X1   g186(.A1(G155gat), .A2(G162gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(G155gat), .A2(G162gat), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n385), .B(new_n387), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G141gat), .B(G148gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT72), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT2), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n393), .A2(new_n394), .B1(G155gat), .B2(G162gat), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n391), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT71), .B1(new_n388), .B2(new_n389), .ZN(new_n397));
  INV_X1    g196(.A(G155gat), .ZN(new_n398));
  INV_X1    g197(.A(G162gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT71), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n401), .A3(new_n386), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n390), .B1(new_n396), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n380), .B1(new_n382), .B2(new_n404), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n381), .B(new_n390), .C1(new_n396), .C2(new_n403), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n324), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n317), .ZN(new_n411));
  NOR2_X1   g210(.A1(G211gat), .A2(G218gat), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT79), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT79), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n321), .A2(new_n414), .A3(new_n317), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n318), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n407), .B1(new_n318), .B2(new_n413), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n381), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n404), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n323), .B1(new_n406), .B2(new_n407), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT80), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI211_X1 g221(.A(KEYINPUT80), .B(new_n323), .C1(new_n407), .C2(new_n406), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n380), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT81), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g225(.A(KEYINPUT81), .B(new_n380), .C1(new_n422), .C2(new_n423), .ZN(new_n427));
  AOI211_X1 g226(.A(G22gat), .B(new_n410), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G22gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n427), .ZN(new_n430));
  INV_X1    g229(.A(new_n410), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(G78gat), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n409), .A2(KEYINPUT80), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n420), .A2(new_n421), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n419), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT81), .B1(new_n436), .B2(new_n380), .ZN(new_n437));
  INV_X1    g236(.A(new_n427), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n431), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(G22gat), .ZN(new_n440));
  INV_X1    g239(.A(G78gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n430), .A2(new_n429), .A3(new_n431), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT31), .B(G50gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n444), .B(G106gat), .Z(new_n445));
  NAND3_X1  g244(.A1(new_n433), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n445), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n428), .A2(new_n432), .A3(G78gat), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n441), .B1(new_n440), .B2(new_n442), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n378), .A2(new_n379), .A3(new_n446), .A4(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT84), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n404), .A2(new_n351), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n453), .A2(KEYINPUT4), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT74), .B1(new_n404), .B2(new_n351), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT74), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n393), .A2(new_n394), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(new_n392), .A3(new_n386), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n385), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(new_n397), .A3(new_n402), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n353), .A2(new_n456), .A3(new_n460), .A4(new_n390), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n454), .B1(KEYINPUT4), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT5), .ZN(new_n464));
  NAND2_X1  g263(.A1(G225gat), .A2(G233gat), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n404), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT73), .B1(new_n404), .B2(KEYINPUT3), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n351), .B(new_n406), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n463), .A2(new_n464), .A3(new_n465), .A4(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n453), .A2(KEYINPUT4), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT4), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n461), .A3(new_n472), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n468), .A2(new_n465), .A3(new_n471), .A4(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT75), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n404), .A2(new_n351), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n455), .A2(new_n461), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n465), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n475), .B1(new_n479), .B2(KEYINPUT5), .ZN(new_n480));
  AOI211_X1 g279(.A(KEYINPUT75), .B(new_n464), .C1(new_n477), .C2(new_n478), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n474), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT76), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT76), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n484), .B(new_n474), .C1(new_n480), .C2(new_n481), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n470), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  XOR2_X1   g285(.A(G1gat), .B(G29gat), .Z(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G57gat), .B(G85gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n452), .B1(new_n493), .B2(KEYINPUT6), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT5), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT75), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n475), .A3(KEYINPUT5), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n484), .B1(new_n498), .B2(new_n474), .ZN(new_n499));
  INV_X1    g298(.A(new_n485), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n469), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(KEYINPUT6), .A3(new_n491), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(new_n486), .B2(new_n492), .ZN(new_n504));
  AOI211_X1 g303(.A(new_n491), .B(new_n470), .C1(new_n483), .C2(new_n485), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n494), .B1(new_n506), .B2(new_n452), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n451), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n335), .A2(new_n377), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n506), .A2(KEYINPUT78), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT78), .B1(new_n506), .B2(new_n509), .ZN(new_n511));
  INV_X1    g310(.A(new_n376), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n450), .A2(new_n446), .A3(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n508), .B1(new_n514), .B2(new_n379), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT37), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n333), .A2(new_n516), .A3(new_n325), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n324), .B1(new_n309), .B2(new_n312), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n328), .B1(new_n329), .B2(new_n311), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n518), .B(KEYINPUT37), .C1(new_n324), .C2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n249), .A2(KEYINPUT38), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n334), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT85), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n516), .B1(new_n333), .B2(new_n325), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n524), .B1(new_n525), .B2(new_n248), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT37), .B1(new_n326), .B2(new_n331), .ZN(new_n527));
  INV_X1    g326(.A(new_n248), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(KEYINPUT85), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n529), .A3(new_n517), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n523), .B1(new_n530), .B2(KEYINPUT38), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n506), .A2(new_n452), .ZN(new_n532));
  INV_X1    g331(.A(new_n494), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n450), .A2(new_n446), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT82), .ZN(new_n536));
  AOI211_X1 g335(.A(KEYINPUT39), .B(new_n465), .C1(new_n463), .C2(new_n468), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(new_n491), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n465), .B1(new_n463), .B2(new_n468), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT39), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n541), .A2(KEYINPUT82), .A3(new_n492), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT39), .B1(new_n477), .B2(new_n478), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n538), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT40), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n545), .A2(KEYINPUT83), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n546), .B1(new_n545), .B2(KEYINPUT83), .ZN(new_n548));
  NOR3_X1   g347(.A1(new_n547), .A2(new_n548), .A3(new_n493), .ZN(new_n549));
  INV_X1    g348(.A(new_n509), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n535), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n535), .B1(new_n510), .B2(new_n511), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT36), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n376), .B(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n244), .B1(new_n515), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G85gat), .A2(G92gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT7), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT91), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n558), .B2(KEYINPUT7), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT7), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n563), .A2(KEYINPUT92), .A3(G85gat), .A4(G92gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT91), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n558), .A2(new_n565), .A3(KEYINPUT7), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n560), .A2(new_n562), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(G85gat), .ZN(new_n569));
  INV_X1    g368(.A(G92gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(KEYINPUT8), .A2(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G99gat), .B(G106gat), .Z(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT93), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n573), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G71gat), .B(G78gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(KEYINPUT87), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(G57gat), .B(G64gat), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n578), .A2(KEYINPUT87), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n572), .A2(KEYINPUT93), .A3(new_n573), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n577), .A2(new_n584), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n585), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(new_n574), .A3(new_n576), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G230gat), .A2(G233gat), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n591), .B(KEYINPUT96), .Z(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(G120gat), .B(G148gat), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT98), .ZN(new_n595));
  XNOR2_X1  g394(.A(G176gat), .B(G204gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n592), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n577), .A2(new_n586), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n588), .A2(KEYINPUT10), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n604), .A3(new_n589), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT94), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n587), .A2(KEYINPUT94), .A3(new_n604), .A4(new_n589), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n603), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n600), .B1(new_n609), .B2(KEYINPUT95), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(KEYINPUT95), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(KEYINPUT97), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT97), .ZN(new_n614));
  INV_X1    g413(.A(new_n612), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n614), .B1(new_n615), .B2(new_n610), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n599), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n607), .A2(new_n608), .ZN(new_n618));
  INV_X1    g417(.A(new_n603), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n592), .B(KEYINPUT99), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n598), .B1(new_n623), .B2(new_n593), .ZN(new_n624));
  OR3_X1    g423(.A1(new_n617), .A2(KEYINPUT100), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(KEYINPUT100), .B1(new_n617), .B2(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n225), .A2(new_n601), .ZN(new_n628));
  NAND3_X1  g427(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n628), .B(new_n629), .C1(new_n223), .C2(new_n601), .ZN(new_n630));
  XNOR2_X1  g429(.A(G190gat), .B(G218gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G134gat), .B(G162gat), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n632), .A2(new_n635), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n206), .B1(new_n588), .B2(KEYINPUT21), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT90), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n588), .A2(KEYINPUT21), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n640), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G127gat), .B(G155gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT20), .ZN(new_n646));
  NAND2_X1  g445(.A1(G231gat), .A2(G233gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n647), .B(KEYINPUT88), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n646), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G183gat), .B(G211gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n644), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n644), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n627), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n557), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n506), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(G1gat), .ZN(G1324gat));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  NAND3_X1  g463(.A1(new_n659), .A2(new_n550), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(G8gat), .B1(new_n658), .B2(new_n509), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n667), .B1(new_n663), .B2(new_n665), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT101), .Z(G1325gat));
  OAI21_X1  g468(.A(G15gat), .B1(new_n658), .B2(new_n555), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n376), .A2(G15gat), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n670), .B1(new_n658), .B2(new_n671), .ZN(G1326gat));
  NAND2_X1  g471(.A1(new_n659), .A2(new_n535), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT102), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT43), .B(G22gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  AND3_X1   g475(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n451), .A2(new_n507), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n506), .A2(new_n509), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT78), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n506), .A2(KEYINPUT78), .A3(new_n509), .ZN(new_n682));
  INV_X1    g481(.A(new_n513), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n678), .B1(new_n684), .B2(KEYINPUT35), .ZN(new_n685));
  OAI211_X1 g484(.A(KEYINPUT105), .B(new_n638), .C1(new_n677), .C2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n515), .A2(new_n556), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n689), .A2(KEYINPUT105), .A3(KEYINPUT44), .A4(new_n638), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n240), .A2(KEYINPUT103), .A3(new_n242), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT103), .B1(new_n240), .B2(new_n242), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n654), .B(KEYINPUT104), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n627), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n688), .A2(new_n690), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n688), .A2(KEYINPUT106), .A3(new_n690), .A4(new_n696), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n660), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(G29gat), .ZN(new_n702));
  INV_X1    g501(.A(new_n654), .ZN(new_n703));
  INV_X1    g502(.A(new_n638), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n627), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n557), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n706), .A2(G29gat), .A3(new_n506), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT45), .Z(new_n708));
  NAND2_X1  g507(.A1(new_n702), .A2(new_n708), .ZN(G1328gat));
  NOR3_X1   g508(.A1(new_n706), .A2(G36gat), .A3(new_n509), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT107), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(KEYINPUT46), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n699), .A2(new_n550), .A3(new_n700), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n715));
  OAI221_X1 g514(.A(new_n713), .B1(new_n218), .B2(new_n714), .C1(new_n711), .C2(new_n715), .ZN(G1329gat));
  INV_X1    g515(.A(new_n706), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n376), .A2(G43gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n555), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n699), .A2(new_n722), .A3(new_n700), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n721), .B1(new_n723), .B2(G43gat), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n688), .A2(new_n722), .A3(new_n690), .A4(new_n696), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n211), .B1(new_n727), .B2(new_n728), .ZN(new_n730));
  AOI22_X1  g529(.A1(new_n729), .A2(new_n730), .B1(new_n717), .B2(new_n718), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n725), .B(new_n726), .C1(new_n720), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n730), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n720), .B1(new_n733), .B2(new_n719), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT110), .B1(new_n734), .B2(new_n724), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(G1330gat));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n737));
  INV_X1    g536(.A(G50gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n717), .A2(new_n738), .A3(new_n535), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n688), .A2(new_n535), .A3(new_n690), .A4(new_n696), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT111), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G50gat), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n740), .A2(KEYINPUT111), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n739), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT48), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n739), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n699), .A2(new_n535), .A3(new_n700), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(G50gat), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n737), .B1(new_n745), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n738), .B1(new_n740), .B2(KEYINPUT111), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n686), .A2(new_n687), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n704), .B1(new_n515), .B2(new_n556), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT44), .B1(new_n754), .B2(KEYINPUT105), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n756), .A2(new_n757), .A3(new_n535), .A4(new_n696), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n752), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n746), .B1(new_n759), .B2(new_n739), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n760), .A2(KEYINPUT112), .A3(new_n749), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n751), .A2(new_n761), .ZN(G1331gat));
  NAND3_X1  g561(.A1(new_n627), .A2(new_n655), .A3(new_n693), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT113), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n764), .A2(new_n689), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n660), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n550), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n769));
  XOR2_X1   g568(.A(KEYINPUT49), .B(G64gat), .Z(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n768), .B2(new_n770), .ZN(G1333gat));
  NAND2_X1  g570(.A1(new_n765), .A2(new_n722), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n376), .A2(G71gat), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n772), .A2(G71gat), .B1(new_n765), .B2(new_n773), .ZN(new_n774));
  XOR2_X1   g573(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1334gat));
  NAND2_X1  g575(.A1(new_n765), .A2(new_n535), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n754), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n693), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n703), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n754), .A2(new_n779), .ZN(new_n785));
  OR3_X1    g584(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n783), .B2(new_n785), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n627), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n660), .A2(new_n569), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n782), .A2(new_n627), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT115), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n756), .A2(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n793), .A2(new_n660), .ZN(new_n794));
  OAI22_X1  g593(.A1(new_n789), .A2(new_n790), .B1(new_n794), .B2(new_n569), .ZN(G1336gat));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n509), .A2(G92gat), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n756), .A2(new_n550), .A3(new_n792), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G92gat), .ZN(new_n803));
  OAI221_X1 g602(.A(new_n796), .B1(new_n789), .B2(new_n798), .C1(new_n801), .C2(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n798), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n799), .A2(G92gat), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT52), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(G1337gat));
  NAND3_X1  g607(.A1(new_n788), .A2(new_n512), .A3(new_n627), .ZN(new_n809));
  INV_X1    g608(.A(G99gat), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n555), .A2(new_n810), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n809), .A2(new_n810), .B1(new_n793), .B2(new_n811), .ZN(G1338gat));
  NAND2_X1  g611(.A1(new_n793), .A2(new_n535), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G106gat), .ZN(new_n814));
  INV_X1    g613(.A(new_n535), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(G106gat), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n788), .A2(new_n627), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n818), .B(new_n819), .ZN(G1339gat));
  OAI21_X1  g619(.A(new_n597), .B1(new_n623), .B2(KEYINPUT54), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n613), .A2(new_n616), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n609), .A2(KEYINPUT120), .A3(new_n621), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT120), .B1(new_n609), .B2(new_n621), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n821), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n617), .B1(new_n827), .B2(KEYINPUT55), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n822), .A2(new_n826), .ZN(new_n829));
  INV_X1    g628(.A(new_n821), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT121), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n827), .A2(new_n834), .A3(KEYINPUT55), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n781), .B(new_n828), .C1(new_n833), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n226), .A2(new_n227), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n231), .A2(new_n232), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n238), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n242), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n625), .B2(new_n626), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n638), .B1(new_n836), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n831), .A2(KEYINPUT121), .A3(new_n832), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n834), .B1(new_n827), .B2(KEYINPUT55), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n704), .A2(new_n840), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n828), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n694), .B1(new_n843), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n693), .A2(new_n625), .A3(new_n655), .A4(new_n626), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT119), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n535), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n854), .A2(new_n660), .A3(new_n378), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n345), .A3(new_n781), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n243), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(G113gat), .ZN(new_n859));
  AOI211_X1 g658(.A(KEYINPUT122), .B(new_n345), .C1(new_n855), .C2(new_n243), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(G1340gat));
  INV_X1    g660(.A(new_n855), .ZN(new_n862));
  INV_X1    g661(.A(new_n627), .ZN(new_n863));
  OAI21_X1  g662(.A(G120gat), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n627), .A2(new_n343), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT123), .Z(new_n866));
  OAI21_X1  g665(.A(new_n864), .B1(new_n862), .B2(new_n866), .ZN(G1341gat));
  OAI21_X1  g666(.A(new_n338), .B1(new_n862), .B2(new_n654), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n695), .A2(G127gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n862), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n855), .A2(KEYINPUT124), .A3(G127gat), .A4(new_n695), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n868), .A2(new_n871), .A3(new_n872), .ZN(G1342gat));
  OAI21_X1  g672(.A(G134gat), .B1(new_n862), .B2(new_n704), .ZN(new_n874));
  INV_X1    g673(.A(new_n854), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(new_n506), .ZN(new_n876));
  NOR4_X1   g675(.A1(new_n704), .A2(G134gat), .A3(new_n550), .A4(new_n376), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n876), .A2(KEYINPUT56), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT56), .B1(new_n876), .B2(new_n877), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n874), .B1(new_n878), .B2(new_n879), .ZN(G1343gat));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n815), .B1(new_n850), .B2(new_n853), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n722), .A2(new_n506), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n509), .ZN(new_n886));
  INV_X1    g685(.A(new_n617), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(new_n831), .B2(new_n832), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n243), .B1(new_n827), .B2(KEYINPUT55), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n704), .B1(new_n890), .B2(new_n841), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n703), .B1(new_n891), .B2(new_n848), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n535), .B1(new_n892), .B2(new_n852), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n886), .B1(new_n893), .B2(KEYINPUT57), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n884), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n881), .B(G141gat), .C1(new_n895), .C2(new_n244), .ZN(new_n896));
  NAND2_X1  g695(.A1(KEYINPUT125), .A2(KEYINPUT58), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n882), .A2(new_n885), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n509), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n244), .A2(G141gat), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n896), .B(new_n897), .C1(new_n899), .C2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n899), .A2(new_n901), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n884), .A2(new_n894), .A3(new_n781), .ZN(new_n904));
  AOI22_X1  g703(.A1(new_n903), .A2(KEYINPUT125), .B1(G141gat), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n902), .B1(new_n905), .B2(new_n881), .ZN(G1344gat));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n627), .A2(new_n243), .A3(new_n656), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n883), .B(new_n535), .C1(new_n892), .C2(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n863), .A2(new_n886), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n909), .B(new_n910), .C1(new_n882), .C2(new_n883), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G148gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n884), .A2(new_n894), .A3(new_n627), .ZN(new_n913));
  INV_X1    g712(.A(G148gat), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(KEYINPUT59), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n912), .A2(KEYINPUT59), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n898), .A2(new_n914), .A3(new_n509), .A4(new_n627), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n907), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n913), .A2(new_n915), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n921), .B1(new_n911), .B2(G148gat), .ZN(new_n922));
  OAI211_X1 g721(.A(KEYINPUT126), .B(new_n917), .C1(new_n920), .C2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n919), .A2(new_n923), .ZN(G1345gat));
  OAI21_X1  g723(.A(G155gat), .B1(new_n895), .B2(new_n694), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n703), .A2(new_n398), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n899), .B2(new_n926), .ZN(G1346gat));
  OAI21_X1  g726(.A(G162gat), .B1(new_n895), .B2(new_n704), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n898), .A2(new_n399), .A3(new_n509), .A4(new_n638), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1347gat));
  NAND2_X1  g729(.A1(new_n550), .A2(new_n506), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n931), .A2(new_n376), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n854), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(G169gat), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n933), .A2(new_n934), .A3(new_n244), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n660), .B1(new_n850), .B2(new_n853), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(new_n550), .A3(new_n683), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n781), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n935), .B1(new_n938), .B2(new_n934), .ZN(G1348gat));
  INV_X1    g738(.A(G176gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n937), .A2(new_n940), .A3(new_n627), .ZN(new_n941));
  OAI21_X1  g740(.A(G176gat), .B1(new_n933), .B2(new_n863), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1349gat));
  NAND3_X1  g742(.A1(new_n937), .A2(new_n258), .A3(new_n703), .ZN(new_n944));
  OAI21_X1  g743(.A(G183gat), .B1(new_n933), .B2(new_n694), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g746(.A1(new_n937), .A2(new_n259), .A3(new_n638), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n949));
  INV_X1    g748(.A(new_n933), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n638), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n949), .B1(new_n951), .B2(G190gat), .ZN(new_n952));
  AOI211_X1 g751(.A(KEYINPUT61), .B(new_n259), .C1(new_n950), .C2(new_n638), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n948), .B1(new_n952), .B2(new_n953), .ZN(G1351gat));
  OR2_X1    g753(.A1(new_n882), .A2(new_n883), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n722), .A2(new_n931), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(new_n909), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n243), .A2(G197gat), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n722), .A2(new_n815), .A3(new_n509), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n936), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n960), .A2(new_n693), .ZN(new_n961));
  OAI22_X1  g760(.A1(new_n957), .A2(new_n958), .B1(new_n961), .B2(G197gat), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(G1352gat));
  OAI21_X1  g762(.A(G204gat), .B1(new_n957), .B2(new_n863), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n960), .A2(G204gat), .A3(new_n863), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n964), .A2(new_n967), .A3(new_n968), .ZN(G1353gat));
  INV_X1    g768(.A(new_n960), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n970), .A2(new_n319), .A3(new_n703), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n955), .A2(new_n703), .A3(new_n909), .A4(new_n956), .ZN(new_n972));
  AND2_X1   g771(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n973));
  OAI21_X1  g772(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n973), .B1(new_n972), .B2(new_n975), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n971), .B1(new_n977), .B2(new_n978), .ZN(G1354gat));
  OAI21_X1  g778(.A(G218gat), .B1(new_n957), .B2(new_n704), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n970), .A2(new_n320), .A3(new_n638), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1355gat));
endmodule


