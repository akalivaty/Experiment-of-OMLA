//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n621, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1205, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(KEYINPUT68), .B(G125), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n461), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n474), .B1(new_n464), .B2(new_n465), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT69), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n474), .B(new_n477), .C1(new_n465), .C2(new_n464), .ZN(new_n478));
  AOI211_X1 g053(.A(new_n463), .B(new_n472), .C1(new_n476), .C2(new_n478), .ZN(G160));
  OR2_X1    g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n461), .B1(new_n480), .B2(new_n481), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n491), .A2(new_n493), .A3(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n464), .B2(new_n465), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT3), .B(G2104), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(new_n497), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n495), .B1(new_n499), .B2(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n504), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT70), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n507), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(G543), .B1(new_n508), .B2(new_n509), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n519), .A2(G651), .B1(new_n521), .B2(G50), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n516), .A2(new_n522), .ZN(G166));
  NAND2_X1  g098(.A1(new_n515), .A2(G89), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n520), .A2(KEYINPUT71), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n526), .B(G543), .C1(new_n508), .C2(new_n509), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n531), .A2(new_n532), .B1(new_n512), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n524), .A2(new_n529), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND2_X1  g111(.A1(new_n515), .A2(G90), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT72), .B(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n528), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G651), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n537), .A2(new_n539), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND2_X1  g119(.A1(new_n528), .A2(G43), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n511), .A2(G81), .A3(new_n514), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n547));
  OAI21_X1  g122(.A(G56), .B1(new_n505), .B2(new_n506), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n547), .B1(new_n550), .B2(G651), .ZN(new_n551));
  AOI211_X1 g126(.A(KEYINPUT73), .B(new_n541), .C1(new_n548), .C2(new_n549), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n545), .B(new_n546), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND3_X1  g134(.A1(new_n511), .A2(G91), .A3(new_n514), .ZN(new_n560));
  NAND2_X1  g135(.A1(KEYINPUT74), .A2(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT9), .B1(new_n520), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(new_n561), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n513), .A2(new_n563), .A3(G543), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n507), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n560), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n560), .A2(new_n566), .A3(KEYINPUT75), .A4(new_n570), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G299));
  NAND2_X1  g151(.A1(new_n516), .A2(new_n522), .ZN(G303));
  NAND2_X1  g152(.A1(new_n515), .A2(G87), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n512), .A2(G74), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(new_n521), .B2(G49), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(G288));
  AND2_X1   g156(.A1(new_n512), .A2(G61), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  OAI211_X1 g159(.A(KEYINPUT76), .B(G651), .C1(new_n582), .C2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT76), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n584), .B1(new_n512), .B2(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n587), .B2(new_n541), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n521), .A2(G48), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n585), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n511), .A2(KEYINPUT77), .A3(G86), .A4(new_n514), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n511), .A2(G86), .A3(new_n514), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n590), .A2(new_n591), .A3(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(new_n515), .A2(G85), .ZN(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT78), .B(G47), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n528), .A2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n541), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n511), .A2(new_n514), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n511), .A2(KEYINPUT10), .A3(G92), .A4(new_n514), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT79), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n541), .B1(new_n609), .B2(new_n610), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n611), .A2(new_n612), .B1(G54), .B2(new_n528), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n602), .B1(new_n615), .B2(G868), .ZN(G284));
  OAI21_X1  g191(.A(new_n602), .B1(new_n615), .B2(G868), .ZN(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n575), .B2(G868), .ZN(G297));
  OAI21_X1  g194(.A(new_n618), .B1(new_n575), .B2(G868), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n615), .B1(new_n621), .B2(G860), .ZN(G148));
  OAI21_X1  g197(.A(KEYINPUT80), .B1(new_n554), .B2(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n615), .A2(new_n621), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  MUX2_X1   g200(.A(KEYINPUT80), .B(new_n623), .S(new_n625), .Z(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n500), .A2(new_n462), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g205(.A(G2100), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  AOI22_X1  g208(.A1(G123), .A2(new_n484), .B1(new_n482), .B2(G135), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  INV_X1    g210(.A(G111), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n635), .A2(KEYINPUT81), .B1(new_n636), .B2(G2105), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(KEYINPUT81), .B2(new_n635), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(G2096), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n632), .A2(new_n633), .A3(new_n641), .ZN(G156));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(G14), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(G401));
  XNOR2_X1  g233(.A(G2072), .B(G2078), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT17), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT82), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n660), .A2(new_n661), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n666), .B(new_n663), .C1(new_n659), .C2(new_n661), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n662), .A2(new_n659), .A3(new_n661), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  NAND3_X1  g244(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n640), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT83), .B(G2100), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1961), .B(G1966), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n677), .A2(new_n678), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n676), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n676), .B2(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(G229));
  NAND2_X1  g266(.A1(new_n482), .A2(G140), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n484), .A2(G128), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n461), .A2(G116), .ZN(new_n694));
  OAI21_X1  g269(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n692), .B(new_n693), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G29), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G26), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT89), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT88), .B(G2067), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT85), .B(G16), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(G19), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n554), .B2(new_n706), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(G1341), .Z(new_n709));
  NOR2_X1   g284(.A1(G4), .A2(G16), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT87), .Z(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n614), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1348), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n704), .A2(new_n709), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n712), .A2(G21), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G168), .B2(new_n712), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G1966), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT92), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n712), .A2(G5), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G171), .B2(new_n712), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(G1961), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n482), .A2(G141), .B1(G105), .B2(new_n462), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n484), .A2(G129), .ZN(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT26), .Z(new_n728));
  NAND3_X1  g303(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT91), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G29), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G29), .B2(G32), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT27), .B(G1996), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AND2_X1   g309(.A1(KEYINPUT24), .A2(G34), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n698), .B1(KEYINPUT24), .B2(G34), .ZN(new_n736));
  OAI22_X1  g311(.A1(G160), .A2(new_n698), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G2084), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n723), .A2(G1961), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n724), .A2(new_n734), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n721), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n715), .A2(new_n716), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n698), .A2(G33), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT25), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n500), .A2(G127), .ZN(new_n746));
  NAND2_X1  g321(.A1(G115), .A2(G2104), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n461), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n745), .B(new_n748), .C1(G139), .C2(new_n482), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n743), .B1(new_n749), .B2(new_n698), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G2072), .Z(new_n751));
  XOR2_X1   g326(.A(KEYINPUT31), .B(G11), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT93), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT30), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n754), .A2(G28), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n698), .B1(new_n754), .B2(G28), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n753), .B1(new_n755), .B2(new_n756), .C1(new_n639), .C2(new_n698), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT94), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n698), .A2(G27), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G164), .B2(new_n698), .ZN(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n751), .A2(new_n758), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n698), .A2(G35), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G162), .B2(new_n698), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT29), .ZN(new_n766));
  OAI22_X1  g341(.A1(G1966), .A2(new_n719), .B1(new_n766), .B2(G2090), .ZN(new_n767));
  OAI22_X1  g342(.A1(new_n733), .A2(new_n732), .B1(new_n737), .B2(G2084), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n763), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n717), .A2(new_n741), .A3(new_n742), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n705), .A2(G20), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT95), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT23), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n575), .B2(new_n712), .ZN(new_n774));
  INV_X1    g349(.A(G1956), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n766), .A2(G2090), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT96), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n770), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n712), .A2(G23), .ZN(new_n781));
  INV_X1    g356(.A(G288), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n712), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT33), .B(G1976), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n706), .A2(G22), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G166), .B2(new_n706), .ZN(new_n787));
  INV_X1    g362(.A(G1971), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(G6), .A2(G16), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G305), .B2(new_n712), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT32), .B(G1981), .Z(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n785), .A2(new_n789), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(KEYINPUT34), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(KEYINPUT34), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n706), .A2(G24), .ZN(new_n798));
  AND3_X1   g373(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n706), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1986), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n698), .A2(G25), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n482), .A2(G131), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n484), .A2(G119), .ZN(new_n804));
  OR2_X1    g379(.A1(G95), .A2(G2105), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n805), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n802), .B1(new_n808), .B2(new_n698), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT35), .B(G1991), .Z(new_n810));
  XOR2_X1   g385(.A(new_n809), .B(new_n810), .Z(new_n811));
  NOR2_X1   g386(.A1(new_n801), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n796), .A2(new_n797), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(KEYINPUT86), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n813), .A2(new_n815), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n780), .B1(new_n816), .B2(new_n817), .ZN(G150));
  INV_X1    g393(.A(KEYINPUT97), .ZN(new_n819));
  XNOR2_X1  g394(.A(G150), .B(new_n819), .ZN(G311));
  NOR2_X1   g395(.A1(new_n614), .A2(new_n621), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT38), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n545), .A2(new_n546), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n551), .A2(new_n552), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n515), .A2(G93), .ZN(new_n825));
  NAND2_X1  g400(.A1(G80), .A2(G543), .ZN(new_n826));
  INV_X1    g401(.A(G67), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n507), .B2(new_n827), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n528), .A2(G55), .B1(new_n828), .B2(G651), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n823), .A2(new_n824), .A3(new_n825), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n526), .B1(new_n513), .B2(G543), .ZN(new_n831));
  INV_X1    g406(.A(new_n527), .ZN(new_n832));
  OAI21_X1  g407(.A(G55), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n828), .A2(G651), .ZN(new_n834));
  INV_X1    g409(.A(G93), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n833), .B(new_n834), .C1(new_n604), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n553), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n830), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n822), .B(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT98), .B(G860), .Z(new_n842));
  NAND3_X1  g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n836), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(new_n842), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n846), .ZN(G145));
  NAND2_X1  g422(.A1(new_n499), .A2(new_n502), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n490), .A2(new_n494), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n696), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n807), .ZN(new_n852));
  AOI22_X1  g427(.A1(G130), .A2(new_n484), .B1(new_n482), .B2(G142), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n854), .A2(KEYINPUT100), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT99), .ZN(new_n856));
  OR3_X1    g431(.A1(new_n856), .A2(new_n461), .A3(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n461), .B2(G118), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n857), .B(new_n858), .C1(KEYINPUT100), .C2(new_n854), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n853), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n629), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n852), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n730), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n749), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n749), .B2(new_n729), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n862), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(G160), .B(new_n639), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(G162), .ZN(new_n869));
  AOI21_X1  g444(.A(G37), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NOR3_X1   g445(.A1(new_n867), .A2(KEYINPUT101), .A3(new_n869), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n872));
  INV_X1    g447(.A(new_n869), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n872), .B1(new_n866), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n870), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g451(.A(G868), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n575), .A2(new_n614), .A3(KEYINPUT102), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT102), .B1(new_n575), .B2(new_n614), .ZN(new_n879));
  OAI21_X1  g454(.A(KEYINPUT103), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n575), .A2(new_n614), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n575), .A2(new_n614), .A3(KEYINPUT102), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(G299), .A2(new_n615), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n880), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n878), .A2(new_n879), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(G299), .B2(new_n615), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n624), .B(new_n838), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n887), .A3(new_n891), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G166), .B(G288), .ZN(new_n899));
  NAND2_X1  g474(.A1(G305), .A2(new_n799), .ZN(new_n900));
  NAND4_X1  g475(.A1(G290), .A2(new_n590), .A3(new_n591), .A4(new_n594), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(G288), .B(G303), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n901), .A3(new_n900), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n906), .A2(KEYINPUT42), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n903), .A2(new_n905), .A3(KEYINPUT104), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT104), .B1(new_n903), .B2(new_n905), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n907), .B1(new_n911), .B2(KEYINPUT42), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n877), .B1(new_n898), .B2(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n911), .A2(KEYINPUT42), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n897), .B(new_n896), .C1(new_n914), .C2(new_n907), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n913), .A2(KEYINPUT105), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(new_n844), .B2(G868), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(new_n913), .B2(new_n915), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n916), .A2(new_n919), .ZN(G295));
  NOR2_X1   g495(.A1(new_n916), .A2(new_n919), .ZN(G331));
  NAND3_X1  g496(.A1(new_n883), .A2(new_n887), .A3(new_n885), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n553), .A2(new_n836), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n553), .A2(new_n836), .ZN(new_n924));
  OAI21_X1  g499(.A(G168), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n830), .A2(G286), .A3(new_n837), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n925), .A2(G171), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(G171), .B1(new_n925), .B2(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n922), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n922), .A2(new_n889), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n925), .A2(new_n926), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(G301), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n925), .A2(G171), .A3(new_n926), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n892), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n880), .A2(new_n886), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n929), .B(new_n930), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(G37), .B1(new_n936), .B2(new_n910), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n938), .B(new_n922), .C1(new_n927), .C2(new_n928), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n929), .A2(KEYINPUT106), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n888), .A2(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n932), .A2(new_n933), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n939), .B(new_n940), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n937), .B1(new_n943), .B2(new_n910), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n942), .B1(new_n890), .B2(new_n893), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n940), .A2(new_n939), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(G37), .B1(new_n950), .B2(new_n911), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n943), .A2(new_n910), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n944), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n947), .A2(KEYINPUT44), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n952), .B1(new_n951), .B2(new_n953), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n937), .B(new_n952), .C1(new_n943), .C2(new_n910), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n957), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n956), .A2(new_n961), .ZN(G397));
  AOI21_X1  g537(.A(KEYINPUT68), .B1(new_n500), .B2(G125), .ZN(new_n963));
  INV_X1    g538(.A(new_n469), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n471), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(G2105), .ZN(new_n966));
  INV_X1    g541(.A(G40), .ZN(new_n967));
  AOI211_X1 g542(.A(new_n967), .B(new_n463), .C1(new_n476), .C2(new_n478), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(new_n968), .A3(KEYINPUT109), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n462), .A2(G101), .ZN(new_n971));
  INV_X1    g546(.A(new_n478), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n477), .B1(new_n500), .B2(new_n474), .ZN(new_n973));
  OAI211_X1 g548(.A(G40), .B(new_n971), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n970), .B1(new_n472), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n969), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(G164), .B2(G1384), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1996), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n730), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G2067), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n696), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n729), .A2(G1996), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n808), .A2(new_n810), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n808), .A2(new_n810), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(G290), .B(G1986), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n981), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n571), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n995), .B(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n978), .B1(new_n850), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  AOI211_X1 g575(.A(new_n1000), .B(G1384), .C1(new_n848), .C2(new_n849), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT56), .B(G2072), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n976), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(G164), .B2(G1384), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n850), .A2(KEYINPUT50), .A3(new_n998), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1956), .B1(new_n976), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n997), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n850), .A2(new_n998), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n969), .B2(new_n975), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n984), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n969), .A2(new_n975), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(G1348), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n615), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT117), .B(new_n997), .C1(new_n1004), .C2(new_n1009), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1012), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n996), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n995), .B(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n976), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1023), .B(new_n1024), .C1(G1956), .C2(new_n1017), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1010), .A2(new_n1025), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT61), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT118), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n1030));
  AOI211_X1 g605(.A(new_n1030), .B(KEYINPUT61), .C1(new_n1010), .C2(new_n1025), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n850), .A2(KEYINPUT45), .A3(new_n998), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n980), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n969), .B2(new_n975), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT109), .B1(new_n966), .B2(new_n968), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n472), .A2(new_n974), .A3(new_n970), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1008), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1035), .A2(new_n1003), .B1(new_n1038), .B2(new_n775), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1028), .B1(new_n1039), .B2(new_n1023), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(new_n1012), .A3(new_n1020), .ZN(new_n1041));
  INV_X1    g616(.A(G1348), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(KEYINPUT60), .A3(new_n1015), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(KEYINPUT119), .A3(new_n614), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n614), .B(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1047), .A2(KEYINPUT60), .A3(new_n1015), .A4(new_n1043), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT60), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1045), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n976), .A2(new_n982), .A3(new_n1002), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT58), .B(G1341), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1014), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n554), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT59), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1057), .B(new_n554), .C1(new_n1052), .C2(new_n1054), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1041), .A2(new_n1051), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1026), .B1(new_n1032), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT120), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1063), .B(new_n1026), .C1(new_n1032), .C2(new_n1060), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n782), .A2(G1976), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT110), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1013), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n976), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1066), .B1(new_n1068), .B2(G8), .ZN(new_n1069));
  INV_X1    g644(.A(G8), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1014), .A2(KEYINPUT110), .A3(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1065), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT52), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1068), .A2(new_n1066), .A3(G8), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT110), .B1(new_n1014), .B2(new_n1070), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1074), .A2(new_n1075), .B1(G1976), .B2(new_n782), .ZN(new_n1076));
  INV_X1    g651(.A(G1976), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT52), .B1(G288), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT49), .ZN(new_n1080));
  INV_X1    g655(.A(G1981), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n587), .A2(new_n541), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n592), .A2(new_n589), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n1083), .B2(KEYINPUT111), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT111), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n592), .A2(new_n1085), .A3(new_n589), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1081), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n594), .A2(new_n591), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n585), .A2(new_n588), .A3(new_n589), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1088), .A2(new_n1089), .A3(G1981), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1080), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n590), .A2(new_n1081), .A3(new_n591), .A4(new_n594), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1086), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1085), .B1(new_n592), .B2(new_n589), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1093), .A2(new_n1094), .A3(new_n1082), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1092), .B(KEYINPUT49), .C1(new_n1095), .C2(new_n1081), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1073), .A2(new_n1079), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n976), .A2(new_n1002), .A3(new_n761), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n1102));
  INV_X1    g677(.A(G1961), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1101), .A2(new_n1102), .B1(new_n1038), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1000), .B1(G164), .B2(G1384), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n850), .A2(new_n998), .A3(new_n978), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(new_n969), .B2(new_n975), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1102), .A2(G2078), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1104), .A2(G301), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT125), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n461), .B1(new_n965), .B2(KEYINPUT124), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(KEYINPUT124), .B2(new_n965), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1002), .A2(new_n968), .A3(new_n1114), .A4(new_n1109), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1104), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(G171), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1104), .A2(new_n1118), .A3(G301), .A4(new_n1110), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1112), .A2(new_n1117), .A3(KEYINPUT54), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT55), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(G166), .B2(new_n1070), .ZN(new_n1122));
  NAND3_X1  g697(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G2090), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n976), .A2(new_n1125), .A3(new_n1008), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1971), .B1(new_n976), .B2(new_n1002), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1124), .B(G8), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n976), .A2(new_n1125), .A3(new_n1008), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1035), .B2(G1971), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1124), .B1(new_n1131), .B2(G8), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1134));
  AND3_X1   g709(.A1(new_n1104), .A2(G301), .A3(new_n1115), .ZN(new_n1135));
  AOI21_X1  g710(.A(G301), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1100), .A2(new_n1120), .A3(new_n1133), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(G286), .A2(G8), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n1140));
  AOI21_X1  g715(.A(G2084), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT113), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n976), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1108), .B2(G1966), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n976), .B2(new_n1141), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1140), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1145), .ZN(new_n1147));
  INV_X1    g722(.A(G1966), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n977), .B2(new_n1107), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1147), .A2(new_n1149), .A3(KEYINPUT121), .A4(new_n1143), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1139), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1146), .A2(G168), .A3(new_n1150), .ZN(new_n1152));
  OAI21_X1  g727(.A(G8), .B1(KEYINPUT122), .B2(KEYINPUT51), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(KEYINPUT122), .B2(KEYINPUT51), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(G8), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1156));
  AOI21_X1  g731(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1151), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1138), .A2(new_n1159), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1062), .A2(new_n1064), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1151), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1152), .A2(new_n1154), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT62), .B1(new_n1166), .B2(new_n1151), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1076), .A2(new_n1078), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1168));
  AND4_X1   g743(.A1(new_n1073), .A2(new_n1168), .A3(new_n1133), .A4(new_n1136), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1165), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  OAI211_X1 g745(.A(G8), .B(G168), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1168), .A2(new_n1133), .A3(new_n1073), .A4(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT114), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1174), .A2(KEYINPUT63), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1173), .B(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n782), .A2(new_n1077), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1177), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1098), .B1(new_n1178), .B2(new_n1090), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1073), .A2(new_n1079), .A3(new_n1099), .A4(new_n1129), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1179), .A2(new_n1180), .A3(KEYINPUT112), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT112), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1170), .A2(new_n1176), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n993), .B1(new_n1161), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n981), .A2(new_n982), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT46), .ZN(new_n1187));
  INV_X1    g762(.A(new_n985), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n981), .B1(new_n729), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT47), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n1192));
  OR2_X1    g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1194));
  NOR2_X1   g769(.A1(G290), .A2(G1986), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n981), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1196), .ZN(new_n1197));
  AOI22_X1  g772(.A1(new_n981), .A2(new_n991), .B1(new_n1197), .B2(KEYINPUT48), .ZN(new_n1198));
  OR2_X1    g773(.A1(new_n1197), .A2(KEYINPUT48), .ZN(new_n1199));
  OAI22_X1  g774(.A1(new_n987), .A2(new_n990), .B1(G2067), .B2(new_n696), .ZN(new_n1200));
  AOI22_X1  g775(.A1(new_n1198), .A2(new_n1199), .B1(new_n981), .B2(new_n1200), .ZN(new_n1201));
  AND3_X1   g776(.A1(new_n1193), .A2(new_n1194), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1185), .A2(new_n1202), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g778(.A(G319), .B1(new_n656), .B2(new_n657), .ZN(new_n1205));
  NOR3_X1   g779(.A1(G229), .A2(G227), .A3(new_n1205), .ZN(new_n1206));
  OAI211_X1 g780(.A(new_n875), .B(new_n1206), .C1(new_n958), .C2(new_n960), .ZN(G225));
  INV_X1    g781(.A(G225), .ZN(G308));
endmodule


