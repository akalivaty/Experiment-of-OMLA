//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT13), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT91), .ZN(new_n204));
  INV_X1    g003(.A(G8gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(G15gat), .A2(G22gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT90), .ZN(new_n208));
  NAND2_X1  g007(.A1(G15gat), .A2(G22gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n209), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT90), .B1(new_n211), .B2(new_n206), .ZN(new_n212));
  INV_X1    g011(.A(G1gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n210), .A2(new_n212), .B1(KEYINPUT16), .B2(new_n213), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n204), .B(new_n205), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n210), .A2(new_n212), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(KEYINPUT16), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n221));
  NAND2_X1  g020(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n214), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G50gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G43gat), .ZN(new_n226));
  INV_X1    g025(.A(G43gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G50gat), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT15), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G29gat), .ZN(new_n230));
  INV_X1    g029(.A(G36gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT14), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT14), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G29gat), .B2(G36gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT88), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT88), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G29gat), .A2(G36gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT89), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n236), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n228), .A3(KEYINPUT15), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n229), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n242), .B1(G29gat), .B2(G36gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(new_n234), .A3(new_n232), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n224), .A2(new_n246), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n217), .A2(new_n223), .B1(new_n243), .B2(new_n245), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n203), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT92), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g050(.A(KEYINPUT92), .B(new_n203), .C1(new_n247), .C2(new_n248), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT18), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT17), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n246), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n243), .A2(KEYINPUT17), .A3(new_n245), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n247), .B1(new_n258), .B2(new_n224), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n254), .B1(new_n259), .B2(new_n202), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n243), .A2(KEYINPUT17), .A3(new_n245), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT17), .B1(new_n243), .B2(new_n245), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n224), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n224), .A2(new_n246), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(new_n202), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n265), .A2(KEYINPUT18), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n253), .B1(new_n260), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT11), .B(G169gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(G197gat), .ZN(new_n269));
  XOR2_X1   g068(.A(G113gat), .B(G141gat), .Z(new_n270));
  XOR2_X1   g069(.A(new_n269), .B(new_n270), .Z(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT12), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n259), .A2(new_n254), .A3(new_n202), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n265), .A2(KEYINPUT18), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n274), .A2(new_n275), .B1(new_n251), .B2(new_n252), .ZN(new_n276));
  INV_X1    g075(.A(new_n272), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G85gat), .A2(G92gat), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n281), .B(KEYINPUT7), .Z(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT98), .ZN(new_n284));
  INV_X1    g083(.A(G85gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT97), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(G92gat), .ZN(new_n287));
  INV_X1    g086(.A(G92gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(KEYINPUT97), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n285), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G99gat), .ZN(new_n291));
  INV_X1    g090(.A(G106gat), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT8), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n284), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n288), .A2(KEYINPUT97), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n286), .A2(G92gat), .ZN(new_n296));
  AOI21_X1  g095(.A(G85gat), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT8), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n298), .B1(G99gat), .B2(G106gat), .ZN(new_n299));
  NOR3_X1   g098(.A1(new_n297), .A2(KEYINPUT98), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n283), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G99gat), .B(G106gat), .Z(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT98), .B1(new_n297), .B2(new_n299), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT97), .B(G92gat), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n284), .B(new_n293), .C1(new_n305), .C2(G85gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n302), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n283), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT95), .ZN(new_n310));
  INV_X1    g109(.A(G57gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(G64gat), .ZN(new_n312));
  INV_X1    g111(.A(G64gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(G57gat), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT94), .ZN(new_n316));
  OAI22_X1  g115(.A1(new_n312), .A2(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G71gat), .A2(G78gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT9), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(G71gat), .A2(G78gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(G71gat), .A2(G78gat), .ZN(new_n322));
  OAI22_X1  g121(.A1(new_n320), .A2(KEYINPUT94), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n310), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n313), .A2(G57gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n311), .A2(G64gat), .ZN(new_n326));
  AOI22_X1  g125(.A1(KEYINPUT94), .A2(new_n320), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OR2_X1    g126(.A1(G71gat), .A2(G78gat), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n318), .A2(new_n328), .B1(new_n315), .B2(new_n316), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT95), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n320), .B1(new_n312), .B2(new_n314), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT93), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT93), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n333), .B1(new_n328), .B2(new_n318), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n324), .A2(new_n330), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n303), .A2(new_n309), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n331), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n317), .A2(new_n323), .A3(new_n310), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT95), .B1(new_n327), .B2(new_n329), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n308), .B1(new_n307), .B2(new_n283), .ZN(new_n342));
  AOI211_X1 g141(.A(new_n302), .B(new_n282), .C1(new_n304), .C2(new_n306), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n337), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G230gat), .A2(G233gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G120gat), .B(G148gat), .ZN(new_n349));
  INV_X1    g148(.A(G176gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G204gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT96), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n341), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n336), .A2(KEYINPUT96), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n303), .A2(KEYINPUT99), .A3(new_n309), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT99), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(new_n342), .B2(new_n343), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n358), .A2(new_n359), .A3(new_n361), .A4(KEYINPUT10), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT10), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n337), .A2(new_n344), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT101), .B1(new_n365), .B2(new_n346), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT101), .ZN(new_n367));
  AOI211_X1 g166(.A(new_n367), .B(new_n347), .C1(new_n362), .C2(new_n364), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n348), .B(new_n354), .C1(new_n366), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n365), .A2(new_n346), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n348), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n353), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n280), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G127gat), .B(G155gat), .ZN(new_n376));
  INV_X1    g175(.A(G211gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n358), .A2(KEYINPUT21), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n224), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G183gat), .ZN(new_n381));
  INV_X1    g180(.A(G183gat), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n379), .A2(new_n382), .A3(new_n224), .ZN(new_n383));
  INV_X1    g182(.A(G231gat), .ZN(new_n384));
  INV_X1    g183(.A(G233gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n381), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n386), .B1(new_n381), .B2(new_n383), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n378), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n389), .ZN(new_n391));
  INV_X1    g190(.A(new_n378), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n387), .A3(new_n392), .ZN(new_n393));
  OR2_X1    g192(.A1(new_n336), .A2(KEYINPUT21), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n394), .B(new_n395), .Z(new_n396));
  AND3_X1   g195(.A1(new_n390), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n396), .B1(new_n390), .B2(new_n393), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n359), .A2(new_n361), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n400), .A2(new_n246), .ZN(new_n401));
  XOR2_X1   g200(.A(G190gat), .B(G218gat), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n400), .A2(new_n258), .B1(KEYINPUT100), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n401), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(G134gat), .B(G162gat), .Z(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n403), .A2(KEYINPUT100), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT41), .ZN(new_n410));
  INV_X1    g209(.A(G232gat), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n410), .B1(new_n411), .B2(new_n385), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n409), .B(new_n412), .Z(new_n413));
  INV_X1    g212(.A(new_n407), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n401), .A2(new_n404), .A3(new_n414), .A4(new_n405), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n408), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n413), .B1(new_n408), .B2(new_n415), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n399), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G190gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n382), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(G183gat), .A2(G190gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(KEYINPUT24), .A3(new_n424), .ZN(new_n425));
  OR2_X1    g224(.A1(new_n424), .A2(KEYINPUT24), .ZN(new_n426));
  NAND2_X1  g225(.A1(G169gat), .A2(G176gat), .ZN(new_n427));
  INV_X1    g226(.A(G169gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(new_n350), .A3(KEYINPUT23), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n425), .A2(new_n426), .A3(new_n427), .A4(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT23), .B1(new_n428), .B2(new_n350), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n430), .A2(KEYINPUT25), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT28), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT27), .B(G183gat), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT67), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n382), .A2(KEYINPUT27), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n422), .B1(new_n437), .B2(KEYINPUT67), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n433), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n434), .A2(KEYINPUT28), .A3(new_n422), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n439), .A2(new_n440), .B1(G183gat), .B2(G190gat), .ZN(new_n441));
  OR3_X1    g240(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n427), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n432), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n425), .A2(new_n426), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(KEYINPUT66), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT64), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n427), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n429), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT65), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n431), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n452), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT25), .B1(new_n447), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n445), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g257(.A(G127gat), .B(G134gat), .Z(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n460));
  XNOR2_X1  g259(.A(G113gat), .B(G120gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(KEYINPUT69), .B(KEYINPUT1), .Z(new_n463));
  XNOR2_X1  g262(.A(G127gat), .B(G134gat), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT68), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n460), .A2(new_n462), .A3(new_n463), .A4(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n459), .B1(KEYINPUT1), .B2(new_n461), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n467), .A2(KEYINPUT70), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT70), .B1(new_n467), .B2(new_n468), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n458), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(G227gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(new_n385), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n469), .A2(new_n470), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(new_n445), .A3(new_n457), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(G15gat), .B(G43gat), .Z(new_n480));
  XNOR2_X1  g279(.A(G71gat), .B(G99gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n476), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n475), .B1(new_n457), .B2(new_n445), .ZN(new_n485));
  OAI22_X1  g284(.A1(new_n484), .A2(new_n485), .B1(new_n473), .B2(new_n385), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(KEYINPUT71), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n474), .B1(new_n472), .B2(new_n476), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT71), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT34), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n477), .A2(KEYINPUT32), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(new_n488), .B2(new_n491), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n483), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n492), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n487), .B1(new_n486), .B2(KEYINPUT71), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT34), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n483), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n495), .A2(new_n502), .A3(KEYINPUT36), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT36), .B1(new_n495), .B2(new_n502), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G141gat), .B(G148gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT77), .ZN(new_n507));
  NAND2_X1  g306(.A1(G155gat), .A2(G162gat), .ZN(new_n508));
  INV_X1    g307(.A(G155gat), .ZN(new_n509));
  INV_X1    g308(.A(G162gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n508), .B1(new_n511), .B2(KEYINPUT2), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n508), .B(new_n511), .C1(new_n506), .C2(KEYINPUT2), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G218gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT22), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT72), .B(G211gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(new_n516), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT73), .ZN(new_n520));
  XNOR2_X1  g319(.A(G197gat), .B(G204gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n520), .B1(new_n519), .B2(new_n521), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n523), .A2(G211gat), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n519), .A2(new_n521), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT73), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n377), .B1(new_n527), .B2(new_n522), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n516), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT29), .ZN(new_n530));
  OAI21_X1  g329(.A(G211gat), .B1(new_n523), .B2(new_n524), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n527), .A2(new_n377), .A3(new_n522), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(G218gat), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT3), .B1(new_n534), .B2(KEYINPUT80), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT80), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n529), .A2(new_n536), .A3(new_n530), .A4(new_n533), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n515), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n529), .A2(new_n533), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT3), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n513), .A2(new_n540), .A3(new_n514), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n539), .B1(KEYINPUT29), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  OAI211_X1 g343(.A(G228gat), .B(G233gat), .C1(new_n538), .C2(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n534), .A2(new_n515), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n513), .A2(new_n514), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT3), .ZN(new_n548));
  NAND2_X1  g347(.A1(G228gat), .A2(G233gat), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n546), .A2(new_n548), .A3(new_n549), .A4(new_n543), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT31), .B(G50gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G78gat), .B(G106gat), .ZN(new_n554));
  INV_X1    g353(.A(G22gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n552), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n535), .A2(new_n537), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n544), .B1(new_n558), .B2(new_n547), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n557), .B(new_n550), .C1(new_n559), .C2(new_n549), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n553), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n556), .ZN(new_n562));
  INV_X1    g361(.A(new_n560), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n557), .B1(new_n545), .B2(new_n550), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n467), .A2(new_n468), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT4), .B1(new_n547), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT79), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT4), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n515), .B(new_n571), .C1(new_n469), .C2(new_n470), .ZN(new_n572));
  OAI211_X1 g371(.A(KEYINPUT79), .B(KEYINPUT4), .C1(new_n547), .C2(new_n567), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT5), .ZN(new_n575));
  NAND2_X1  g374(.A1(G225gat), .A2(G233gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n548), .A2(new_n567), .A3(new_n541), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n547), .B(new_n567), .ZN(new_n579));
  INV_X1    g378(.A(new_n576), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n575), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n515), .B(KEYINPUT4), .C1(new_n469), .C2(new_n470), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n547), .A2(new_n567), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n580), .A2(new_n571), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n577), .B(new_n582), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n578), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G1gat), .B(G29gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(G57gat), .B(G85gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT6), .ZN(new_n594));
  INV_X1    g393(.A(new_n592), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n578), .A2(new_n586), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n587), .A2(KEYINPUT6), .A3(new_n592), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G8gat), .B(G36gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G92gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT76), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(new_n313), .ZN(new_n604));
  NAND2_X1  g403(.A1(G226gat), .A2(G233gat), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n606), .B1(new_n458), .B2(new_n530), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n605), .B1(new_n445), .B2(new_n457), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(KEYINPUT74), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(KEYINPUT74), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n539), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n539), .B1(new_n607), .B2(new_n608), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n611), .A2(new_n612), .B1(new_n613), .B2(KEYINPUT75), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n458), .A2(new_n530), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n605), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n458), .A2(KEYINPUT74), .A3(new_n606), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n608), .A2(KEYINPUT74), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n616), .B(new_n612), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT75), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n604), .B1(new_n614), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n609), .A2(new_n610), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n623), .A2(KEYINPUT75), .A3(new_n612), .A4(new_n616), .ZN(new_n624));
  INV_X1    g423(.A(new_n604), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n613), .A2(KEYINPUT75), .ZN(new_n626));
  INV_X1    g425(.A(new_n619), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n624), .B(new_n625), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n622), .A2(KEYINPUT30), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n614), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT30), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n630), .A2(new_n631), .A3(new_n624), .A4(new_n625), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n600), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n505), .B1(new_n566), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT81), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT83), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n574), .A2(new_n577), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(new_n637), .B2(new_n580), .ZN(new_n638));
  AOI211_X1 g437(.A(KEYINPUT83), .B(new_n576), .C1(new_n574), .C2(new_n577), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n640), .B(KEYINPUT39), .C1(new_n580), .C2(new_n579), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(new_n638), .B2(new_n639), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT84), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n592), .B(KEYINPUT82), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n644), .B1(new_n643), .B2(new_n646), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n641), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT85), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(KEYINPUT40), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n629), .A2(new_n632), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n587), .A2(new_n645), .ZN(new_n654));
  INV_X1    g453(.A(new_n651), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n655), .B(new_n641), .C1(new_n647), .C2(new_n648), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n652), .A2(new_n653), .A3(new_n654), .A4(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n616), .B(new_n539), .C1(new_n617), .C2(new_n618), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n612), .B1(new_n607), .B2(new_n608), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(KEYINPUT37), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT38), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT37), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n624), .B(new_n663), .C1(new_n626), .C2(new_n627), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n662), .A2(new_n664), .A3(new_n604), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n654), .A2(new_n594), .A3(new_n596), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n598), .A2(KEYINPUT86), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT86), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n587), .A2(new_n668), .A3(KEYINPUT6), .A4(new_n592), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n628), .A2(new_n666), .A3(new_n667), .A4(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT87), .B1(new_n665), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n663), .B1(new_n630), .B2(new_n624), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n664), .A2(new_n604), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT38), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n662), .A2(new_n664), .A3(new_n604), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT87), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n675), .A2(new_n676), .A3(new_n677), .A4(new_n628), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n671), .A2(new_n674), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n657), .A2(new_n679), .A3(new_n566), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT81), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n505), .B(new_n681), .C1(new_n566), .C2(new_n633), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n635), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n495), .A2(new_n502), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n566), .A2(new_n633), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT35), .ZN(new_n686));
  INV_X1    g485(.A(new_n684), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(new_n561), .B2(new_n565), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n629), .A2(new_n632), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n675), .A2(KEYINPUT35), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  AOI211_X1 g491(.A(new_n375), .B(new_n421), .C1(new_n683), .C2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n600), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G1gat), .ZN(G1324gat));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n683), .A2(new_n692), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(new_n374), .A3(new_n420), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n698), .B2(new_n689), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n693), .A2(KEYINPUT102), .A3(new_n653), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT105), .B1(new_n701), .B2(new_n205), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n699), .A2(new_n700), .A3(new_n703), .A4(G8gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT16), .B(G8gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT103), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT104), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n708), .A2(KEYINPUT104), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n701), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT42), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n693), .A2(KEYINPUT42), .A3(new_n653), .A4(new_n708), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n705), .A2(new_n713), .A3(new_n714), .ZN(G1325gat));
  AOI21_X1  g514(.A(G15gat), .B1(new_n693), .B2(new_n684), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n698), .A2(new_n505), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n716), .B1(G15gat), .B2(new_n717), .ZN(G1326gat));
  AND2_X1   g517(.A1(new_n561), .A2(new_n565), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n693), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT43), .B(G22gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1327gat));
  AOI21_X1  g521(.A(new_n418), .B1(new_n683), .B2(new_n692), .ZN(new_n723));
  INV_X1    g522(.A(new_n399), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n375), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n230), .A3(new_n600), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT45), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n697), .A2(KEYINPUT44), .A3(new_n419), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731));
  INV_X1    g530(.A(new_n634), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n680), .A2(new_n732), .B1(new_n686), .B2(new_n691), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n733), .B2(new_n418), .ZN(new_n734));
  AND4_X1   g533(.A1(new_n600), .A2(new_n730), .A3(new_n725), .A4(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n729), .B1(new_n230), .B2(new_n735), .ZN(G1328gat));
  NOR3_X1   g535(.A1(new_n726), .A2(G36gat), .A3(new_n689), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  AND4_X1   g539(.A1(new_n653), .A2(new_n730), .A3(new_n725), .A4(new_n734), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n739), .B(new_n740), .C1(new_n231), .C2(new_n741), .ZN(G1329gat));
  OAI21_X1  g541(.A(new_n227), .B1(new_n726), .B2(new_n687), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n730), .A2(new_n725), .A3(new_n734), .ZN(new_n744));
  INV_X1    g543(.A(new_n505), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G43gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n743), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g547(.A1(KEYINPUT107), .A2(KEYINPUT48), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT107), .A2(KEYINPUT48), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT108), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n730), .A2(new_n734), .A3(new_n719), .A4(new_n725), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n752), .A2(G50gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n719), .A2(new_n225), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT106), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n727), .A2(new_n755), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n749), .B(new_n751), .C1(new_n753), .C2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n751), .ZN(new_n758));
  AOI22_X1  g557(.A1(new_n752), .A2(G50gat), .B1(new_n727), .B2(new_n755), .ZN(new_n759));
  INV_X1    g558(.A(new_n749), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n757), .A2(new_n761), .ZN(G1331gat));
  OAI211_X1 g561(.A(new_n280), .B(new_n418), .C1(new_n397), .C2(new_n398), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n689), .B1(new_n651), .B2(new_n649), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n656), .A2(new_n654), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n719), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n634), .B1(new_n767), .B2(new_n679), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n566), .A2(new_n689), .A3(new_n684), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n769), .A2(new_n690), .B1(new_n685), .B2(KEYINPUT35), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n373), .B(new_n764), .C1(new_n768), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n599), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(new_n311), .ZN(G1332gat));
  NAND2_X1  g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n373), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n680), .A2(new_n732), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n692), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT109), .B1(new_n779), .B2(new_n764), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n653), .B(new_n774), .C1(new_n776), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(KEYINPUT110), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n771), .A2(new_n775), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n779), .A2(KEYINPUT109), .A3(new_n764), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n689), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n783), .B1(new_n786), .B2(new_n774), .ZN(new_n787));
  OAI22_X1  g586(.A1(new_n782), .A2(new_n787), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n781), .A2(KEYINPUT110), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n786), .A2(new_n783), .A3(new_n774), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT49), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n789), .A2(new_n790), .A3(new_n791), .A4(new_n313), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n788), .A2(new_n792), .ZN(G1333gat));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n784), .A2(new_n785), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n745), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G71gat), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT111), .B1(new_n771), .B2(new_n687), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n779), .A2(new_n799), .A3(new_n684), .A4(new_n764), .ZN(new_n800));
  AOI21_X1  g599(.A(G71gat), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n794), .B1(new_n797), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(G71gat), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n804), .B1(new_n795), .B2(new_n745), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n805), .A2(new_n801), .A3(KEYINPUT50), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n803), .A2(new_n806), .ZN(G1334gat));
  NAND2_X1  g606(.A1(new_n795), .A2(new_n719), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g608(.A1(new_n724), .A2(new_n279), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n730), .A2(new_n734), .A3(new_n373), .A4(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G85gat), .B1(new_n811), .B2(new_n599), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n418), .B1(new_n778), .B2(new_n692), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n813), .A2(KEYINPUT51), .A3(new_n810), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT51), .B1(new_n813), .B2(new_n810), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n777), .A2(new_n599), .A3(G85gat), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT112), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n812), .B1(new_n816), .B2(new_n818), .ZN(G1336gat));
  OAI21_X1  g618(.A(new_n305), .B1(new_n811), .B2(new_n689), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n777), .A2(G92gat), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n653), .B(new_n821), .C1(new_n814), .C2(new_n815), .ZN(new_n822));
  NAND2_X1  g621(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n820), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT114), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n820), .A2(new_n826), .A3(new_n822), .A4(new_n823), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1337gat));
  XOR2_X1   g629(.A(KEYINPUT115), .B(G99gat), .Z(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n811), .B2(new_n505), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n373), .B(new_n684), .C1(new_n814), .C2(new_n815), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n831), .B2(new_n833), .ZN(G1338gat));
  NAND2_X1  g633(.A1(KEYINPUT116), .A2(G106gat), .ZN(new_n835));
  OR2_X1    g634(.A1(KEYINPUT116), .A2(G106gat), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n835), .B(new_n836), .C1(new_n811), .C2(new_n566), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n719), .A2(new_n292), .A3(new_n373), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n838), .B(KEYINPUT117), .Z(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n814), .B2(new_n815), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT53), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n837), .B(new_n843), .C1(new_n816), .C2(new_n838), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(G1339gat));
  NOR2_X1   g644(.A1(new_n763), .A2(new_n373), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT54), .B1(new_n365), .B2(new_n346), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n370), .A2(new_n367), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n347), .B1(new_n362), .B2(new_n364), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT101), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n849), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n354), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n848), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n366), .A2(new_n368), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT55), .B(new_n855), .C1(new_n858), .C2(new_n849), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n857), .A2(new_n369), .A3(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n271), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n247), .A2(new_n248), .ZN(new_n862));
  OAI22_X1  g661(.A1(new_n259), .A2(new_n202), .B1(new_n862), .B2(new_n203), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n276), .A2(new_n277), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n416), .B2(new_n417), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n857), .A2(new_n279), .A3(new_n369), .A4(new_n859), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n373), .A2(new_n864), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n373), .A2(new_n864), .A3(KEYINPUT118), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n867), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n866), .B1(new_n872), .B2(new_n418), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n847), .B1(new_n873), .B2(new_n724), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n874), .A2(new_n600), .A3(new_n769), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n279), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n373), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(G120gat), .ZN(G1341gat));
  NAND3_X1  g678(.A1(new_n875), .A2(G127gat), .A3(new_n724), .ZN(new_n880));
  XOR2_X1   g679(.A(new_n880), .B(KEYINPUT119), .Z(new_n881));
  AOI21_X1  g680(.A(G127gat), .B1(new_n875), .B2(new_n724), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(G1342gat));
  NAND2_X1  g682(.A1(new_n875), .A2(new_n419), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(G134gat), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT56), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(G134gat), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1343gat));
  NOR3_X1   g687(.A1(new_n745), .A2(new_n599), .A3(new_n653), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n419), .B1(new_n867), .B2(new_n868), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n399), .B1(new_n890), .B2(new_n866), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n847), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n719), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XOR2_X1   g694(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n896));
  AOI21_X1  g695(.A(new_n896), .B1(new_n874), .B2(new_n719), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n889), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G141gat), .B1(new_n898), .B2(new_n280), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n874), .A2(new_n719), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n889), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n901), .A2(G141gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n899), .B1(new_n280), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT58), .ZN(G1344gat));
  OR3_X1    g703(.A1(new_n901), .A2(G148gat), .A3(new_n777), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n872), .A2(new_n418), .ZN(new_n907));
  INV_X1    g706(.A(new_n866), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n724), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n719), .B(new_n896), .C1(new_n909), .C2(new_n846), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT121), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n893), .A2(new_n894), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n874), .A2(new_n913), .A3(new_n719), .A4(new_n896), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n373), .A3(new_n889), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n906), .B1(new_n916), .B2(G148gat), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n373), .B(new_n889), .C1(new_n895), .C2(new_n897), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n918), .A2(new_n906), .A3(G148gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n905), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g721(.A(KEYINPUT122), .B(new_n905), .C1(new_n917), .C2(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1345gat));
  OR3_X1    g723(.A1(new_n898), .A2(new_n509), .A3(new_n399), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n900), .A2(new_n724), .A3(new_n889), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n926), .B1(new_n509), .B2(new_n927), .ZN(G1346gat));
  OR3_X1    g727(.A1(new_n898), .A2(new_n510), .A3(new_n418), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n510), .B1(new_n901), .B2(new_n418), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(G1347gat));
  NOR2_X1   g730(.A1(new_n689), .A2(new_n600), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n874), .A2(new_n688), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT123), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n874), .A2(new_n688), .A3(new_n932), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(G169gat), .B1(new_n938), .B2(new_n280), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n933), .A2(new_n428), .A3(new_n279), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1348gat));
  NAND2_X1  g740(.A1(new_n934), .A2(new_n937), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(G176gat), .A3(new_n373), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(KEYINPUT124), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(KEYINPUT124), .ZN(new_n945));
  AOI21_X1  g744(.A(G176gat), .B1(new_n933), .B2(new_n373), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(G1349gat));
  OAI21_X1  g746(.A(G183gat), .B1(new_n938), .B2(new_n399), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n933), .A2(new_n724), .A3(new_n434), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n952), .B(G190gat), .C1(new_n938), .C2(new_n418), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n418), .B1(new_n934), .B2(new_n937), .ZN(new_n954));
  OAI21_X1  g753(.A(KEYINPUT125), .B1(new_n954), .B2(new_n422), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n933), .A2(new_n422), .A3(new_n419), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n953), .A2(KEYINPUT61), .A3(new_n955), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(G1351gat));
  AND2_X1   g760(.A1(new_n505), .A2(new_n932), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n915), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(new_n279), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G197gat), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n900), .A2(new_n962), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n966), .A2(G197gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n965), .B1(new_n280), .B2(new_n967), .ZN(G1352gat));
  NOR3_X1   g767(.A1(new_n966), .A2(G204gat), .A3(new_n777), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT62), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n915), .A2(new_n373), .A3(new_n962), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n352), .B2(new_n971), .ZN(G1353gat));
  NAND2_X1  g771(.A1(new_n963), .A2(new_n724), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n724), .A2(new_n518), .ZN(new_n976));
  OAI22_X1  g775(.A1(new_n974), .A2(new_n975), .B1(new_n966), .B2(new_n976), .ZN(G1354gat));
  OAI21_X1  g776(.A(new_n516), .B1(new_n966), .B2(new_n418), .ZN(new_n978));
  XOR2_X1   g777(.A(new_n978), .B(KEYINPUT126), .Z(new_n979));
  NAND2_X1  g778(.A1(new_n419), .A2(G218gat), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT127), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n979), .B1(new_n963), .B2(new_n981), .ZN(G1355gat));
endmodule


