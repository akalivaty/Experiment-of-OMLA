

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595;

  NOR2_X2 U325 ( .A1(n589), .A2(n575), .ZN(n577) );
  XNOR2_X1 U326 ( .A(n294), .B(KEYINPUT13), .ZN(n327) );
  XNOR2_X2 U327 ( .A(G57GAT), .B(KEYINPUT69), .ZN(n294) );
  XOR2_X1 U328 ( .A(n434), .B(n433), .Z(n293) );
  NOR2_X1 U329 ( .A1(n567), .A2(n366), .ZN(n368) );
  INV_X1 U330 ( .A(KEYINPUT80), .ZN(n437) );
  INV_X1 U331 ( .A(n380), .ZN(n321) );
  XNOR2_X1 U332 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U333 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U334 ( .A(n440), .B(n439), .ZN(n444) );
  XNOR2_X1 U335 ( .A(n315), .B(n309), .ZN(n310) );
  XNOR2_X1 U336 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U337 ( .A(n311), .B(n310), .ZN(n345) );
  XNOR2_X1 U338 ( .A(n412), .B(KEYINPUT65), .ZN(n580) );
  XNOR2_X1 U339 ( .A(n483), .B(KEYINPUT38), .ZN(n511) );
  XNOR2_X1 U340 ( .A(n458), .B(KEYINPUT58), .ZN(n459) );
  XNOR2_X1 U341 ( .A(n488), .B(KEYINPUT39), .ZN(n489) );
  XNOR2_X1 U342 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  XNOR2_X1 U343 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  XOR2_X1 U344 ( .A(G120GAT), .B(G71GAT), .Z(n434) );
  XNOR2_X1 U345 ( .A(n327), .B(n434), .ZN(n296) );
  AND2_X1 U346 ( .A1(G230GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n299) );
  INV_X1 U348 ( .A(n299), .ZN(n297) );
  NAND2_X1 U349 ( .A1(n297), .A2(KEYINPUT71), .ZN(n301) );
  INV_X1 U350 ( .A(KEYINPUT71), .ZN(n298) );
  NAND2_X1 U351 ( .A1(n299), .A2(n298), .ZN(n300) );
  NAND2_X1 U352 ( .A1(n301), .A2(n300), .ZN(n304) );
  XNOR2_X1 U353 ( .A(G78GAT), .B(G204GAT), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n302), .B(G148GAT), .ZN(n419) );
  XNOR2_X1 U355 ( .A(n419), .B(KEYINPUT31), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U357 ( .A(G176GAT), .B(G64GAT), .Z(n377) );
  XOR2_X1 U358 ( .A(n305), .B(n377), .Z(n311) );
  XOR2_X1 U359 ( .A(KEYINPUT70), .B(G92GAT), .Z(n307) );
  XNOR2_X1 U360 ( .A(G99GAT), .B(G85GAT), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U362 ( .A(G106GAT), .B(n308), .Z(n315) );
  XNOR2_X1 U363 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n309) );
  XNOR2_X1 U364 ( .A(KEYINPUT41), .B(n345), .ZN(n560) );
  XOR2_X1 U365 ( .A(n560), .B(KEYINPUT108), .Z(n543) );
  XOR2_X1 U366 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n313) );
  XNOR2_X1 U367 ( .A(KEYINPUT67), .B(KEYINPUT11), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n326) );
  XOR2_X1 U370 ( .A(G29GAT), .B(G43GAT), .Z(n317) );
  XNOR2_X1 U371 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n357) );
  XOR2_X1 U373 ( .A(n357), .B(KEYINPUT9), .Z(n319) );
  NAND2_X1 U374 ( .A1(G232GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U375 ( .A(n319), .B(n318), .ZN(n324) );
  XOR2_X1 U376 ( .A(G50GAT), .B(G162GAT), .Z(n423) );
  XOR2_X1 U377 ( .A(G134GAT), .B(KEYINPUT74), .Z(n402) );
  XNOR2_X1 U378 ( .A(n423), .B(n402), .ZN(n322) );
  XNOR2_X1 U379 ( .A(G36GAT), .B(G190GAT), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n320), .B(G218GAT), .ZN(n380) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n567) );
  XNOR2_X1 U382 ( .A(KEYINPUT75), .B(n567), .ZN(n551) );
  XNOR2_X1 U383 ( .A(KEYINPUT36), .B(n551), .ZN(n461) );
  XOR2_X1 U384 ( .A(G8GAT), .B(G183GAT), .Z(n375) );
  XOR2_X1 U385 ( .A(n375), .B(n327), .Z(n329) );
  XNOR2_X1 U386 ( .A(G71GAT), .B(G127GAT), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n334) );
  XNOR2_X1 U388 ( .A(G15GAT), .B(G22GAT), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n330), .B(G1GAT), .ZN(n356) );
  XOR2_X1 U390 ( .A(n356), .B(KEYINPUT77), .Z(n332) );
  NAND2_X1 U391 ( .A1(G231GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U393 ( .A(n334), .B(n333), .Z(n342) );
  XOR2_X1 U394 ( .A(G64GAT), .B(G211GAT), .Z(n336) );
  XNOR2_X1 U395 ( .A(G155GAT), .B(G78GAT), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U397 ( .A(KEYINPUT12), .B(KEYINPUT76), .Z(n338) );
  XNOR2_X1 U398 ( .A(KEYINPUT14), .B(KEYINPUT15), .ZN(n337) );
  XNOR2_X1 U399 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n589) );
  NOR2_X1 U402 ( .A1(n461), .A2(n589), .ZN(n344) );
  XNOR2_X1 U403 ( .A(KEYINPUT45), .B(KEYINPUT66), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n346) );
  BUF_X1 U405 ( .A(n345), .Z(n586) );
  NAND2_X1 U406 ( .A1(n346), .A2(n586), .ZN(n347) );
  XNOR2_X1 U407 ( .A(KEYINPUT115), .B(n347), .ZN(n362) );
  XOR2_X1 U408 ( .A(G50GAT), .B(G36GAT), .Z(n349) );
  NAND2_X1 U409 ( .A1(G229GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n361) );
  XOR2_X1 U411 ( .A(KEYINPUT29), .B(G8GAT), .Z(n351) );
  XNOR2_X1 U412 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U414 ( .A(G141GAT), .B(G197GAT), .Z(n353) );
  XNOR2_X1 U415 ( .A(G169GAT), .B(G113GAT), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U417 ( .A(n355), .B(n354), .Z(n359) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U419 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U420 ( .A(n361), .B(n360), .Z(n581) );
  NAND2_X1 U421 ( .A1(n362), .A2(n581), .ZN(n370) );
  INV_X1 U422 ( .A(n581), .ZN(n558) );
  NAND2_X1 U423 ( .A1(n560), .A2(n558), .ZN(n364) );
  INV_X1 U424 ( .A(KEYINPUT46), .ZN(n363) );
  XOR2_X1 U425 ( .A(n364), .B(n363), .Z(n365) );
  NAND2_X1 U426 ( .A1(n365), .A2(n589), .ZN(n366) );
  XNOR2_X1 U427 ( .A(KEYINPUT114), .B(KEYINPUT47), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n369) );
  NAND2_X1 U429 ( .A1(n370), .A2(n369), .ZN(n372) );
  XOR2_X1 U430 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n555) );
  XOR2_X1 U432 ( .A(G92GAT), .B(KEYINPUT94), .Z(n374) );
  NAND2_X1 U433 ( .A1(G226GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n374), .B(n373), .ZN(n376) );
  XOR2_X1 U435 ( .A(n376), .B(n375), .Z(n379) );
  XNOR2_X1 U436 ( .A(G204GAT), .B(n377), .ZN(n378) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n381) );
  XOR2_X1 U438 ( .A(n381), .B(n380), .Z(n387) );
  XOR2_X1 U439 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n383) );
  XNOR2_X1 U440 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n383), .B(n382), .ZN(n436) );
  XOR2_X1 U442 ( .A(G211GAT), .B(KEYINPUT86), .Z(n385) );
  XNOR2_X1 U443 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n422) );
  XNOR2_X1 U445 ( .A(n436), .B(n422), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n387), .B(n386), .ZN(n529) );
  NOR2_X1 U447 ( .A1(n555), .A2(n529), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n388), .B(KEYINPUT54), .ZN(n411) );
  XOR2_X1 U449 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n390) );
  XNOR2_X1 U450 ( .A(KEYINPUT4), .B(KEYINPUT6), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n390), .B(n389), .ZN(n410) );
  XOR2_X1 U452 ( .A(G85GAT), .B(G162GAT), .Z(n392) );
  XNOR2_X1 U453 ( .A(G120GAT), .B(G148GAT), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U455 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n394) );
  XNOR2_X1 U456 ( .A(G1GAT), .B(G57GAT), .ZN(n393) );
  XNOR2_X1 U457 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U458 ( .A(n396), .B(n395), .Z(n408) );
  XOR2_X1 U459 ( .A(KEYINPUT87), .B(G155GAT), .Z(n398) );
  XNOR2_X1 U460 ( .A(G141GAT), .B(KEYINPUT88), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n400) );
  XOR2_X1 U462 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n399) );
  XNOR2_X1 U463 ( .A(n400), .B(n399), .ZN(n431) );
  INV_X1 U464 ( .A(n431), .ZN(n406) );
  XNOR2_X1 U465 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n401) );
  XNOR2_X1 U466 ( .A(n401), .B(G127GAT), .ZN(n433) );
  XOR2_X1 U467 ( .A(n402), .B(n433), .Z(n404) );
  NAND2_X1 U468 ( .A1(G225GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U469 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U470 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n410), .B(n409), .ZN(n484) );
  XNOR2_X1 U473 ( .A(G29GAT), .B(n484), .ZN(n556) );
  NAND2_X1 U474 ( .A1(n411), .A2(n556), .ZN(n412) );
  XOR2_X1 U475 ( .A(KEYINPUT84), .B(KEYINPUT90), .Z(n414) );
  XNOR2_X1 U476 ( .A(KEYINPUT22), .B(KEYINPUT89), .ZN(n413) );
  XNOR2_X1 U477 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U478 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n416) );
  XNOR2_X1 U479 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n415) );
  XNOR2_X1 U480 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U481 ( .A(n418), .B(n417), .Z(n429) );
  XOR2_X1 U482 ( .A(n419), .B(KEYINPUT85), .Z(n421) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n427) );
  XOR2_X1 U485 ( .A(n422), .B(G106GAT), .Z(n425) );
  XNOR2_X1 U486 ( .A(G218GAT), .B(n423), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U489 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n471) );
  NAND2_X1 U491 ( .A1(n580), .A2(n471), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n432), .B(KEYINPUT55), .ZN(n453) );
  NAND2_X1 U493 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n293), .B(n435), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n436), .B(KEYINPUT79), .ZN(n438) );
  XOR2_X1 U496 ( .A(G190GAT), .B(G134GAT), .Z(n442) );
  XNOR2_X1 U497 ( .A(G43GAT), .B(G99GAT), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n452) );
  XOR2_X1 U500 ( .A(KEYINPUT83), .B(KEYINPUT78), .Z(n446) );
  XNOR2_X1 U501 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U503 ( .A(G176GAT), .B(G183GAT), .Z(n448) );
  XNOR2_X1 U504 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U506 ( .A(n450), .B(n449), .Z(n451) );
  XNOR2_X1 U507 ( .A(n452), .B(n451), .ZN(n541) );
  AND2_X2 U508 ( .A1(n453), .A2(n541), .ZN(n454) );
  XNOR2_X2 U509 ( .A(n454), .B(KEYINPUT121), .ZN(n575) );
  NOR2_X1 U510 ( .A1(n543), .A2(n575), .ZN(n457) );
  XNOR2_X1 U511 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n455) );
  XNOR2_X1 U512 ( .A(n455), .B(G176GAT), .ZN(n456) );
  XNOR2_X1 U513 ( .A(n457), .B(n456), .ZN(G1349GAT) );
  NOR2_X1 U514 ( .A1(n551), .A2(n575), .ZN(n460) );
  INV_X1 U515 ( .A(G190GAT), .ZN(n458) );
  XOR2_X1 U516 ( .A(n529), .B(KEYINPUT27), .Z(n473) );
  XNOR2_X1 U517 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n463) );
  NOR2_X1 U518 ( .A1(n541), .A2(n471), .ZN(n462) );
  XNOR2_X1 U519 ( .A(n463), .B(n462), .ZN(n579) );
  NAND2_X1 U520 ( .A1(n473), .A2(n579), .ZN(n554) );
  XNOR2_X1 U521 ( .A(n554), .B(KEYINPUT97), .ZN(n468) );
  INV_X1 U522 ( .A(n529), .ZN(n505) );
  NAND2_X1 U523 ( .A1(n505), .A2(n541), .ZN(n464) );
  NAND2_X1 U524 ( .A1(n464), .A2(n471), .ZN(n465) );
  XNOR2_X1 U525 ( .A(n465), .B(KEYINPUT25), .ZN(n466) );
  XNOR2_X1 U526 ( .A(KEYINPUT98), .B(n466), .ZN(n467) );
  NOR2_X1 U527 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U528 ( .A(KEYINPUT99), .B(n469), .ZN(n470) );
  NAND2_X1 U529 ( .A1(n470), .A2(n556), .ZN(n476) );
  XOR2_X1 U530 ( .A(n471), .B(KEYINPUT28), .Z(n510) );
  NOR2_X1 U531 ( .A1(n556), .A2(n510), .ZN(n472) );
  NAND2_X1 U532 ( .A1(n473), .A2(n472), .ZN(n539) );
  XNOR2_X1 U533 ( .A(n539), .B(KEYINPUT95), .ZN(n474) );
  INV_X1 U534 ( .A(n541), .ZN(n532) );
  NAND2_X1 U535 ( .A1(n474), .A2(n532), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U537 ( .A(KEYINPUT100), .B(n477), .ZN(n493) );
  NAND2_X1 U538 ( .A1(n493), .A2(n589), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n478), .B(KEYINPUT104), .ZN(n479) );
  NOR2_X1 U540 ( .A1(n461), .A2(n479), .ZN(n481) );
  XOR2_X1 U541 ( .A(KEYINPUT105), .B(KEYINPUT37), .Z(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(n524) );
  NAND2_X1 U543 ( .A1(n586), .A2(n558), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n482), .B(KEYINPUT72), .ZN(n494) );
  NOR2_X1 U545 ( .A1(n524), .A2(n494), .ZN(n483) );
  NOR2_X1 U546 ( .A1(G29GAT), .A2(n511), .ZN(n487) );
  INV_X1 U547 ( .A(n511), .ZN(n485) );
  NOR2_X1 U548 ( .A1(n485), .A2(n484), .ZN(n486) );
  NOR2_X1 U549 ( .A1(n487), .A2(n486), .ZN(n490) );
  INV_X1 U550 ( .A(KEYINPUT106), .ZN(n488) );
  INV_X1 U551 ( .A(n589), .ZN(n564) );
  NAND2_X1 U552 ( .A1(n551), .A2(n564), .ZN(n491) );
  XOR2_X1 U553 ( .A(KEYINPUT16), .B(n491), .Z(n492) );
  NAND2_X1 U554 ( .A1(n493), .A2(n492), .ZN(n513) );
  OR2_X1 U555 ( .A1(n494), .A2(n513), .ZN(n503) );
  NOR2_X1 U556 ( .A1(n556), .A2(n503), .ZN(n496) );
  XNOR2_X1 U557 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G1GAT), .B(n497), .ZN(G1324GAT) );
  NOR2_X1 U560 ( .A1(n529), .A2(n503), .ZN(n498) );
  XOR2_X1 U561 ( .A(G8GAT), .B(n498), .Z(G1325GAT) );
  NOR2_X1 U562 ( .A1(n503), .A2(n532), .ZN(n502) );
  XOR2_X1 U563 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n500) );
  XNOR2_X1 U564 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(G1326GAT) );
  INV_X1 U567 ( .A(n510), .ZN(n535) );
  NOR2_X1 U568 ( .A1(n535), .A2(n503), .ZN(n504) );
  XOR2_X1 U569 ( .A(G22GAT), .B(n504), .Z(G1327GAT) );
  XOR2_X1 U570 ( .A(G36GAT), .B(KEYINPUT107), .Z(n507) );
  NAND2_X1 U571 ( .A1(n511), .A2(n505), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(G1329GAT) );
  NAND2_X1 U573 ( .A1(n511), .A2(n541), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(KEYINPUT40), .ZN(n509) );
  XNOR2_X1 U575 ( .A(G43GAT), .B(n509), .ZN(G1330GAT) );
  NAND2_X1 U576 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U578 ( .A1(n543), .A2(n558), .ZN(n525) );
  INV_X1 U579 ( .A(n513), .ZN(n514) );
  NAND2_X1 U580 ( .A1(n525), .A2(n514), .ZN(n519) );
  NOR2_X1 U581 ( .A1(n556), .A2(n519), .ZN(n515) );
  XOR2_X1 U582 ( .A(n515), .B(KEYINPUT42), .Z(n516) );
  XNOR2_X1 U583 ( .A(G57GAT), .B(n516), .ZN(G1332GAT) );
  NOR2_X1 U584 ( .A1(n529), .A2(n519), .ZN(n517) );
  XOR2_X1 U585 ( .A(G64GAT), .B(n517), .Z(G1333GAT) );
  NOR2_X1 U586 ( .A1(n532), .A2(n519), .ZN(n518) );
  XOR2_X1 U587 ( .A(G71GAT), .B(n518), .Z(G1334GAT) );
  NOR2_X1 U588 ( .A1(n519), .A2(n535), .ZN(n523) );
  XOR2_X1 U589 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n521) );
  XNOR2_X1 U590 ( .A(G78GAT), .B(KEYINPUT110), .ZN(n520) );
  XNOR2_X1 U591 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U592 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  INV_X1 U593 ( .A(n524), .ZN(n526) );
  NAND2_X1 U594 ( .A1(n526), .A2(n525), .ZN(n534) );
  NOR2_X1 U595 ( .A1(n556), .A2(n534), .ZN(n528) );
  XNOR2_X1 U596 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n527) );
  XNOR2_X1 U597 ( .A(n528), .B(n527), .ZN(G1336GAT) );
  NOR2_X1 U598 ( .A1(n529), .A2(n534), .ZN(n530) );
  XOR2_X1 U599 ( .A(KEYINPUT112), .B(n530), .Z(n531) );
  XNOR2_X1 U600 ( .A(G92GAT), .B(n531), .ZN(G1337GAT) );
  NOR2_X1 U601 ( .A1(n532), .A2(n534), .ZN(n533) );
  XOR2_X1 U602 ( .A(G99GAT), .B(n533), .Z(G1338GAT) );
  NOR2_X1 U603 ( .A1(n535), .A2(n534), .ZN(n537) );
  XNOR2_X1 U604 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U606 ( .A(G106GAT), .B(n538), .ZN(G1339GAT) );
  NOR2_X1 U607 ( .A1(n555), .A2(n539), .ZN(n540) );
  NAND2_X1 U608 ( .A1(n541), .A2(n540), .ZN(n550) );
  NOR2_X1 U609 ( .A1(n581), .A2(n550), .ZN(n542) );
  XOR2_X1 U610 ( .A(G113GAT), .B(n542), .Z(G1340GAT) );
  NOR2_X1 U611 ( .A1(n543), .A2(n550), .ZN(n545) );
  XNOR2_X1 U612 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U614 ( .A(G120GAT), .B(n546), .ZN(G1341GAT) );
  NOR2_X1 U615 ( .A1(n589), .A2(n550), .ZN(n548) );
  XNOR2_X1 U616 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U618 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  NOR2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  OR2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n557) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n568) );
  AND2_X1 U624 ( .A1(n558), .A2(n568), .ZN(n559) );
  XOR2_X1 U625 ( .A(G141GAT), .B(n559), .Z(G1344GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n562) );
  NAND2_X1 U627 ( .A1(n568), .A2(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(n563), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n568), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT118), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G155GAT), .B(n566), .ZN(G1346GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n570) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G162GAT), .B(n571), .ZN(G1347GAT) );
  NOR2_X1 U637 ( .A1(n581), .A2(n575), .ZN(n574) );
  XNOR2_X1 U638 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(KEYINPUT123), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1348GAT) );
  INV_X1 U641 ( .A(KEYINPUT124), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n593) );
  NOR2_X1 U645 ( .A1(n593), .A2(n581), .ZN(n585) );
  XOR2_X1 U646 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n583) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n593), .ZN(n588) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n593), .ZN(n591) );
  XNOR2_X1 U654 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G211GAT), .B(n592), .ZN(G1354GAT) );
  NOR2_X1 U657 ( .A1(n461), .A2(n593), .ZN(n594) );
  XOR2_X1 U658 ( .A(KEYINPUT62), .B(n594), .Z(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

