//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1097, new_n1098;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT68), .B(G2105), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n463), .A2(G2105), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n469), .A2(new_n471), .B1(G101), .B2(new_n472), .ZN(new_n473));
  AND3_X1   g048(.A1(new_n463), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT69), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n464), .B2(new_n475), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n476), .A2(KEYINPUT70), .A3(G137), .A4(new_n470), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n463), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n480), .B1(new_n465), .B2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n465), .A2(G2104), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n470), .A2(G137), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n478), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n473), .A2(new_n477), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G160));
  INV_X1    g062(.A(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n476), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT71), .Z(new_n492));
  NOR2_X1   g067(.A1(new_n483), .A2(new_n470), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G124), .ZN(new_n494));
  NOR2_X1   g069(.A1(G100), .A2(G2105), .ZN(new_n495));
  XNOR2_X1  g070(.A(new_n495), .B(KEYINPUT72), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n492), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G162));
  AND2_X1   g074(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(KEYINPUT4), .B(G138), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  AND2_X1   g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT73), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(new_n476), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n479), .B(new_n503), .C1(new_n481), .C2(new_n482), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n510));
  OAI21_X1  g085(.A(G138), .B1(new_n500), .B2(new_n501), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(new_n467), .ZN(new_n512));
  OR2_X1    g087(.A1(G102), .A2(G2105), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT74), .B(G114), .ZN(new_n514));
  OAI211_X1 g089(.A(G2104), .B(new_n513), .C1(new_n514), .C2(new_n488), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n506), .A2(new_n509), .A3(new_n512), .A4(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(G164));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT75), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT5), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G543), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n526), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n518), .ZN(new_n529));
  INV_X1    g104(.A(G88), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OR3_X1    g106(.A1(new_n521), .A2(KEYINPUT76), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT76), .B1(new_n521), .B2(new_n531), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(G166));
  NAND2_X1  g109(.A1(new_n519), .A2(G51), .ZN(new_n535));
  INV_X1    g110(.A(G89), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n523), .A2(new_n525), .ZN(new_n537));
  NAND2_X1  g112(.A1(G63), .A2(G651), .ZN(new_n538));
  OAI221_X1 g113(.A(new_n535), .B1(new_n536), .B2(new_n529), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT77), .ZN(new_n541));
  XOR2_X1   g116(.A(new_n541), .B(KEYINPUT7), .Z(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G168));
  AOI22_X1  g118(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n528), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n518), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n529), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n545), .A2(new_n549), .ZN(G171));
  INV_X1    g125(.A(new_n529), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(G81), .B1(G43), .B2(new_n519), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n528), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT78), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n547), .A2(KEYINPUT9), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n547), .B2(new_n563), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT79), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n526), .B(KEYINPUT80), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(G91), .B2(new_n551), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n567), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  XNOR2_X1  g149(.A(G168), .B(KEYINPUT81), .ZN(G286));
  AND2_X1   g150(.A1(new_n532), .A2(new_n533), .ZN(G303));
  NAND2_X1  g151(.A1(new_n551), .A2(G87), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n519), .A2(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  AOI22_X1  g155(.A1(new_n526), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n528), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n529), .A2(new_n583), .B1(new_n547), .B2(new_n584), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n582), .A2(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n528), .ZN(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n529), .A2(new_n589), .B1(new_n547), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  AND2_X1   g168(.A1(G301), .A2(G868), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n569), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G79), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n522), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n596), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  OAI221_X1 g176(.A(KEYINPUT83), .B1(new_n599), .B2(new_n522), .C1(new_n569), .C2(new_n597), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n601), .A2(G651), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n519), .A2(G54), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n551), .A2(G92), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT10), .Z(new_n606));
  NAND3_X1  g181(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n595), .B1(new_n608), .B2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(KEYINPUT82), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(KEYINPUT82), .B2(new_n594), .ZN(G284));
  OAI21_X1  g186(.A(new_n610), .B1(KEYINPUT82), .B2(new_n594), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G299), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(G868), .B2(new_n614), .ZN(G297));
  OAI21_X1  g190(.A(new_n613), .B1(G868), .B2(new_n614), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n608), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n608), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n490), .A2(G135), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n493), .A2(G123), .ZN(new_n624));
  OAI221_X1 g199(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n470), .C2(G111), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  NAND3_X1  g202(.A1(new_n488), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n627), .A2(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT15), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2435), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n637));
  XOR2_X1   g212(.A(G2443), .B(G2446), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G1341), .B(G1348), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n642), .B(new_n643), .Z(new_n644));
  AND2_X1   g219(.A1(new_n644), .A2(G14), .ZN(G401));
  XOR2_X1   g220(.A(G2072), .B(G2078), .Z(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2067), .B(G2678), .Z(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2096), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(G2100), .Z(new_n654));
  INV_X1    g229(.A(KEYINPUT17), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n648), .B2(new_n649), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n651), .B1(new_n650), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n660), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n669), .B(new_n670), .C1(new_n668), .C2(new_n667), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G1981), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT86), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT21), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n672), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT85), .B(G1986), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n677), .B(new_n678), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G229));
  NOR2_X1   g255(.A1(G16), .A2(G22), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(G166), .B2(G16), .ZN(new_n682));
  INV_X1    g257(.A(G1971), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  MUX2_X1   g259(.A(G6), .B(G305), .S(G16), .Z(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT32), .B(G1981), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT88), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G23), .ZN(new_n690));
  INV_X1    g265(.A(G288), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT33), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1976), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n684), .A2(new_n688), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT34), .Z(new_n696));
  NOR2_X1   g271(.A1(G25), .A2(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n490), .A2(G131), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n493), .A2(G119), .ZN(new_n699));
  OAI221_X1 g274(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n470), .C2(G107), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n697), .B1(new_n702), .B2(G29), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT87), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT35), .B(G1991), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G1986), .ZN(new_n708));
  NOR2_X1   g283(.A1(G16), .A2(G24), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n592), .B2(G16), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n707), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n696), .B(new_n712), .C1(new_n708), .C2(new_n711), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT36), .Z(new_n714));
  INV_X1    g289(.A(KEYINPUT94), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n716), .A2(G35), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n715), .B(new_n717), .C1(new_n498), .C2(G29), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n715), .B2(new_n717), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT29), .B(G2090), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(G115), .A2(G2104), .ZN(new_n722));
  INV_X1    g297(.A(G127), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n467), .B2(new_n723), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n490), .A2(G139), .B1(new_n471), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT25), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  MUX2_X1   g303(.A(G33), .B(new_n728), .S(G29), .Z(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(G2072), .Z(new_n730));
  INV_X1    g305(.A(G1966), .ZN(new_n731));
  NOR2_X1   g306(.A1(G16), .A2(G21), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G168), .B2(G16), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n730), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n689), .A2(G19), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n555), .B2(new_n689), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(G1341), .Z(new_n738));
  NAND2_X1  g313(.A1(G171), .A2(G16), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G5), .B2(G16), .ZN(new_n740));
  INV_X1    g315(.A(G1961), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT93), .B(KEYINPUT30), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G28), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n740), .A2(new_n741), .B1(new_n716), .B2(new_n743), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n738), .B(new_n744), .C1(G1966), .C2(new_n733), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n721), .A2(new_n735), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n740), .A2(new_n741), .ZN(new_n747));
  INV_X1    g322(.A(G11), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(KEYINPUT31), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n748), .A2(KEYINPUT31), .ZN(new_n750));
  NOR3_X1   g325(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(KEYINPUT24), .A2(G34), .ZN(new_n752));
  NAND2_X1  g327(.A1(KEYINPUT24), .A2(G34), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n752), .A2(new_n716), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G160), .B2(new_n716), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n755), .A2(G2084), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(G2084), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n716), .A2(G27), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G164), .B2(new_n716), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(G2078), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n756), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n746), .A2(new_n751), .A3(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n626), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n762), .B1(G29), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n689), .A2(G4), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n608), .B2(new_n689), .ZN(new_n766));
  INV_X1    g341(.A(G1348), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n493), .A2(G129), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n472), .A2(G105), .ZN(new_n770));
  INV_X1    g345(.A(G141), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n769), .B(new_n770), .C1(new_n771), .C2(new_n489), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT91), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT26), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G29), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n778), .B(KEYINPUT92), .C1(G29), .C2(G32), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(KEYINPUT92), .B2(new_n778), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT27), .B(G1996), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G2078), .B2(new_n759), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n493), .A2(G128), .ZN(new_n784));
  OAI221_X1 g359(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n470), .C2(G116), .ZN(new_n785));
  INV_X1    g360(.A(G140), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n784), .B(new_n785), .C1(new_n786), .C2(new_n489), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G29), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n716), .A2(G26), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT89), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT28), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT90), .B(G2067), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n689), .A2(KEYINPUT23), .A3(G20), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT23), .ZN(new_n796));
  INV_X1    g371(.A(G20), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G16), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n795), .B(new_n798), .C1(new_n614), .C2(new_n689), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT95), .B(G1956), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n783), .A2(new_n794), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n764), .A2(new_n768), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(KEYINPUT96), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT96), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n764), .A2(new_n806), .A3(new_n768), .A4(new_n803), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n714), .B1(new_n805), .B2(new_n807), .ZN(G311));
  INV_X1    g383(.A(G311), .ZN(G150));
  NAND2_X1  g384(.A1(G80), .A2(G543), .ZN(new_n810));
  INV_X1    g385(.A(G67), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n537), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT97), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n813), .A2(G651), .ZN(new_n814));
  INV_X1    g389(.A(G93), .ZN(new_n815));
  INV_X1    g390(.A(G55), .ZN(new_n816));
  OAI22_X1  g391(.A1(new_n529), .A2(new_n815), .B1(new_n547), .B2(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G860), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT37), .Z(new_n820));
  NOR2_X1   g395(.A1(new_n607), .A2(new_n617), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT38), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT39), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n555), .B1(new_n818), .B2(KEYINPUT98), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n814), .A2(new_n817), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n825), .A2(new_n826), .A3(new_n555), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n823), .B(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n820), .B1(new_n831), .B2(G860), .ZN(G145));
  NAND2_X1  g407(.A1(new_n490), .A2(G142), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT100), .Z(new_n834));
  OAI221_X1 g409(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n470), .C2(G118), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n493), .A2(G130), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n701), .B(new_n629), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT101), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n728), .A2(KEYINPUT99), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G164), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n777), .B(new_n787), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n840), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n626), .B(new_n486), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n498), .B(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G37), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n847), .B1(new_n840), .B2(new_n844), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n844), .B2(new_n839), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g428(.A1(new_n818), .A2(G868), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n608), .A2(G299), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n607), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(KEYINPUT41), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT102), .B1(new_n614), .B2(new_n607), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(new_n857), .B2(KEYINPUT102), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n859), .B1(new_n861), .B2(KEYINPUT41), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n830), .B(new_n619), .Z(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(G166), .B(G305), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n592), .B(G288), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT42), .Z(new_n868));
  OAI221_X1 g443(.A(new_n864), .B1(new_n863), .B2(new_n858), .C1(new_n868), .C2(KEYINPUT103), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(KEYINPUT103), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n869), .B(new_n870), .Z(new_n871));
  AOI21_X1  g446(.A(new_n854), .B1(new_n871), .B2(G868), .ZN(G295));
  AOI21_X1  g447(.A(new_n854), .B1(new_n871), .B2(G868), .ZN(G331));
  NOR3_X1   g448(.A1(new_n539), .A2(G171), .A3(new_n542), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(G286), .B2(G171), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n830), .B(new_n875), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n876), .B(new_n859), .C1(KEYINPUT41), .C2(new_n861), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n857), .B2(new_n876), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n879));
  INV_X1    g454(.A(new_n867), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n879), .B1(new_n878), .B2(new_n880), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n876), .A2(KEYINPUT41), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(new_n861), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n858), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n867), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n885), .A2(KEYINPUT105), .A3(new_n867), .A4(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n883), .A2(new_n891), .A3(new_n892), .A4(new_n849), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n878), .A2(new_n880), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT104), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n878), .A2(new_n880), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n849), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT43), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n883), .A2(new_n891), .A3(KEYINPUT43), .A4(new_n849), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n892), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  MUX2_X1   g478(.A(new_n900), .B(new_n903), .S(KEYINPUT44), .Z(G397));
  INV_X1    g479(.A(G1384), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT45), .B1(new_n516), .B2(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n473), .A2(new_n477), .A3(G40), .A4(new_n485), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n909), .A2(G1996), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n777), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT107), .ZN(new_n912));
  INV_X1    g487(.A(new_n909), .ZN(new_n913));
  INV_X1    g488(.A(new_n777), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n914), .A2(G1996), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n787), .B(G2067), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n912), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n701), .B(new_n706), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n918), .B1(new_n909), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n592), .A2(new_n708), .ZN(new_n921));
  XOR2_X1   g496(.A(new_n921), .B(KEYINPUT106), .Z(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(new_n708), .B2(new_n592), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n920), .B1(new_n913), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT55), .ZN(new_n928));
  INV_X1    g503(.A(G8), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n928), .B1(G166), .B2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(G303), .A2(KEYINPUT109), .A3(KEYINPUT55), .A4(G8), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n516), .A2(new_n905), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n516), .A2(KEYINPUT45), .A3(new_n905), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n908), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n683), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(KEYINPUT108), .A3(new_n683), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n933), .A2(KEYINPUT50), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT50), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n516), .A2(new_n943), .A3(new_n905), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n908), .A3(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n945), .A2(G2090), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n940), .A2(new_n941), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n932), .A2(G8), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n933), .A2(new_n907), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(new_n929), .ZN(new_n950));
  INV_X1    g525(.A(G1976), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n950), .B1(new_n951), .B2(G288), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n952), .A2(KEYINPUT52), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n691), .A2(G1976), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n952), .A2(KEYINPUT52), .A3(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(G305), .B(G1981), .ZN(new_n956));
  NOR2_X1   g531(.A1(KEYINPUT110), .A2(KEYINPUT49), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n956), .B(new_n957), .Z(new_n958));
  AOI211_X1 g533(.A(new_n953), .B(new_n955), .C1(new_n950), .C2(new_n958), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n948), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n932), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n946), .A2(new_n938), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n962), .A2(KEYINPUT112), .ZN(new_n963));
  OAI21_X1  g538(.A(G8), .B1(new_n962), .B2(KEYINPUT112), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n942), .A2(new_n908), .A3(new_n944), .ZN(new_n967));
  INV_X1    g542(.A(G2084), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n967), .A2(new_n968), .B1(new_n937), .B2(new_n731), .ZN(new_n969));
  OAI21_X1  g544(.A(G8), .B1(new_n539), .B2(new_n542), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT119), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT120), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n974), .B(new_n971), .C1(new_n969), .C2(new_n929), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT122), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n942), .A2(new_n968), .A3(new_n908), .A4(new_n944), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n516), .A2(KEYINPUT45), .A3(new_n905), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n979), .A2(new_n906), .A3(new_n907), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n980), .B2(G1966), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(G8), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n982), .A2(KEYINPUT122), .A3(new_n974), .A4(new_n971), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n977), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n971), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n937), .A2(new_n731), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n929), .B1(new_n986), .B2(new_n978), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT121), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n982), .A2(KEYINPUT121), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n974), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n973), .B(KEYINPUT123), .C1(new_n984), .C2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n981), .A2(new_n988), .A3(G8), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n971), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n987), .A2(new_n988), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT51), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(new_n977), .A3(new_n983), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT123), .B1(new_n998), .B2(new_n973), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT62), .B1(new_n993), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n1001));
  OR3_X1    g576(.A1(new_n937), .A2(new_n1001), .A3(G2078), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n945), .A2(new_n741), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n937), .B2(G2078), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(G171), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n973), .B1(new_n984), .B2(new_n991), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT123), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT62), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(new_n992), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1000), .A2(new_n1007), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(new_n992), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1002), .A2(G301), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1006), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT124), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT60), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n933), .A2(new_n907), .A3(G2067), .ZN(new_n1021));
  AOI211_X1 g596(.A(new_n1020), .B(new_n1021), .C1(new_n945), .C2(new_n767), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1019), .B1(new_n1022), .B2(new_n607), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n945), .A2(new_n767), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1021), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(KEYINPUT60), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT117), .B1(new_n1026), .B2(new_n608), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1022), .A2(new_n1028), .A3(new_n607), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1026), .A2(KEYINPUT118), .A3(new_n608), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1023), .A2(new_n1027), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1021), .B1(new_n945), .B2(new_n767), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1032), .A2(KEYINPUT60), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT58), .B(G1341), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n937), .A2(G1996), .B1(new_n949), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(new_n1037), .A3(new_n555), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1038), .B(KEYINPUT59), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT56), .B(G2072), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n980), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n935), .A2(new_n908), .A3(new_n936), .A4(new_n1041), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT115), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT114), .B(G1956), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1042), .A2(new_n1044), .B1(new_n945), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT57), .B1(new_n564), .B2(new_n565), .ZN(new_n1047));
  AOI22_X1  g622(.A1(G299), .A2(KEYINPUT57), .B1(new_n572), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT61), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1049), .A2(KEYINPUT61), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1034), .A2(new_n1039), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1032), .A2(new_n607), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1049), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1018), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1016), .A2(KEYINPUT124), .A3(new_n1017), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1006), .B(KEYINPUT125), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(KEYINPUT54), .A3(new_n1015), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1014), .A2(new_n1056), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n966), .B1(new_n1013), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n982), .A2(G286), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1062), .B(KEYINPUT113), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n947), .A2(G8), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(new_n961), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n960), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n960), .A2(new_n965), .A3(new_n1063), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1067), .B1(new_n1068), .B2(KEYINPUT63), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n959), .A2(G8), .A3(new_n932), .A4(new_n947), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n958), .A2(new_n950), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1071), .A2(new_n951), .A3(new_n691), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(G1981), .B2(G305), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(KEYINPUT111), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n950), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1069), .A2(new_n1070), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n924), .B1(new_n1061), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n918), .A2(new_n706), .A3(new_n702), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n787), .A2(G2067), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n909), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1080), .B(KEYINPUT126), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n910), .A2(KEYINPUT46), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n913), .B1(new_n916), .B2(new_n914), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n910), .A2(KEYINPUT46), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(KEYINPUT47), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n922), .A2(new_n909), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1087), .B(KEYINPUT48), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1081), .B(new_n1086), .C1(new_n920), .C2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1077), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT127), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT127), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1077), .A2(new_n1093), .A3(new_n1090), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g670(.A1(G401), .A2(G227), .ZN(new_n1097));
  AND2_X1   g671(.A1(new_n1097), .A2(new_n852), .ZN(new_n1098));
  NAND4_X1  g672(.A1(new_n900), .A2(new_n1098), .A3(G319), .A4(new_n679), .ZN(G225));
  INV_X1    g673(.A(G225), .ZN(G308));
endmodule


