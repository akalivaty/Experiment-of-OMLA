

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764;

  XNOR2_X1 U372 ( .A(n561), .B(KEYINPUT32), .ZN(n599) );
  INV_X1 U373 ( .A(G953), .ZN(n430) );
  XNOR2_X2 U374 ( .A(KEYINPUT64), .B(G143), .ZN(n414) );
  NAND2_X2 U375 ( .A1(n635), .A2(n754), .ZN(n399) );
  OR2_X1 U376 ( .A1(n548), .A2(n547), .ZN(n550) );
  NAND2_X1 U377 ( .A1(n407), .A2(n405), .ZN(n528) );
  AND2_X1 U378 ( .A1(n409), .A2(n408), .ZN(n407) );
  XNOR2_X1 U379 ( .A(n536), .B(n535), .ZN(n684) );
  XNOR2_X1 U380 ( .A(n550), .B(n549), .ZN(n564) );
  NAND2_X1 U381 ( .A1(n356), .A2(n368), .ZN(n610) );
  OR2_X2 U382 ( .A1(n399), .A2(n729), .ZN(n359) );
  XNOR2_X2 U383 ( .A(n753), .B(G146), .ZN(n374) );
  XNOR2_X2 U384 ( .A(n437), .B(n436), .ZN(n753) );
  XNOR2_X2 U385 ( .A(n469), .B(n357), .ZN(n437) );
  NAND2_X1 U386 ( .A1(n599), .A2(n565), .ZN(n569) );
  XNOR2_X1 U387 ( .A(n591), .B(KEYINPUT38), .ZN(n708) );
  NAND2_X1 U388 ( .A1(n591), .A2(n519), .ZN(n372) );
  AND2_X1 U389 ( .A1(n396), .A2(n390), .ZN(n389) );
  NAND2_X1 U390 ( .A1(n393), .A2(n391), .ZN(n390) );
  NAND2_X1 U391 ( .A1(n388), .A2(n360), .ZN(n387) );
  XNOR2_X1 U392 ( .A(n438), .B(G125), .ZN(n449) );
  NOR2_X1 U393 ( .A1(n569), .A2(KEYINPUT65), .ZN(n567) );
  AND2_X1 U394 ( .A1(n532), .A2(n531), .ZN(n558) );
  XNOR2_X1 U395 ( .A(n449), .B(n448), .ZN(n476) );
  INV_X1 U396 ( .A(KEYINPUT10), .ZN(n448) );
  XOR2_X1 U397 ( .A(G137), .B(G140), .Z(n474) );
  XNOR2_X1 U398 ( .A(n518), .B(n517), .ZN(n706) );
  INV_X1 U399 ( .A(KEYINPUT33), .ZN(n517) );
  NOR2_X1 U400 ( .A1(n533), .A2(n551), .ZN(n518) );
  XNOR2_X1 U401 ( .A(n508), .B(n507), .ZN(n562) );
  OR2_X1 U402 ( .A1(n661), .A2(G902), .ZN(n508) );
  XNOR2_X1 U403 ( .A(KEYINPUT3), .B(G119), .ZN(n422) );
  XNOR2_X1 U404 ( .A(n382), .B(n381), .ZN(n433) );
  XNOR2_X1 U405 ( .A(G104), .B(G101), .ZN(n382) );
  XNOR2_X1 U406 ( .A(G110), .B(G107), .ZN(n381) );
  XNOR2_X1 U407 ( .A(n386), .B(n385), .ZN(n723) );
  XNOR2_X1 U408 ( .A(KEYINPUT41), .B(KEYINPUT104), .ZN(n385) );
  NAND2_X1 U409 ( .A1(n714), .A2(n711), .ZN(n386) );
  AND2_X1 U410 ( .A1(n589), .A2(n593), .ZN(n380) );
  NOR2_X1 U411 ( .A1(n410), .A2(n358), .ZN(n409) );
  NOR2_X1 U412 ( .A1(n534), .A2(n526), .ZN(n410) );
  NOR2_X1 U413 ( .A1(n655), .A2(n426), .ZN(n428) );
  XNOR2_X1 U414 ( .A(n489), .B(n488), .ZN(n514) );
  OR2_X1 U415 ( .A1(n545), .A2(n541), .ZN(n596) );
  AND2_X2 U416 ( .A1(n400), .A2(n359), .ZN(n746) );
  NAND2_X1 U417 ( .A1(n404), .A2(n401), .ZN(n400) );
  NAND2_X1 U418 ( .A1(n403), .A2(n402), .ZN(n401) );
  XNOR2_X1 U419 ( .A(n640), .B(KEYINPUT87), .ZN(n745) );
  NAND2_X1 U420 ( .A1(n395), .A2(n394), .ZN(n393) );
  NAND2_X1 U421 ( .A1(n392), .A2(n604), .ZN(n391) );
  OR2_X1 U422 ( .A1(n603), .A2(KEYINPUT79), .ZN(n392) );
  INV_X1 U423 ( .A(KEYINPUT79), .ZN(n394) );
  AND2_X1 U424 ( .A1(n398), .A2(n397), .ZN(n612) );
  NAND2_X1 U425 ( .A1(n389), .A2(n387), .ZN(n397) );
  NOR2_X1 U426 ( .A1(G237), .A2(G953), .ZN(n442) );
  INV_X1 U427 ( .A(KEYINPUT69), .ZN(n435) );
  XNOR2_X1 U428 ( .A(G113), .B(G143), .ZN(n451) );
  XNOR2_X1 U429 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n416) );
  XNOR2_X1 U430 ( .A(n621), .B(KEYINPUT103), .ZN(n714) );
  INV_X1 U431 ( .A(n605), .ZN(n375) );
  BUF_X1 U432 ( .A(n562), .Z(n537) );
  XNOR2_X1 U433 ( .A(n476), .B(n475), .ZN(n751) );
  XNOR2_X1 U434 ( .A(G119), .B(G128), .ZN(n478) );
  XOR2_X1 U435 ( .A(G107), .B(G122), .Z(n460) );
  INV_X1 U436 ( .A(G128), .ZN(n413) );
  INV_X1 U437 ( .A(KEYINPUT80), .ZN(n402) );
  NAND2_X1 U438 ( .A1(n384), .A2(n729), .ZN(n383) );
  NAND2_X1 U439 ( .A1(n376), .A2(n707), .ZN(n587) );
  NAND2_X1 U440 ( .A1(n370), .A2(n369), .ZN(n368) );
  NOR2_X1 U441 ( .A1(n519), .A2(n585), .ZN(n369) );
  XNOR2_X1 U442 ( .A(n562), .B(n377), .ZN(n376) );
  INV_X1 U443 ( .A(KEYINPUT100), .ZN(n377) );
  XNOR2_X1 U444 ( .A(KEYINPUT16), .B(G122), .ZN(n421) );
  NAND2_X1 U445 ( .A1(n399), .A2(n730), .ZN(n731) );
  AND2_X1 U446 ( .A1(n622), .A2(n723), .ZN(n623) );
  XNOR2_X1 U447 ( .A(n378), .B(n598), .ZN(n624) );
  NAND2_X1 U448 ( .A1(n406), .A2(KEYINPUT34), .ZN(n405) );
  NAND2_X1 U449 ( .A1(n560), .A2(n411), .ZN(n561) );
  NAND2_X1 U450 ( .A1(n622), .A2(n610), .ZN(n678) );
  XNOR2_X1 U451 ( .A(n596), .B(n473), .ZN(n680) );
  XNOR2_X1 U452 ( .A(n737), .B(n740), .ZN(n741) );
  AND2_X1 U453 ( .A1(n590), .A2(n589), .ZN(n351) );
  OR2_X1 U454 ( .A1(n678), .A2(n713), .ZN(n352) );
  AND2_X1 U455 ( .A1(n754), .A2(n426), .ZN(n353) );
  NOR2_X1 U456 ( .A1(n376), .A2(n592), .ZN(n354) );
  INV_X1 U457 ( .A(G146), .ZN(n438) );
  AND2_X1 U458 ( .A1(n429), .A2(G210), .ZN(n355) );
  AND2_X1 U459 ( .A1(n372), .A2(n371), .ZN(n356) );
  XOR2_X1 U460 ( .A(KEYINPUT68), .B(KEYINPUT4), .Z(n357) );
  XOR2_X1 U461 ( .A(n601), .B(KEYINPUT77), .Z(n358) );
  AND2_X1 U462 ( .A1(n604), .A2(n394), .ZN(n360) );
  AND2_X1 U463 ( .A1(n534), .A2(n526), .ZN(n361) );
  XNOR2_X1 U464 ( .A(n525), .B(KEYINPUT0), .ZN(n548) );
  NOR2_X1 U465 ( .A1(n680), .A2(n605), .ZN(n362) );
  OR2_X1 U466 ( .A1(n761), .A2(KEYINPUT44), .ZN(n363) );
  XOR2_X1 U467 ( .A(n543), .B(KEYINPUT99), .Z(n364) );
  AND2_X1 U468 ( .A1(n603), .A2(KEYINPUT79), .ZN(n365) );
  XOR2_X1 U469 ( .A(n678), .B(n611), .Z(n366) );
  AND2_X1 U470 ( .A1(n754), .A2(KEYINPUT80), .ZN(n367) );
  XNOR2_X1 U471 ( .A(KEYINPUT15), .B(G902), .ZN(n636) );
  NAND2_X1 U472 ( .A1(n370), .A2(n707), .ZN(n373) );
  INV_X1 U473 ( .A(n591), .ZN(n370) );
  NAND2_X1 U474 ( .A1(n585), .A2(n519), .ZN(n371) );
  NOR2_X1 U475 ( .A1(n613), .A2(n373), .ZN(n616) );
  NAND2_X1 U476 ( .A1(n353), .A2(n635), .ZN(n403) );
  NAND2_X1 U477 ( .A1(n367), .A2(n635), .ZN(n384) );
  XNOR2_X1 U478 ( .A(n399), .B(KEYINPUT78), .ZN(n690) );
  XNOR2_X1 U479 ( .A(n374), .B(n506), .ZN(n661) );
  XNOR2_X1 U480 ( .A(n374), .B(n439), .ZN(n737) );
  NAND2_X1 U481 ( .A1(n376), .A2(n375), .ZN(n607) );
  NOR2_X1 U482 ( .A1(n624), .A2(n764), .ZN(n625) );
  NAND2_X1 U483 ( .A1(n379), .A2(n597), .ZN(n378) );
  INV_X1 U484 ( .A(n631), .ZN(n379) );
  NAND2_X1 U485 ( .A1(n590), .A2(n380), .ZN(n595) );
  NAND2_X1 U486 ( .A1(n383), .A2(n426), .ZN(n404) );
  XNOR2_X2 U487 ( .A(n574), .B(KEYINPUT45), .ZN(n635) );
  NAND2_X1 U488 ( .A1(n351), .A2(n603), .ZN(n677) );
  INV_X1 U489 ( .A(n351), .ZN(n388) );
  INV_X1 U490 ( .A(n604), .ZN(n395) );
  NAND2_X1 U491 ( .A1(n351), .A2(n365), .ZN(n396) );
  NAND2_X1 U492 ( .A1(n352), .A2(n366), .ZN(n398) );
  INV_X1 U493 ( .A(n706), .ZN(n406) );
  NAND2_X1 U494 ( .A1(n706), .A2(n361), .ZN(n408) );
  BUF_X1 U495 ( .A(n706), .Z(n724) );
  AND2_X1 U496 ( .A1(n617), .A2(n514), .ZN(n411) );
  AND2_X1 U497 ( .A1(n490), .A2(G217), .ZN(n412) );
  INV_X1 U498 ( .A(KEYINPUT65), .ZN(n566) );
  INV_X1 U499 ( .A(n474), .ZN(n475) );
  XNOR2_X1 U500 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U501 ( .A(n456), .B(n455), .ZN(n645) );
  XNOR2_X1 U502 ( .A(KEYINPUT31), .B(KEYINPUT91), .ZN(n535) );
  XNOR2_X2 U503 ( .A(n414), .B(n413), .ZN(n469) );
  INV_X1 U504 ( .A(n437), .ZN(n420) );
  NAND2_X1 U505 ( .A1(n430), .A2(G224), .ZN(n415) );
  XNOR2_X1 U506 ( .A(n415), .B(KEYINPUT76), .ZN(n418) );
  XNOR2_X1 U507 ( .A(n449), .B(n416), .ZN(n417) );
  XNOR2_X1 U508 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U509 ( .A(n420), .B(n419), .ZN(n425) );
  XNOR2_X1 U510 ( .A(n433), .B(n421), .ZN(n424) );
  XNOR2_X1 U511 ( .A(G116), .B(G113), .ZN(n423) );
  XNOR2_X1 U512 ( .A(n423), .B(n422), .ZN(n504) );
  XNOR2_X1 U513 ( .A(n424), .B(n504), .ZN(n580) );
  XNOR2_X1 U514 ( .A(n425), .B(n580), .ZN(n655) );
  INV_X1 U515 ( .A(n636), .ZN(n426) );
  INV_X1 U516 ( .A(G902), .ZN(n485) );
  INV_X1 U517 ( .A(G237), .ZN(n427) );
  NAND2_X1 U518 ( .A1(n485), .A2(n427), .ZN(n429) );
  XNOR2_X2 U519 ( .A(n428), .B(n355), .ZN(n591) );
  AND2_X1 U520 ( .A1(n429), .A2(G214), .ZN(n585) );
  INV_X1 U521 ( .A(n585), .ZN(n707) );
  XOR2_X1 U522 ( .A(n474), .B(KEYINPUT75), .Z(n432) );
  NAND2_X1 U523 ( .A1(G227), .A2(n430), .ZN(n431) );
  XNOR2_X1 U524 ( .A(n432), .B(n431), .ZN(n434) );
  XNOR2_X1 U525 ( .A(n434), .B(n433), .ZN(n439) );
  XNOR2_X1 U526 ( .A(n435), .B(G131), .ZN(n450) );
  XNOR2_X1 U527 ( .A(n450), .B(G134), .ZN(n436) );
  OR2_X2 U528 ( .A1(n737), .A2(G902), .ZN(n440) );
  XNOR2_X2 U529 ( .A(n440), .B(G469), .ZN(n538) );
  INV_X1 U530 ( .A(KEYINPUT1), .ZN(n441) );
  XNOR2_X1 U531 ( .A(n538), .B(n441), .ZN(n515) );
  INV_X1 U532 ( .A(n515), .ZN(n553) );
  XNOR2_X1 U533 ( .A(KEYINPUT74), .B(n442), .ZN(n500) );
  NAND2_X1 U534 ( .A1(n500), .A2(G214), .ZN(n446) );
  XOR2_X1 U535 ( .A(KEYINPUT92), .B(KEYINPUT11), .Z(n444) );
  XNOR2_X1 U536 ( .A(G140), .B(KEYINPUT93), .ZN(n443) );
  XNOR2_X1 U537 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U538 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U539 ( .A(n447), .B(KEYINPUT12), .Z(n456) );
  XNOR2_X1 U540 ( .A(n450), .B(n476), .ZN(n454) );
  XOR2_X1 U541 ( .A(G104), .B(G122), .Z(n452) );
  XNOR2_X1 U542 ( .A(n452), .B(n451), .ZN(n453) );
  NAND2_X1 U543 ( .A1(n645), .A2(n485), .ZN(n458) );
  XNOR2_X1 U544 ( .A(KEYINPUT13), .B(G475), .ZN(n457) );
  XNOR2_X1 U545 ( .A(n458), .B(n457), .ZN(n545) );
  XNOR2_X1 U546 ( .A(G116), .B(G134), .ZN(n459) );
  XNOR2_X1 U547 ( .A(n460), .B(n459), .ZN(n464) );
  XOR2_X1 U548 ( .A(KEYINPUT94), .B(KEYINPUT7), .Z(n462) );
  XNOR2_X1 U549 ( .A(KEYINPUT9), .B(KEYINPUT95), .ZN(n461) );
  XNOR2_X1 U550 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U551 ( .A(n464), .B(n463), .Z(n467) );
  NAND2_X1 U552 ( .A1(G234), .A2(n430), .ZN(n465) );
  XOR2_X1 U553 ( .A(KEYINPUT8), .B(n465), .Z(n477) );
  NAND2_X1 U554 ( .A1(G217), .A2(n477), .ZN(n466) );
  XNOR2_X1 U555 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U556 ( .A(n469), .B(n468), .ZN(n748) );
  NAND2_X1 U557 ( .A1(n748), .A2(n485), .ZN(n472) );
  XNOR2_X1 U558 ( .A(G478), .B(KEYINPUT97), .ZN(n470) );
  XNOR2_X1 U559 ( .A(n470), .B(KEYINPUT96), .ZN(n471) );
  XNOR2_X1 U560 ( .A(n472), .B(n471), .ZN(n544) );
  INV_X1 U561 ( .A(n544), .ZN(n541) );
  INV_X1 U562 ( .A(KEYINPUT101), .ZN(n473) );
  XNOR2_X1 U563 ( .A(n751), .B(KEYINPUT24), .ZN(n484) );
  NAND2_X1 U564 ( .A1(n477), .A2(G221), .ZN(n482) );
  XOR2_X1 U565 ( .A(KEYINPUT89), .B(G110), .Z(n479) );
  XNOR2_X1 U566 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U567 ( .A(n480), .B(KEYINPUT23), .Z(n481) );
  XNOR2_X1 U568 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U569 ( .A(n484), .B(n483), .ZN(n637) );
  NAND2_X1 U570 ( .A1(n637), .A2(n485), .ZN(n489) );
  XOR2_X1 U571 ( .A(KEYINPUT90), .B(KEYINPUT25), .Z(n487) );
  NAND2_X1 U572 ( .A1(n636), .A2(G234), .ZN(n486) );
  XNOR2_X1 U573 ( .A(n486), .B(KEYINPUT20), .ZN(n490) );
  XNOR2_X1 U574 ( .A(n487), .B(n412), .ZN(n488) );
  AND2_X1 U575 ( .A1(n490), .A2(G221), .ZN(n492) );
  INV_X1 U576 ( .A(KEYINPUT21), .ZN(n491) );
  XNOR2_X1 U577 ( .A(n492), .B(n491), .ZN(n695) );
  NAND2_X1 U578 ( .A1(G234), .A2(G237), .ZN(n493) );
  XNOR2_X1 U579 ( .A(n493), .B(KEYINPUT14), .ZN(n494) );
  NAND2_X1 U580 ( .A1(G952), .A2(n494), .ZN(n722) );
  OR2_X1 U581 ( .A1(n722), .A2(G953), .ZN(n522) );
  INV_X1 U582 ( .A(n522), .ZN(n497) );
  NAND2_X1 U583 ( .A1(G902), .A2(n494), .ZN(n520) );
  OR2_X1 U584 ( .A1(n430), .A2(n520), .ZN(n495) );
  NOR2_X1 U585 ( .A1(n495), .A2(G900), .ZN(n496) );
  NOR2_X1 U586 ( .A1(n497), .A2(n496), .ZN(n498) );
  NOR2_X1 U587 ( .A1(n695), .A2(n498), .ZN(n588) );
  XNOR2_X1 U588 ( .A(n588), .B(KEYINPUT70), .ZN(n499) );
  NAND2_X1 U589 ( .A1(n514), .A2(n499), .ZN(n605) );
  NAND2_X1 U590 ( .A1(n500), .A2(G210), .ZN(n503) );
  XNOR2_X1 U591 ( .A(G101), .B(KEYINPUT5), .ZN(n501) );
  XNOR2_X1 U592 ( .A(n501), .B(G137), .ZN(n502) );
  XNOR2_X1 U593 ( .A(n503), .B(n502), .ZN(n505) );
  XNOR2_X1 U594 ( .A(n505), .B(n504), .ZN(n506) );
  INV_X1 U595 ( .A(G472), .ZN(n507) );
  INV_X1 U596 ( .A(KEYINPUT6), .ZN(n509) );
  XNOR2_X1 U597 ( .A(n537), .B(n509), .ZN(n551) );
  INV_X1 U598 ( .A(n551), .ZN(n510) );
  NAND2_X1 U599 ( .A1(n362), .A2(n510), .ZN(n613) );
  NOR2_X1 U600 ( .A1(n553), .A2(n613), .ZN(n511) );
  NAND2_X1 U601 ( .A1(n707), .A2(n511), .ZN(n512) );
  XNOR2_X1 U602 ( .A(n512), .B(KEYINPUT43), .ZN(n513) );
  NAND2_X1 U603 ( .A1(n591), .A2(n513), .ZN(n632) );
  XNOR2_X1 U604 ( .A(n632), .B(G140), .ZN(G42) );
  OR2_X1 U605 ( .A1(n514), .A2(n695), .ZN(n692) );
  NOR2_X1 U606 ( .A1(n515), .A2(n692), .ZN(n516) );
  XNOR2_X1 U607 ( .A(n516), .B(KEYINPUT73), .ZN(n533) );
  XNOR2_X1 U608 ( .A(KEYINPUT66), .B(KEYINPUT19), .ZN(n519) );
  INV_X1 U609 ( .A(G898), .ZN(n577) );
  NAND2_X1 U610 ( .A1(G953), .A2(n577), .ZN(n581) );
  OR2_X1 U611 ( .A1(n520), .A2(n581), .ZN(n521) );
  NAND2_X1 U612 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U613 ( .A(n523), .B(KEYINPUT88), .ZN(n524) );
  NAND2_X1 U614 ( .A1(n610), .A2(n524), .ZN(n525) );
  INV_X1 U615 ( .A(n548), .ZN(n534) );
  INV_X1 U616 ( .A(KEYINPUT34), .ZN(n526) );
  INV_X1 U617 ( .A(n545), .ZN(n527) );
  NAND2_X1 U618 ( .A1(n527), .A2(n541), .ZN(n601) );
  XNOR2_X2 U619 ( .A(n528), .B(KEYINPUT35), .ZN(n761) );
  INV_X1 U620 ( .A(n761), .ZN(n529) );
  NAND2_X1 U621 ( .A1(n529), .A2(KEYINPUT44), .ZN(n532) );
  INV_X1 U622 ( .A(KEYINPUT44), .ZN(n530) );
  NAND2_X1 U623 ( .A1(n530), .A2(n566), .ZN(n531) );
  NOR2_X1 U624 ( .A1(n533), .A2(n537), .ZN(n703) );
  NAND2_X1 U625 ( .A1(n703), .A2(n534), .ZN(n536) );
  INV_X1 U626 ( .A(n537), .ZN(n697) );
  NOR2_X1 U627 ( .A1(n697), .A2(n692), .ZN(n539) );
  NAND2_X1 U628 ( .A1(n539), .A2(n538), .ZN(n540) );
  OR2_X1 U629 ( .A1(n548), .A2(n540), .ZN(n668) );
  NAND2_X1 U630 ( .A1(n684), .A2(n668), .ZN(n542) );
  NAND2_X1 U631 ( .A1(n545), .A2(n541), .ZN(n685) );
  XNOR2_X1 U632 ( .A(n685), .B(KEYINPUT98), .ZN(n630) );
  AND2_X1 U633 ( .A1(n630), .A2(n596), .ZN(n600) );
  INV_X1 U634 ( .A(n600), .ZN(n713) );
  NAND2_X1 U635 ( .A1(n542), .A2(n713), .ZN(n543) );
  AND2_X1 U636 ( .A1(n545), .A2(n544), .ZN(n711) );
  INV_X1 U637 ( .A(n695), .ZN(n546) );
  NAND2_X1 U638 ( .A1(n711), .A2(n546), .ZN(n547) );
  XNOR2_X1 U639 ( .A(KEYINPUT71), .B(KEYINPUT22), .ZN(n549) );
  NAND2_X1 U640 ( .A1(n564), .A2(n551), .ZN(n559) );
  INV_X1 U641 ( .A(KEYINPUT82), .ZN(n552) );
  XNOR2_X1 U642 ( .A(n559), .B(n552), .ZN(n555) );
  INV_X1 U643 ( .A(n553), .ZN(n691) );
  INV_X1 U644 ( .A(n514), .ZN(n592) );
  AND2_X1 U645 ( .A1(n691), .A2(n592), .ZN(n554) );
  AND2_X1 U646 ( .A1(n555), .A2(n554), .ZN(n666) );
  INV_X1 U647 ( .A(n666), .ZN(n556) );
  NAND2_X1 U648 ( .A1(n364), .A2(n556), .ZN(n557) );
  NOR2_X1 U649 ( .A1(n558), .A2(n557), .ZN(n573) );
  INV_X1 U650 ( .A(n559), .ZN(n560) );
  XNOR2_X1 U651 ( .A(n691), .B(KEYINPUT85), .ZN(n617) );
  AND2_X1 U652 ( .A1(n354), .A2(n691), .ZN(n563) );
  AND2_X1 U653 ( .A1(n564), .A2(n563), .ZN(n674) );
  INV_X1 U654 ( .A(n674), .ZN(n565) );
  NAND2_X1 U655 ( .A1(n363), .A2(n567), .ZN(n571) );
  NAND2_X1 U656 ( .A1(n566), .A2(KEYINPUT44), .ZN(n568) );
  NAND2_X1 U657 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U658 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U659 ( .A1(n573), .A2(n572), .ZN(n574) );
  AND2_X1 U660 ( .A1(n635), .A2(n430), .ZN(n579) );
  NAND2_X1 U661 ( .A1(G953), .A2(G224), .ZN(n575) );
  XOR2_X1 U662 ( .A(KEYINPUT61), .B(n575), .Z(n576) );
  NOR2_X1 U663 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U664 ( .A1(n579), .A2(n578), .ZN(n584) );
  INV_X1 U665 ( .A(n580), .ZN(n582) );
  NAND2_X1 U666 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U667 ( .A(n584), .B(n583), .ZN(G69) );
  INV_X1 U668 ( .A(KEYINPUT30), .ZN(n586) );
  XNOR2_X1 U669 ( .A(n587), .B(n586), .ZN(n590) );
  AND2_X1 U670 ( .A1(n538), .A2(n588), .ZN(n589) );
  AND2_X1 U671 ( .A1(n592), .A2(n708), .ZN(n593) );
  INV_X1 U672 ( .A(KEYINPUT39), .ZN(n594) );
  XNOR2_X1 U673 ( .A(n595), .B(n594), .ZN(n631) );
  INV_X1 U674 ( .A(n596), .ZN(n597) );
  INV_X1 U675 ( .A(KEYINPUT40), .ZN(n598) );
  XOR2_X1 U676 ( .A(G131), .B(n624), .Z(G33) );
  XNOR2_X1 U677 ( .A(n599), .B(G119), .ZN(G21) );
  NAND2_X1 U678 ( .A1(KEYINPUT47), .A2(n600), .ZN(n604) );
  OR2_X1 U679 ( .A1(n601), .A2(n514), .ZN(n602) );
  NOR2_X1 U680 ( .A1(n602), .A2(n591), .ZN(n603) );
  INV_X1 U681 ( .A(KEYINPUT28), .ZN(n606) );
  XNOR2_X1 U682 ( .A(n607), .B(n606), .ZN(n609) );
  XNOR2_X1 U683 ( .A(n538), .B(KEYINPUT102), .ZN(n608) );
  AND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n622) );
  INV_X1 U685 ( .A(KEYINPUT47), .ZN(n611) );
  XNOR2_X1 U686 ( .A(n612), .B(KEYINPUT72), .ZN(n620) );
  XNOR2_X1 U687 ( .A(KEYINPUT105), .B(KEYINPUT36), .ZN(n614) );
  XNOR2_X1 U688 ( .A(n614), .B(KEYINPUT83), .ZN(n615) );
  XNOR2_X1 U689 ( .A(n616), .B(n615), .ZN(n618) );
  NAND2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U691 ( .A(n619), .B(KEYINPUT106), .ZN(n762) );
  AND2_X1 U692 ( .A1(n620), .A2(n762), .ZN(n627) );
  NAND2_X1 U693 ( .A1(n708), .A2(n707), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n623), .B(KEYINPUT42), .ZN(n764) );
  XNOR2_X1 U695 ( .A(n625), .B(KEYINPUT46), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n627), .A2(n626), .ZN(n629) );
  INV_X1 U697 ( .A(KEYINPUT48), .ZN(n628) );
  XNOR2_X1 U698 ( .A(n629), .B(n628), .ZN(n634) );
  OR2_X1 U699 ( .A1(n631), .A2(n630), .ZN(n687) );
  AND2_X1 U700 ( .A1(n687), .A2(n632), .ZN(n633) );
  AND2_X2 U701 ( .A1(n634), .A2(n633), .ZN(n754) );
  NAND2_X1 U702 ( .A1(n746), .A2(G217), .ZN(n639) );
  XNOR2_X1 U703 ( .A(n637), .B(KEYINPUT124), .ZN(n638) );
  XNOR2_X1 U704 ( .A(n639), .B(n638), .ZN(n641) );
  NOR2_X1 U705 ( .A1(n430), .A2(G952), .ZN(n640) );
  NAND2_X1 U706 ( .A1(n641), .A2(n745), .ZN(n642) );
  XNOR2_X1 U707 ( .A(n642), .B(KEYINPUT125), .ZN(G66) );
  NAND2_X1 U708 ( .A1(n746), .A2(G475), .ZN(n647) );
  XNOR2_X1 U709 ( .A(KEYINPUT86), .B(KEYINPUT122), .ZN(n643) );
  XOR2_X1 U710 ( .A(n643), .B(KEYINPUT59), .Z(n644) );
  XNOR2_X1 U711 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U712 ( .A(n647), .B(n646), .ZN(n648) );
  NAND2_X1 U713 ( .A1(n648), .A2(n745), .ZN(n651) );
  XNOR2_X1 U714 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n649) );
  XOR2_X1 U715 ( .A(n649), .B(KEYINPUT67), .Z(n650) );
  XNOR2_X1 U716 ( .A(n651), .B(n650), .ZN(G60) );
  NAND2_X1 U717 ( .A1(n746), .A2(G210), .ZN(n657) );
  XNOR2_X1 U718 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n653) );
  XNOR2_X1 U719 ( .A(KEYINPUT55), .B(KEYINPUT84), .ZN(n652) );
  XNOR2_X1 U720 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U721 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U722 ( .A(n657), .B(n656), .ZN(n658) );
  NAND2_X1 U723 ( .A1(n658), .A2(n745), .ZN(n660) );
  XNOR2_X1 U724 ( .A(KEYINPUT81), .B(KEYINPUT56), .ZN(n659) );
  XNOR2_X1 U725 ( .A(n660), .B(n659), .ZN(G51) );
  NAND2_X1 U726 ( .A1(n746), .A2(G472), .ZN(n663) );
  XOR2_X1 U727 ( .A(KEYINPUT62), .B(n661), .Z(n662) );
  XNOR2_X1 U728 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U729 ( .A1(n664), .A2(n745), .ZN(n665) );
  XNOR2_X1 U730 ( .A(n665), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U731 ( .A(G101), .B(n666), .Z(G3) );
  NOR2_X1 U732 ( .A1(n680), .A2(n668), .ZN(n667) );
  XOR2_X1 U733 ( .A(G104), .B(n667), .Z(G6) );
  NOR2_X1 U734 ( .A1(n685), .A2(n668), .ZN(n673) );
  XOR2_X1 U735 ( .A(KEYINPUT108), .B(KEYINPUT27), .Z(n670) );
  XNOR2_X1 U736 ( .A(G107), .B(KEYINPUT26), .ZN(n669) );
  XNOR2_X1 U737 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U738 ( .A(KEYINPUT107), .B(n671), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n673), .B(n672), .ZN(G9) );
  XOR2_X1 U740 ( .A(G110), .B(n674), .Z(G12) );
  XOR2_X1 U741 ( .A(G128), .B(KEYINPUT29), .Z(n676) );
  OR2_X1 U742 ( .A1(n678), .A2(n685), .ZN(n675) );
  XNOR2_X1 U743 ( .A(n676), .B(n675), .ZN(G30) );
  XNOR2_X1 U744 ( .A(G143), .B(n677), .ZN(G45) );
  OR2_X1 U745 ( .A1(n678), .A2(n680), .ZN(n679) );
  XNOR2_X1 U746 ( .A(n679), .B(G146), .ZN(G48) );
  NOR2_X1 U747 ( .A1(n680), .A2(n684), .ZN(n682) );
  XNOR2_X1 U748 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n681) );
  XNOR2_X1 U749 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U750 ( .A(G113), .B(n683), .ZN(G15) );
  NOR2_X1 U751 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U752 ( .A(G116), .B(n686), .Z(G18) );
  XOR2_X1 U753 ( .A(G134), .B(n687), .Z(n688) );
  XNOR2_X1 U754 ( .A(n688), .B(KEYINPUT111), .ZN(G36) );
  XOR2_X1 U755 ( .A(KEYINPUT117), .B(KEYINPUT53), .Z(n689) );
  XNOR2_X1 U756 ( .A(KEYINPUT116), .B(n689), .ZN(n736) );
  NOR2_X1 U757 ( .A1(n690), .A2(KEYINPUT2), .ZN(n734) );
  NAND2_X1 U758 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U759 ( .A(n693), .B(KEYINPUT113), .ZN(n694) );
  XNOR2_X1 U760 ( .A(KEYINPUT50), .B(n694), .ZN(n701) );
  AND2_X1 U761 ( .A1(n514), .A2(n695), .ZN(n696) );
  XOR2_X1 U762 ( .A(KEYINPUT49), .B(n696), .Z(n698) );
  NOR2_X1 U763 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U764 ( .A(KEYINPUT112), .B(n699), .Z(n700) );
  NOR2_X1 U765 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U767 ( .A(n704), .B(KEYINPUT51), .ZN(n705) );
  NAND2_X1 U768 ( .A1(n705), .A2(n723), .ZN(n719) );
  NOR2_X1 U769 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U770 ( .A(KEYINPUT114), .B(n709), .Z(n710) );
  NAND2_X1 U771 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U772 ( .A(KEYINPUT115), .B(n712), .Z(n716) );
  NAND2_X1 U773 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U774 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U775 ( .A1(n724), .A2(n717), .ZN(n718) );
  NAND2_X1 U776 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U777 ( .A(KEYINPUT52), .B(n720), .Z(n721) );
  NOR2_X1 U778 ( .A1(n722), .A2(n721), .ZN(n727) );
  NAND2_X1 U779 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U780 ( .A1(n430), .A2(n725), .ZN(n726) );
  NOR2_X1 U781 ( .A1(n727), .A2(n726), .ZN(n732) );
  INV_X1 U782 ( .A(KEYINPUT2), .ZN(n729) );
  INV_X1 U783 ( .A(KEYINPUT78), .ZN(n728) );
  NOR2_X1 U784 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U785 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U786 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U787 ( .A(n736), .B(n735), .ZN(G75) );
  NAND2_X1 U788 ( .A1(n746), .A2(G469), .ZN(n742) );
  XOR2_X1 U789 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n739) );
  XNOR2_X1 U790 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n738) );
  XNOR2_X1 U791 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U792 ( .A(n742), .B(n741), .ZN(n743) );
  NAND2_X1 U793 ( .A1(n743), .A2(n745), .ZN(n744) );
  XNOR2_X1 U794 ( .A(n744), .B(KEYINPUT121), .ZN(G54) );
  INV_X1 U795 ( .A(n745), .ZN(n750) );
  NAND2_X1 U796 ( .A1(n746), .A2(G478), .ZN(n747) );
  XOR2_X1 U797 ( .A(n748), .B(n747), .Z(n749) );
  NOR2_X1 U798 ( .A1(n750), .A2(n749), .ZN(G63) );
  XNOR2_X1 U799 ( .A(n751), .B(KEYINPUT126), .ZN(n752) );
  XNOR2_X1 U800 ( .A(n753), .B(n752), .ZN(n756) );
  XNOR2_X1 U801 ( .A(n754), .B(n756), .ZN(n755) );
  NAND2_X1 U802 ( .A1(n755), .A2(n430), .ZN(n760) );
  XOR2_X1 U803 ( .A(G227), .B(n756), .Z(n757) );
  NAND2_X1 U804 ( .A1(n757), .A2(G900), .ZN(n758) );
  NAND2_X1 U805 ( .A1(G953), .A2(n758), .ZN(n759) );
  NAND2_X1 U806 ( .A1(n760), .A2(n759), .ZN(G72) );
  XOR2_X1 U807 ( .A(n761), .B(G122), .Z(G24) );
  XOR2_X1 U808 ( .A(G125), .B(n762), .Z(n763) );
  XNOR2_X1 U809 ( .A(KEYINPUT37), .B(n763), .ZN(G27) );
  XOR2_X1 U810 ( .A(G137), .B(n764), .Z(G39) );
endmodule

