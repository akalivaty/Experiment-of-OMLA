//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1221, new_n1222, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n209));
  XNOR2_X1  g0009(.A(new_n208), .B(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G77), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  AND3_X1   g0024(.A1(KEYINPUT66), .A2(G1), .A3(G13), .ZN(new_n225));
  AOI21_X1  g0025(.A(KEYINPUT66), .B1(G1), .B2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n202), .A2(KEYINPUT67), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n202), .A2(KEYINPUT67), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n231), .A2(G50), .A3(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n210), .B(new_n224), .C1(new_n230), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n219), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  INV_X1    g0044(.A(G50), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n218), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n256), .A3(G274), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n227), .A2(new_n255), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT3), .B(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G222), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G223), .A2(G1698), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI211_X1 g0067(.A(new_n259), .B(new_n264), .C1(new_n212), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n254), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n256), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI211_X1 g0071(.A(new_n258), .B(new_n268), .C1(G226), .C2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G169), .ZN(new_n273));
  INV_X1    g0073(.A(G179), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(new_n272), .ZN(new_n275));
  INV_X1    g0075(.A(G13), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n276), .A2(new_n229), .A3(G1), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G50), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  OAI22_X1  g0080(.A1(new_n225), .A2(new_n226), .B1(new_n280), .B2(new_n206), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n282), .B1(G1), .B2(new_n229), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n279), .B1(new_n284), .B2(G50), .ZN(new_n285));
  NOR2_X1   g0085(.A1(KEYINPUT8), .A2(G58), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT68), .B(G58), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(KEYINPUT8), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n229), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n288), .A2(new_n290), .B1(G150), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT69), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n203), .A2(G20), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT70), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n292), .A2(new_n293), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n285), .B1(new_n298), .B2(new_n282), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n275), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n272), .A2(G190), .ZN(new_n301));
  INV_X1    g0101(.A(G200), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(new_n272), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n299), .A2(KEYINPUT9), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT9), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n307), .B(new_n285), .C1(new_n298), .C2(new_n282), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n304), .A2(new_n305), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n305), .B1(new_n304), .B2(new_n309), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n300), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT13), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n257), .B1(new_n270), .B2(new_n221), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G97), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n280), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n267), .A2(new_n261), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(G232), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n261), .A2(G226), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT71), .B1(new_n267), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT71), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n260), .A2(new_n322), .A3(G226), .A4(new_n261), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n313), .B(new_n315), .C1(new_n325), .C2(new_n259), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n259), .B1(new_n319), .B2(new_n324), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT13), .B1(new_n327), .B2(new_n314), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G190), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n220), .A2(G20), .ZN(new_n332));
  INV_X1    g0132(.A(new_n291), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n332), .B1(new_n289), .B2(new_n212), .C1(new_n333), .C2(new_n245), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(KEYINPUT11), .A3(new_n281), .ZN(new_n335));
  INV_X1    g0135(.A(G1), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT12), .A3(G13), .ZN(new_n337));
  OAI221_X1 g0137(.A(new_n335), .B1(KEYINPUT12), .B2(new_n277), .C1(new_n332), .C2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n220), .B1(new_n283), .B2(KEYINPUT12), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT11), .B1(new_n334), .B2(new_n281), .ZN(new_n340));
  OR3_X1    g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n302), .B1(new_n326), .B2(new_n328), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n331), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n326), .A2(G179), .A3(new_n328), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT72), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n326), .A2(KEYINPUT72), .A3(new_n328), .A4(G179), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n329), .A2(KEYINPUT14), .A3(G169), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT14), .B1(new_n329), .B2(G169), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n343), .B1(new_n352), .B2(new_n341), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G238), .A2(G1698), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n260), .B(new_n354), .C1(new_n219), .C2(G1698), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(G107), .B2(new_n260), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n257), .B1(new_n213), .B2(new_n270), .C1(new_n356), .C2(new_n259), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G200), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n330), .B2(new_n357), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(new_n290), .B1(G20), .B2(G77), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT8), .B(G58), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n362), .B1(new_n333), .B2(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(new_n281), .B1(new_n212), .B2(new_n277), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n212), .B2(new_n283), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n359), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n357), .A2(G179), .ZN(new_n368));
  INV_X1    g0168(.A(G169), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n357), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n366), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n353), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n287), .A2(G68), .ZN(new_n373));
  INV_X1    g0173(.A(new_n202), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n375), .A2(G20), .B1(G159), .B2(new_n291), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n260), .A2(new_n377), .A3(G20), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n260), .A2(KEYINPUT73), .ZN(new_n379));
  OR2_X1    g0179(.A1(KEYINPUT3), .A2(G33), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT73), .ZN(new_n381));
  NAND2_X1  g0181(.A1(KEYINPUT3), .A2(G33), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n379), .A2(new_n229), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n378), .B1(new_n384), .B2(new_n377), .ZN(new_n385));
  OAI211_X1 g0185(.A(KEYINPUT16), .B(new_n376), .C1(new_n385), .C2(new_n220), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n202), .B1(new_n287), .B2(G68), .ZN(new_n388));
  INV_X1    g0188(.A(G159), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n388), .A2(new_n229), .B1(new_n389), .B2(new_n333), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n377), .B1(new_n260), .B2(G20), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n220), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n387), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n386), .A2(new_n281), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n288), .A2(new_n277), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n283), .B2(new_n288), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n257), .B1(new_n270), .B2(new_n219), .ZN(new_n400));
  INV_X1    g0200(.A(G226), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G1698), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n402), .B1(G223), .B2(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G87), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n259), .B1(new_n405), .B2(KEYINPUT74), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT74), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n403), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  AOI211_X1 g0208(.A(G179), .B(new_n400), .C1(new_n406), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(KEYINPUT74), .ZN(new_n410));
  INV_X1    g0210(.A(new_n259), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n408), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n400), .ZN(new_n413));
  AOI21_X1  g0213(.A(G169), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n409), .A2(new_n414), .A3(KEYINPUT75), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT75), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n403), .A2(new_n407), .A3(new_n404), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n407), .B1(new_n403), .B2(new_n404), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n417), .A2(new_n418), .A3(new_n259), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n369), .B1(new_n419), .B2(new_n400), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n412), .A2(new_n274), .A3(new_n413), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n416), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n399), .B1(new_n415), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT18), .ZN(new_n424));
  OAI21_X1  g0224(.A(G200), .B1(new_n419), .B2(new_n400), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n400), .B1(new_n406), .B2(new_n408), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G190), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n395), .A2(new_n398), .A3(new_n425), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT17), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n302), .B1(new_n412), .B2(new_n413), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(G190), .B2(new_n426), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT17), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(new_n395), .A4(new_n398), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT75), .B1(new_n409), .B2(new_n414), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n420), .A2(new_n416), .A3(new_n421), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n435), .A2(new_n436), .B1(new_n395), .B2(new_n398), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT18), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n424), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n312), .A2(new_n372), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G116), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n277), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n277), .B1(new_n336), .B2(G33), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n282), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n444), .B1(new_n446), .B2(new_n443), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G283), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n448), .B(new_n229), .C1(G33), .C2(new_n316), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n443), .A2(G20), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n281), .A2(KEYINPUT80), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT80), .B1(new_n281), .B2(new_n450), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT20), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(KEYINPUT20), .B(new_n449), .C1(new_n451), .C2(new_n452), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n447), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n256), .A2(G274), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n253), .A2(G1), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT5), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G41), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  OR2_X1    g0264(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n261), .A2(G257), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G264), .A2(G1698), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n466), .B(new_n467), .C1(new_n265), .C2(new_n266), .ZN(new_n468));
  INV_X1    g0268(.A(G303), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n380), .A2(new_n469), .A3(new_n382), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n468), .A2(new_n227), .A3(new_n470), .A4(new_n255), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n464), .A2(G270), .A3(new_n256), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n465), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G200), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n330), .B2(new_n473), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n458), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT21), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n473), .A2(G169), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n478), .B1(new_n457), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT81), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT81), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n482), .B(new_n478), .C1(new_n457), .C2(new_n479), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n473), .A2(new_n274), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n479), .A2(new_n478), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n458), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n477), .A2(new_n481), .A3(new_n483), .A4(new_n486), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n445), .A2(new_n282), .A3(G107), .ZN(new_n488));
  INV_X1    g0288(.A(G107), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n336), .A2(new_n489), .A3(G13), .A4(G20), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT25), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n492), .B(KEYINPUT84), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n277), .A2(KEYINPUT83), .A3(KEYINPUT25), .A4(new_n489), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT83), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n490), .B2(new_n491), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n488), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT23), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(new_n229), .B2(G107), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n489), .A2(KEYINPUT23), .A3(G20), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n229), .A2(G33), .A3(G116), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT82), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT24), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n229), .B(G87), .C1(new_n265), .C2(new_n266), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT22), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT22), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n260), .A2(new_n511), .A3(new_n229), .A4(G87), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n508), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n506), .A2(KEYINPUT24), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n281), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n510), .A2(new_n512), .ZN(new_n517));
  INV_X1    g0317(.A(new_n508), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n514), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n500), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n459), .A2(new_n464), .ZN(new_n522));
  OAI211_X1 g0322(.A(G250), .B(new_n261), .C1(new_n265), .C2(new_n266), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT85), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n260), .A2(KEYINPUT85), .A3(G250), .A4(new_n261), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G294), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n260), .A2(G257), .A3(G1698), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n525), .A2(new_n526), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n522), .B1(new_n529), .B2(new_n411), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n336), .B(G45), .C1(new_n252), .C2(KEYINPUT5), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n462), .A2(G41), .ZN(new_n532));
  OAI211_X1 g0332(.A(G264), .B(new_n256), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT86), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n464), .A2(KEYINPUT86), .A3(G264), .A4(new_n256), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n530), .A2(G179), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n369), .B1(new_n530), .B2(new_n533), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n521), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI22_X1  g0340(.A1(new_n493), .A2(new_n498), .B1(new_n446), .B2(new_n489), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n282), .B1(new_n519), .B2(new_n514), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n513), .A2(new_n515), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n530), .A2(new_n330), .A3(new_n533), .ZN(new_n545));
  AOI21_X1  g0345(.A(G200), .B1(new_n530), .B2(new_n537), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n260), .A2(G250), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n261), .B1(new_n549), .B2(KEYINPUT4), .ZN(new_n550));
  AND2_X1   g0350(.A1(KEYINPUT4), .A2(G244), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n261), .B(new_n551), .C1(new_n265), .C2(new_n266), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n213), .B1(new_n380), .B2(new_n382), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n448), .B(new_n552), .C1(new_n553), .C2(KEYINPUT4), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n411), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n464), .A2(new_n256), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n522), .B1(new_n556), .B2(G257), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT76), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n302), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n555), .A2(KEYINPUT76), .A3(new_n557), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n555), .A2(G190), .A3(new_n557), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT6), .ZN(new_n564));
  NOR3_X1   g0364(.A1(new_n564), .A2(new_n316), .A3(G107), .ZN(new_n565));
  XNOR2_X1  g0365(.A(G97), .B(G107), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n565), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n567), .A2(new_n229), .B1(new_n212), .B2(new_n333), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n489), .B1(new_n391), .B2(new_n392), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n281), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  MUX2_X1   g0370(.A(new_n278), .B(new_n446), .S(G97), .Z(new_n571));
  AND3_X1   g0371(.A1(new_n563), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n555), .A2(new_n557), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n570), .A2(new_n571), .B1(new_n573), .B2(new_n369), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n555), .A2(new_n557), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n274), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n562), .A2(new_n572), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n260), .A2(new_n229), .A3(G68), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n214), .A2(new_n316), .A3(new_n489), .ZN(new_n579));
  OAI211_X1 g0379(.A(KEYINPUT19), .B(new_n579), .C1(new_n317), .C2(G20), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n289), .A2(new_n316), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n578), .B(new_n580), .C1(KEYINPUT19), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n281), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n360), .A2(new_n277), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n445), .A2(new_n282), .A3(G87), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G274), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n460), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n215), .B1(new_n253), .B2(G1), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n256), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(G244), .B(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT77), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT77), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n260), .A2(new_n594), .A3(G244), .A4(G1698), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G116), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n260), .A2(G238), .A3(new_n261), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n593), .A2(new_n595), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n591), .B1(new_n598), .B2(new_n411), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G190), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n586), .B(new_n600), .C1(new_n302), .C2(new_n599), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n274), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n361), .A2(KEYINPUT78), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT78), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n360), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n583), .B(new_n584), .C1(new_n446), .C2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n602), .B(new_n607), .C1(G169), .C2(new_n599), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT79), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT79), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n601), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n577), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NOR4_X1   g0413(.A1(new_n442), .A2(new_n487), .A3(new_n548), .A4(new_n613), .ZN(G372));
  NAND2_X1  g0414(.A1(new_n574), .A2(new_n576), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n610), .A2(new_n612), .A3(KEYINPUT26), .A4(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n609), .A2(new_n615), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n617), .B1(KEYINPUT26), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n608), .B(KEYINPUT87), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n560), .A2(new_n558), .A3(new_n302), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n571), .A2(new_n570), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n563), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n615), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n547), .A2(new_n608), .A3(new_n601), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n481), .A2(new_n483), .A3(new_n486), .A4(new_n540), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n620), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n619), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n441), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n630), .B(KEYINPUT88), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n310), .A2(new_n311), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n435), .A2(new_n436), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n633), .A2(new_n438), .A3(new_n399), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n438), .B1(new_n633), .B2(new_n399), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n343), .ZN(new_n637));
  INV_X1    g0437(.A(new_n371), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n341), .A2(new_n352), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n434), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n632), .A2(new_n641), .B1(new_n299), .B2(new_n275), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n631), .A2(new_n642), .ZN(G369));
  NAND3_X1  g0443(.A1(new_n481), .A2(new_n483), .A3(new_n486), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n336), .A2(new_n229), .A3(G13), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT27), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n647), .A2(new_n336), .A3(new_n229), .A4(G13), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(G213), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g0449(.A(new_n649), .B(KEYINPUT89), .Z(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT90), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n649), .B(KEYINPUT89), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT90), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n654), .A3(G343), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(new_n457), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n644), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n487), .B2(new_n657), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n656), .A2(new_n544), .ZN(new_n662));
  OAI22_X1  g0462(.A1(new_n548), .A2(new_n662), .B1(new_n540), .B2(new_n656), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n644), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n540), .A2(new_n547), .A3(new_n656), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n540), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n667), .B1(new_n668), .B2(new_n656), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n664), .A2(new_n669), .ZN(G399));
  INV_X1    g0470(.A(KEYINPUT91), .ZN(new_n671));
  INV_X1    g0471(.A(new_n207), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n671), .B1(new_n672), .B2(G41), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n207), .A2(KEYINPUT91), .A3(new_n252), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n579), .A2(G116), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G1), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n233), .B2(new_n675), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  INV_X1    g0479(.A(G330), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n529), .A2(new_n411), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(new_n537), .A3(new_n465), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n473), .A2(new_n274), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n682), .A2(new_n573), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n598), .A2(new_n411), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n590), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT92), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT92), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n599), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n684), .A2(new_n690), .A3(KEYINPUT93), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT93), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n688), .B1(new_n685), .B2(new_n590), .ZN(new_n693));
  AOI211_X1 g0493(.A(KEYINPUT92), .B(new_n591), .C1(new_n598), .C2(new_n411), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n682), .A2(new_n573), .A3(new_n683), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n692), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT30), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n575), .A2(new_n599), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n484), .A2(new_n681), .A3(new_n537), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n484), .A2(new_n681), .A3(new_n537), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n702), .A2(KEYINPUT30), .A3(new_n599), .A4(new_n575), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n691), .A2(new_n697), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n656), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT31), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n656), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n701), .B(new_n703), .C1(new_n695), .C2(new_n696), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n706), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n613), .A2(new_n666), .ZN(new_n711));
  INV_X1    g0511(.A(new_n487), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n680), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n618), .A2(KEYINPUT26), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n610), .A2(new_n612), .A3(new_n616), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(KEYINPUT26), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n628), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(KEYINPUT29), .A3(new_n656), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT95), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n705), .B1(new_n717), .B2(new_n628), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT95), .A3(KEYINPUT29), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT29), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT94), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n629), .B2(new_n656), .ZN(new_n727));
  AOI211_X1 g0527(.A(KEYINPUT94), .B(new_n705), .C1(new_n619), .C2(new_n628), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n714), .B1(new_n724), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n679), .B1(new_n730), .B2(G1), .ZN(G364));
  AOI21_X1  g0531(.A(new_n228), .B1(G20), .B2(new_n369), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G13), .A2(G33), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n247), .A2(G45), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n379), .A2(new_n383), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n672), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n738), .B(new_n740), .C1(G45), .C2(new_n233), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n260), .A2(new_n207), .ZN(new_n742));
  INV_X1    g0542(.A(G355), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n742), .A2(new_n743), .B1(G116), .B2(new_n207), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT96), .Z(new_n745));
  AOI21_X1  g0545(.A(new_n737), .B1(new_n741), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n732), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n229), .A2(G190), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G179), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G159), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT32), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n302), .A2(G179), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G107), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n274), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n748), .ZN(new_n759));
  INV_X1    g0559(.A(new_n287), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n229), .A2(new_n330), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n758), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n757), .B1(new_n212), .B2(new_n759), .C1(new_n760), .C2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G190), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n764), .A2(new_n330), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n766), .A2(new_n220), .B1(new_n768), .B2(new_n245), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n761), .A2(new_n754), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G87), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n229), .B1(new_n749), .B2(G190), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n772), .B(new_n260), .C1(new_n316), .C2(new_n773), .ZN(new_n774));
  OR4_X1    g0574(.A1(new_n753), .A2(new_n763), .A3(new_n769), .A4(new_n774), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n767), .A2(G326), .ZN(new_n776));
  INV_X1    g0576(.A(new_n762), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n260), .B(new_n776), .C1(G322), .C2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n759), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G283), .A2(new_n756), .B1(new_n779), .B2(G311), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G303), .A2(new_n771), .B1(new_n751), .B2(G329), .ZN(new_n781));
  INV_X1    g0581(.A(new_n773), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT33), .B(G317), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n782), .A2(G294), .B1(new_n765), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n778), .A2(new_n780), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n747), .B1(new_n775), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n675), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n276), .A2(G20), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n336), .B1(new_n788), .B2(G45), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n746), .A2(new_n786), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n735), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n659), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n660), .A2(new_n792), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n659), .A2(G330), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(G396));
  NOR2_X1   g0598(.A1(new_n371), .A2(new_n705), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n705), .A2(new_n366), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n367), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n799), .B1(new_n371), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n727), .B2(new_n728), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n629), .A2(new_n656), .A3(new_n802), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n714), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n791), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n804), .A2(new_n714), .A3(new_n805), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n732), .A2(new_n733), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n267), .B1(new_n773), .B2(new_n316), .C1(new_n489), .C2(new_n770), .ZN(new_n812));
  INV_X1    g0612(.A(G283), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n766), .A2(new_n813), .B1(new_n768), .B2(new_n469), .ZN(new_n814));
  INV_X1    g0614(.A(G294), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n762), .A2(new_n815), .B1(new_n759), .B2(new_n443), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n755), .A2(new_n214), .B1(new_n750), .B2(new_n817), .ZN(new_n818));
  NOR4_X1   g0618(.A1(new_n812), .A2(new_n814), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G143), .A2(new_n777), .B1(new_n779), .B2(G159), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  INV_X1    g0621(.A(G150), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n768), .B2(new_n821), .C1(new_n822), .C2(new_n766), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT34), .ZN(new_n824));
  INV_X1    g0624(.A(new_n739), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G68), .A2(new_n756), .B1(new_n751), .B2(G132), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n245), .B2(new_n770), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n825), .B(new_n827), .C1(new_n287), .C2(new_n782), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n819), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n791), .B1(G77), .B2(new_n811), .C1(new_n829), .C2(new_n747), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT97), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n734), .B2(new_n802), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n809), .A2(new_n832), .ZN(G384));
  NOR2_X1   g0633(.A1(new_n788), .A2(new_n336), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n724), .A2(new_n441), .A3(new_n729), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n642), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT100), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n636), .A2(new_n653), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n376), .B1(new_n385), .B2(new_n220), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n387), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n840), .A2(new_n281), .A3(new_n386), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n650), .B1(new_n841), .B2(new_n398), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n440), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n386), .A2(new_n281), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n397), .B1(new_n844), .B2(new_n840), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n428), .B1(new_n845), .B2(new_n650), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n435), .A2(new_n436), .B1(new_n841), .B2(new_n398), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT37), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n650), .B1(new_n395), .B2(new_n398), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n423), .A2(new_n849), .A3(new_n428), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n843), .A2(KEYINPUT38), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT38), .B1(new_n843), .B2(new_n853), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT39), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n843), .A2(KEYINPUT38), .A3(new_n853), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT39), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n423), .A2(new_n428), .A3(new_n851), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n440), .A2(new_n850), .B1(new_n860), .B2(new_n852), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n857), .B(new_n858), .C1(new_n861), .C2(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n351), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n864), .A2(new_n349), .B1(new_n346), .B2(new_n347), .ZN(new_n865));
  INV_X1    g0665(.A(new_n341), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n865), .A2(new_n866), .A3(new_n705), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n838), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n866), .A2(new_n656), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT99), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT99), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n352), .A2(new_n872), .A3(new_n869), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n871), .A2(new_n873), .B1(new_n353), .B2(new_n870), .ZN(new_n874));
  INV_X1    g0674(.A(new_n799), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n874), .B1(new_n805), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  INV_X1    g0677(.A(new_n842), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n636), .B2(new_n434), .ZN(new_n879));
  AND4_X1   g0679(.A1(new_n395), .A2(new_n398), .A3(new_n425), .A4(new_n427), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n842), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n841), .A2(new_n398), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n633), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n849), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NOR4_X1   g0684(.A1(new_n437), .A2(new_n880), .A3(KEYINPUT37), .A4(new_n850), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n877), .B1(new_n879), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n857), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n876), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n868), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n837), .B(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n874), .A2(new_n803), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n540), .A2(new_n547), .A3(new_n656), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n893), .A2(new_n612), .A3(new_n610), .A4(new_n577), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n706), .A2(KEYINPUT101), .B1(new_n894), .B2(new_n487), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n704), .A2(new_n708), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT102), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT102), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n704), .A2(new_n899), .A3(new_n708), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n898), .A2(new_n900), .B1(new_n706), .B2(KEYINPUT101), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT103), .B1(new_n896), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n704), .A2(new_n705), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(KEYINPUT101), .A3(new_n707), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n899), .B1(new_n704), .B2(new_n708), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n704), .A2(new_n899), .A3(new_n708), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT103), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n907), .A2(new_n895), .A3(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n888), .B(new_n892), .C1(new_n902), .C2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n637), .B(new_n870), .C1(new_n865), .C2(new_n866), .ZN(new_n912));
  INV_X1    g0712(.A(new_n873), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n872), .B1(new_n352), .B2(new_n869), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n802), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n896), .A2(KEYINPUT103), .A3(new_n901), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n908), .B1(new_n907), .B2(new_n895), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n857), .B1(new_n861), .B2(KEYINPUT38), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n920), .A2(KEYINPUT40), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n910), .A2(new_n911), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n442), .B1(new_n918), .B2(new_n917), .ZN(new_n923));
  OAI21_X1  g0723(.A(G330), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT104), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n924), .A2(new_n925), .B1(new_n922), .B2(new_n923), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n925), .B2(new_n924), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n834), .B1(new_n891), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n891), .B2(new_n927), .ZN(new_n929));
  INV_X1    g0729(.A(new_n567), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n930), .A2(KEYINPUT35), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(KEYINPUT35), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n931), .A2(G116), .A3(new_n230), .A4(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT36), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n201), .A2(G68), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT98), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n212), .B1(new_n287), .B2(G68), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n234), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n276), .A2(G1), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n929), .B(new_n934), .C1(new_n938), .C2(new_n939), .ZN(G367));
  OAI21_X1  g0740(.A(new_n577), .B1(new_n622), .B2(new_n656), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n616), .A2(new_n705), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n667), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT106), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT42), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n615), .B1(new_n941), .B2(new_n540), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n945), .A2(KEYINPUT42), .B1(new_n656), .B2(new_n947), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n608), .B(new_n601), .C1(new_n656), .C2(new_n586), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT105), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n586), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n620), .A2(new_n952), .A3(new_n705), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n949), .A2(new_n950), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n946), .A2(new_n948), .B1(KEYINPUT43), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n956), .B(new_n957), .Z(new_n958));
  INV_X1    g0758(.A(new_n943), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n664), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n958), .A2(new_n961), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n675), .B(KEYINPUT41), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n669), .A2(new_n943), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT107), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT45), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n967), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n669), .A2(new_n943), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT44), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n664), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n665), .A2(new_n705), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n975), .A2(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n661), .B(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n730), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n968), .A2(new_n664), .A3(new_n969), .A4(new_n971), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n974), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n964), .B1(new_n981), .B2(new_n730), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n962), .B(new_n963), .C1(new_n982), .C2(new_n790), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n736), .B1(new_n207), .B2(new_n360), .ZN(new_n984));
  INV_X1    g0784(.A(new_n740), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(new_n242), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n791), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n762), .A2(new_n469), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n316), .A2(new_n755), .B1(new_n759), .B2(new_n813), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(G317), .C2(new_n751), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT46), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n770), .B2(new_n443), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT108), .Z(new_n993));
  OAI22_X1  g0793(.A1(new_n766), .A2(new_n815), .B1(new_n773), .B2(new_n489), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n770), .A2(new_n991), .A3(new_n443), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n739), .B1(G311), .B2(new_n767), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n990), .A2(new_n993), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n760), .A2(new_n770), .B1(new_n750), .B2(new_n821), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n762), .A2(new_n822), .B1(new_n755), .B2(new_n212), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G143), .A2(new_n767), .B1(new_n765), .B2(G159), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n773), .A2(new_n220), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n201), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n267), .B1(new_n1005), .B2(new_n779), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n998), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n987), .B1(new_n1010), .B2(new_n732), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n955), .B2(new_n794), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n983), .A2(new_n1012), .ZN(G387));
  OR2_X1    g0813(.A1(new_n663), .A2(new_n794), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n742), .A2(new_n676), .B1(G107), .B2(new_n207), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n239), .A2(G45), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n676), .ZN(new_n1017));
  AOI211_X1 g0817(.A(G45), .B(new_n1017), .C1(G68), .C2(G77), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n363), .A2(G50), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT50), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n985), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1015), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n791), .B1(new_n1022), .B2(new_n737), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n771), .A2(G77), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n220), .B2(new_n759), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n606), .A2(new_n773), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(G150), .C2(new_n751), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n762), .A2(new_n245), .B1(new_n755), .B2(new_n316), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1028), .B(new_n825), .C1(G159), .C2(new_n767), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n288), .A2(new_n765), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G317), .A2(new_n777), .B1(new_n779), .B2(G303), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1032), .A2(KEYINPUT110), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(KEYINPUT110), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G311), .A2(new_n765), .B1(new_n767), .B2(G322), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT48), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n770), .A2(new_n815), .B1(new_n773), .B2(new_n813), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(KEYINPUT49), .A3(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G116), .A2(new_n756), .B1(new_n751), .B2(G326), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1041), .A2(new_n825), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(KEYINPUT49), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1031), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1023), .B1(new_n1045), .B2(new_n732), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n977), .A2(new_n790), .B1(new_n1014), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n978), .A2(new_n787), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n730), .A2(new_n977), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(G393));
  INV_X1    g0850(.A(KEYINPUT111), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n974), .A2(new_n1051), .A3(new_n980), .ZN(new_n1052));
  OR3_X1    g0852(.A1(new_n972), .A2(new_n1051), .A3(new_n973), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n787), .B(new_n981), .C1(new_n1054), .C2(new_n979), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n777), .A2(G159), .B1(G150), .B2(new_n767), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT112), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT51), .Z(new_n1058));
  AOI22_X1  g0858(.A1(G87), .A2(new_n756), .B1(new_n751), .B2(G143), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n220), .B2(new_n770), .C1(new_n363), .C2(new_n759), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n766), .A2(new_n201), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n782), .A2(G77), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n739), .A2(new_n1062), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n766), .A2(new_n469), .B1(new_n773), .B2(new_n443), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1065), .A2(KEYINPUT113), .B1(G294), .B2(new_n779), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(KEYINPUT113), .B2(new_n1065), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT114), .Z(new_n1068));
  AOI22_X1  g0868(.A1(new_n777), .A2(G311), .B1(G317), .B2(new_n767), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT52), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G283), .A2(new_n771), .B1(new_n751), .B2(G322), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1071), .A2(new_n267), .A3(new_n757), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1068), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n732), .B1(new_n1064), .B2(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n250), .A2(new_n740), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n736), .B1(new_n316), .B2(new_n207), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1074), .B(new_n791), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n959), .B2(new_n735), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n1054), .B2(new_n790), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1055), .A2(new_n1079), .ZN(G390));
  OAI21_X1  g0880(.A(new_n791), .B1(new_n811), .B2(new_n288), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G116), .A2(new_n777), .B1(new_n751), .B2(G294), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n220), .B2(new_n755), .C1(new_n316), .C2(new_n759), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G107), .A2(new_n765), .B1(new_n767), .B2(G283), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n772), .A2(new_n1084), .A3(new_n1062), .A4(new_n267), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n782), .A2(G159), .B1(G137), .B2(new_n765), .ZN(new_n1086));
  INV_X1    g0886(.A(G128), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n770), .A2(new_n822), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1086), .B1(new_n1087), .B2(new_n768), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(KEYINPUT54), .B(G143), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n777), .A2(G132), .B1(new_n779), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1005), .A2(new_n756), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n267), .B1(new_n751), .B2(G125), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1083), .A2(new_n1085), .B1(new_n1090), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1081), .B1(new_n1098), .B2(new_n732), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n863), .B2(new_n734), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n867), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n801), .A2(new_n371), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n799), .B1(new_n722), .B2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1101), .B(new_n920), .C1(new_n1103), .C2(new_n874), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n876), .A2(new_n867), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n863), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n802), .A2(G330), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n874), .B(new_n1107), .C1(new_n917), .C2(new_n918), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n714), .A2(new_n802), .A3(new_n915), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1104), .B(new_n1110), .C1(new_n1105), .C2(new_n863), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1100), .B1(new_n1112), .B2(new_n789), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT116), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n441), .B(G330), .C1(new_n902), .C2(new_n909), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n835), .A2(new_n642), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1107), .B1(new_n917), .B2(new_n918), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1110), .B(new_n1103), .C1(new_n1118), .C2(new_n915), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n915), .B1(new_n714), .B2(new_n802), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1118), .B2(new_n915), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n805), .A2(new_n875), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1119), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n1112), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1117), .A2(new_n1124), .A3(new_n1109), .A4(new_n1111), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n787), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1115), .A2(new_n1128), .A3(new_n1129), .ZN(G378));
  NAND2_X1  g0930(.A1(new_n910), .A2(new_n911), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n919), .A2(new_n921), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(G330), .A3(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n312), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n312), .A2(new_n1134), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1136), .A2(new_n299), .A3(new_n653), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n299), .A2(new_n653), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1137), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1139), .B1(new_n1140), .B2(new_n1135), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1133), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n890), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n922), .A2(G330), .A3(new_n1142), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1145), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n790), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1143), .A2(new_n733), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n791), .B1(new_n811), .B2(new_n1005), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1004), .B1(new_n766), .B2(new_n316), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n739), .A2(G41), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n756), .A2(new_n287), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G107), .A2(new_n777), .B1(new_n751), .B2(G283), .ZN(new_n1155));
  AND4_X1   g0955(.A1(new_n1024), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n606), .B2(new_n759), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1152), .B(new_n1157), .C1(G116), .C2(new_n767), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1158), .A2(KEYINPUT58), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n767), .A2(G125), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n822), .B2(new_n773), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G128), .A2(new_n777), .B1(new_n771), .B2(new_n1092), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n821), .B2(new_n759), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1161), .B(new_n1163), .C1(G132), .C2(new_n765), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1165), .A2(KEYINPUT59), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(KEYINPUT59), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n755), .A2(new_n389), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n280), .A2(new_n252), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT117), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT118), .B(G124), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1168), .B(new_n1170), .C1(new_n751), .C2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1166), .A2(new_n1167), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1158), .A2(KEYINPUT58), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n245), .B(new_n1170), .C1(new_n739), .C2(G41), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1159), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1151), .B1(new_n1176), .B2(new_n732), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1150), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1149), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1124), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1117), .B1(new_n1112), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT57), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n675), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1133), .A2(new_n1143), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1142), .B1(new_n922), .B2(G330), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n890), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1187), .A2(new_n1188), .B1(new_n1117), .B2(new_n1127), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT57), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1179), .B1(new_n1184), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(G375));
  AOI21_X1  g0992(.A(new_n1026), .B1(G283), .B2(new_n777), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT119), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n267), .B1(new_n755), .B2(new_n212), .C1(new_n768), .C2(new_n815), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G116), .B2(new_n765), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G97), .A2(new_n771), .B1(new_n751), .B2(G303), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(new_n489), .C2(new_n759), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1194), .A2(new_n1198), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n770), .A2(new_n389), .B1(new_n750), .B2(new_n1087), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT120), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n782), .A2(G50), .B1(G132), .B2(new_n767), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1202), .B(new_n739), .C1(new_n766), .C2(new_n1091), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n762), .A2(new_n821), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1154), .B1(new_n822), .B2(new_n759), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1201), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n732), .B1(new_n1199), .B2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1207), .B(new_n791), .C1(G68), .C2(new_n811), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n874), .B2(new_n733), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1124), .B2(new_n790), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n964), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1125), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1210), .B1(new_n1212), .B2(new_n1213), .ZN(G381));
  NOR2_X1   g1014(.A1(G387), .A2(G390), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1128), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1216), .A2(new_n1113), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1191), .A3(new_n1217), .A4(new_n1218), .ZN(G407));
  NAND2_X1  g1019(.A1(new_n651), .A2(G213), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1191), .A2(new_n1217), .A3(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(G407), .A2(G213), .A3(new_n1222), .ZN(G409));
  INV_X1    g1023(.A(KEYINPUT126), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT60), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1117), .B2(new_n1124), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n675), .B1(new_n1117), .B2(new_n1124), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n835), .A2(new_n642), .A3(new_n1116), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1122), .B1(new_n1108), .B2(new_n1120), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1228), .A2(new_n1229), .A3(KEYINPUT60), .A4(new_n1119), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1226), .A2(new_n1227), .A3(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1231), .A2(G384), .A3(new_n1210), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1210), .ZN(new_n1233));
  INV_X1    g1033(.A(G384), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1232), .B1(new_n1235), .B2(KEYINPUT122), .ZN(new_n1236));
  INV_X1    g1036(.A(G2897), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1220), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(G384), .B1(new_n1231), .B2(new_n1210), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT122), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1236), .A2(KEYINPUT123), .A3(new_n1238), .A4(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1238), .A2(KEYINPUT123), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1238), .A2(KEYINPUT123), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1241), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1231), .A2(G384), .A3(new_n1210), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1243), .B(new_n1244), .C1(new_n1245), .C2(new_n1247), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1242), .A2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1181), .B(new_n1211), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT121), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1252), .A2(new_n790), .B1(new_n1150), .B2(new_n1177), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT121), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1252), .A2(new_n1254), .A3(new_n1211), .A4(new_n1181), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1251), .A2(new_n1253), .A3(new_n1255), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1191), .A2(G378), .B1(new_n1256), .B2(new_n1217), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT125), .B1(new_n1257), .B2(new_n1221), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1256), .A2(new_n1217), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n787), .B1(new_n1189), .B2(KEYINPUT57), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G378), .B(new_n1253), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT125), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1220), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1249), .B1(new_n1258), .B2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1224), .B1(new_n1266), .B2(KEYINPUT61), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1242), .A2(new_n1248), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1264), .B1(new_n1263), .B2(new_n1220), .ZN(new_n1269));
  AOI211_X1 g1069(.A(KEYINPUT125), .B(new_n1221), .C1(new_n1259), .C2(new_n1262), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1268), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT61), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(KEYINPUT126), .A3(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1258), .A2(KEYINPUT62), .A3(new_n1265), .A4(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1263), .A2(new_n1220), .A3(new_n1274), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1267), .A2(new_n1273), .A3(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1215), .ZN(new_n1281));
  XOR2_X1   g1081(.A(G393), .B(G396), .Z(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n983), .A2(new_n1012), .B1(new_n1055), .B2(new_n1079), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1281), .A2(new_n1283), .A3(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1282), .B1(new_n1215), .B2(new_n1284), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1280), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1276), .A2(new_n1290), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1288), .A2(new_n1291), .A3(KEYINPUT61), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1258), .A2(KEYINPUT63), .A3(new_n1265), .A4(new_n1274), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1249), .B1(new_n1220), .B2(new_n1263), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT124), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1292), .B(new_n1293), .C1(new_n1296), .C2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1289), .A2(new_n1298), .ZN(G405));
  INV_X1    g1099(.A(new_n1217), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1262), .B1(new_n1191), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1288), .A2(KEYINPUT127), .A3(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT127), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1286), .B(new_n1287), .C1(new_n1304), .C2(new_n1301), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1274), .B1(new_n1301), .B2(new_n1304), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1306), .B(new_n1307), .ZN(G402));
endmodule


