//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1307, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n205), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT66), .ZN(new_n214));
  AND2_X1   g0014(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  NOR3_X1   g0017(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT65), .Z(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(G20), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n205), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT0), .ZN(new_n226));
  AND4_X1   g0026(.A1(new_n214), .A2(new_n222), .A3(new_n223), .A4(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(KEYINPUT16), .ZN(new_n243));
  INV_X1    g0043(.A(G68), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT7), .ZN(new_n245));
  OR2_X1    g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n245), .B1(new_n248), .B2(G20), .ZN(new_n249));
  AND2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G20), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n244), .B1(new_n249), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G58), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(new_n244), .ZN(new_n257));
  OAI21_X1  g0057(.A(G20), .B1(new_n257), .B2(new_n201), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G159), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n243), .B1(new_n255), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT7), .B1(new_n252), .B2(new_n253), .ZN(new_n263));
  NOR4_X1   g0063(.A1(new_n250), .A2(new_n251), .A3(new_n245), .A4(G20), .ZN(new_n264));
  OAI21_X1  g0064(.A(G68), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n265), .A2(KEYINPUT16), .A3(new_n260), .A4(new_n258), .ZN(new_n266));
  NAND3_X1  g0066(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT68), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n267), .A2(new_n268), .A3(new_n220), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n268), .B1(new_n267), .B2(new_n220), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n262), .A2(new_n266), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n221), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g0074(.A(G226), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT77), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT77), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n248), .A2(new_n277), .A3(G226), .A4(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G87), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT78), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  OAI211_X1 g0083(.A(G223), .B(new_n283), .C1(new_n250), .C2(new_n251), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n274), .B1(new_n279), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n273), .A2(KEYINPUT67), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT67), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(G33), .A3(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(new_n290), .A3(new_n221), .ZN(new_n291));
  INV_X1    g0091(.A(G41), .ZN(new_n292));
  INV_X1    g0092(.A(G45), .ZN(new_n293));
  AOI21_X1  g0093(.A(G1), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(G274), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n294), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n291), .A2(G232), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(G200), .B1(new_n287), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G13), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(G1), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G20), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT69), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(new_n269), .B2(new_n270), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n267), .A2(new_n220), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT68), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n267), .A2(new_n268), .A3(new_n220), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(KEYINPUT69), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n303), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT8), .B(G58), .ZN(new_n311));
  INV_X1    g0111(.A(G1), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(G20), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n310), .A2(new_n313), .B1(new_n311), .B2(new_n303), .ZN(new_n314));
  INV_X1    g0114(.A(new_n298), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n285), .B1(new_n278), .B2(new_n276), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n315), .B(G190), .C1(new_n316), .C2(new_n274), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n272), .A2(new_n299), .A3(new_n314), .A4(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT17), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT18), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n272), .A2(new_n314), .ZN(new_n322));
  OAI21_X1  g0122(.A(G169), .B1(new_n287), .B2(new_n298), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n315), .B(G179), .C1(new_n316), .C2(new_n274), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n321), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n322), .A2(new_n325), .A3(new_n321), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n318), .A2(new_n319), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n320), .A2(new_n327), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n271), .A2(new_n303), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n312), .A2(G20), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(G77), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT73), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n334), .B(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n311), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n337), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT15), .B(G87), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT72), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n253), .A2(G33), .ZN(new_n341));
  OR3_X1    g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n340), .B1(new_n339), .B2(new_n341), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n338), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G77), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n344), .A2(new_n271), .B1(new_n345), .B2(new_n303), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n336), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G238), .A2(G1698), .ZN(new_n348));
  INV_X1    g0148(.A(G232), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(G1698), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n248), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G107), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(new_n248), .ZN(new_n353));
  OR2_X1    g0153(.A1(new_n353), .A2(KEYINPUT71), .ZN(new_n354));
  INV_X1    g0154(.A(new_n274), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(KEYINPUT71), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n288), .A2(new_n290), .A3(new_n221), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n294), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G244), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n360), .A2(new_n295), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G169), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G179), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n357), .A2(new_n365), .A3(new_n361), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n347), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n347), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n362), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n357), .B2(new_n361), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n367), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n305), .A2(new_n309), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n259), .A2(G50), .B1(G20), .B2(new_n244), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n345), .B2(new_n341), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(KEYINPUT11), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n305), .A2(new_n309), .A3(new_n378), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT11), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n244), .B1(new_n312), .B2(G20), .ZN(new_n383));
  OR3_X1    g0183(.A1(new_n302), .A2(KEYINPUT12), .A3(G68), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT12), .B1(new_n302), .B2(G68), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n332), .A2(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n379), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n283), .B1(new_n246), .B2(new_n247), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n388), .A2(KEYINPUT75), .A3(G232), .ZN(new_n389));
  OAI211_X1 g0189(.A(G232), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT75), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g0193(.A(G226), .B(new_n283), .C1(new_n250), .C2(new_n251), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G33), .A2(G97), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n274), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n291), .A2(G238), .A3(new_n296), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n295), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT13), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n400), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT13), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n396), .B1(new_n389), .B2(new_n392), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n402), .B(new_n403), .C1(new_n404), .C2(new_n274), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT14), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(new_n407), .A3(G169), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n401), .A2(G179), .A3(new_n405), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n407), .B1(new_n406), .B2(G169), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n387), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT76), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n401), .A2(G190), .A3(new_n405), .ZN(new_n414));
  INV_X1    g0214(.A(new_n387), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n371), .B1(new_n401), .B2(new_n405), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n413), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n417), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n419), .A2(KEYINPUT76), .A3(new_n415), .A4(new_n414), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n331), .A2(new_n374), .A3(new_n412), .A4(new_n421), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n388), .A2(G223), .B1(new_n252), .B2(G77), .ZN(new_n423));
  AOI21_X1  g0223(.A(G1698), .B1(new_n246), .B2(new_n247), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G222), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n355), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n359), .A2(G226), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n428), .A3(new_n295), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(new_n369), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(G200), .B2(new_n429), .ZN(new_n431));
  OAI21_X1  g0231(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n259), .A2(G150), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n432), .B(new_n433), .C1(new_n341), .C2(new_n311), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n376), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT70), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT70), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n376), .A2(new_n437), .A3(new_n434), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n303), .A2(new_n217), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n310), .A2(G50), .A3(new_n333), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n436), .A2(new_n438), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n441), .A2(KEYINPUT9), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(KEYINPUT9), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n431), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n441), .B(KEYINPUT9), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n429), .A2(G200), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT74), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT10), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n429), .B2(new_n369), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT74), .B1(new_n429), .B2(G200), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n448), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n444), .A2(KEYINPUT10), .B1(new_n445), .B2(new_n452), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n429), .A2(G179), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n429), .A2(new_n363), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n441), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n422), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT87), .ZN(new_n459));
  INV_X1    g0259(.A(G116), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(new_n312), .B2(G33), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n302), .B(new_n461), .C1(new_n269), .C2(new_n270), .ZN(new_n462));
  INV_X1    g0262(.A(new_n301), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n460), .A2(G20), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n267), .A2(new_n220), .B1(G20), .B2(new_n460), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  INV_X1    g0266(.A(G97), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n466), .B(new_n253), .C1(G33), .C2(new_n467), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n465), .A2(KEYINPUT20), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT20), .B1(new_n465), .B2(new_n468), .ZN(new_n470));
  OAI221_X1 g0270(.A(new_n462), .B1(new_n463), .B2(new_n464), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n312), .A2(G45), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(new_n291), .A3(G274), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n293), .A2(G1), .ZN(new_n478));
  INV_X1    g0278(.A(new_n475), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(new_n473), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n291), .A2(new_n480), .A3(G270), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT85), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n424), .A2(new_n483), .A3(G257), .ZN(new_n484));
  OAI211_X1 g0284(.A(G257), .B(new_n283), .C1(new_n250), .C2(new_n251), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT85), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(G264), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n488));
  INV_X1    g0288(.A(G303), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(new_n248), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n482), .B1(new_n492), .B2(new_n355), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n471), .B1(new_n493), .B2(G190), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n274), .B1(new_n487), .B2(new_n491), .ZN(new_n495));
  OAI21_X1  g0295(.A(G200), .B1(new_n495), .B2(new_n482), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n459), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n471), .ZN(new_n498));
  INV_X1    g0298(.A(new_n482), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n490), .B1(new_n484), .B2(new_n486), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n499), .B(G190), .C1(new_n500), .C2(new_n274), .ZN(new_n501));
  AND4_X1   g0301(.A1(new_n459), .A2(new_n496), .A3(new_n498), .A4(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n492), .A2(new_n355), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n363), .B1(new_n504), .B2(new_n499), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(KEYINPUT86), .A3(KEYINPUT21), .A4(new_n471), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT86), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n471), .B(G169), .C1(new_n495), .C2(new_n482), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT21), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n509), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n499), .B1(new_n500), .B2(new_n274), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(new_n365), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n471), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n506), .A2(new_n510), .A3(new_n511), .A4(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n503), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n339), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n312), .A2(G33), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n310), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n517), .A2(new_n302), .ZN(new_n520));
  XNOR2_X1  g0320(.A(KEYINPUT82), .B(G87), .ZN(new_n521));
  NOR2_X1   g0321(.A1(G97), .A2(G107), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT19), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n253), .B1(new_n395), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n248), .A2(new_n253), .A3(G68), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n524), .B1(new_n341), .B2(new_n467), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n520), .B1(new_n529), .B2(new_n271), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n519), .A2(new_n530), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n293), .A2(G1), .A3(G274), .ZN(new_n532));
  AOI21_X1  g0332(.A(G250), .B1(new_n312), .B2(G45), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n534), .A2(KEYINPUT81), .A3(new_n291), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT81), .B1(new_n534), .B2(new_n291), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(G238), .B(new_n283), .C1(new_n250), .C2(new_n251), .ZN(new_n538));
  OAI211_X1 g0338(.A(G244), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n539));
  INV_X1    g0339(.A(G33), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(new_n460), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n355), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n537), .A2(new_n365), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT81), .ZN(new_n546));
  INV_X1    g0346(.A(G274), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n312), .A2(new_n547), .A3(G45), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n478), .B2(G250), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n546), .B1(new_n358), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n534), .A2(KEYINPUT81), .A3(new_n291), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n544), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n363), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n531), .A2(new_n545), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(G200), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n375), .A2(G87), .A3(new_n302), .A4(new_n518), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n530), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT84), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n544), .A2(G190), .A3(new_n550), .A4(new_n551), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT83), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT83), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n537), .A2(new_n561), .A3(G190), .A4(new_n544), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n557), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n560), .A2(new_n562), .A3(KEYINPUT84), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n554), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n291), .A2(new_n480), .A3(G257), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT80), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT80), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n291), .A2(new_n480), .A3(new_n569), .A4(G257), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(G250), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n572));
  OAI211_X1 g0372(.A(G244), .B(new_n283), .C1(new_n250), .C2(new_n251), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT4), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n466), .B(new_n572), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT4), .B1(new_n424), .B2(G244), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n355), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n571), .A2(new_n577), .A3(new_n477), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G200), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n302), .A2(G97), .ZN(new_n580));
  OAI21_X1  g0380(.A(G107), .B1(new_n263), .B2(new_n264), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n259), .A2(G77), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT6), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n583), .A2(G97), .A3(G107), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n467), .A2(KEYINPUT6), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT79), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n586), .A2(G107), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n352), .A2(KEYINPUT79), .ZN(new_n588));
  OAI22_X1  g0388(.A1(new_n584), .A2(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n522), .A2(KEYINPUT6), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n583), .A2(G97), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n352), .A2(KEYINPUT79), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n586), .A2(G107), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n590), .A2(new_n591), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n589), .A2(G20), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n581), .A2(new_n582), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n580), .B1(new_n596), .B2(new_n271), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n310), .A2(G97), .A3(new_n518), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n571), .A2(new_n577), .A3(G190), .A4(new_n477), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n579), .A2(new_n597), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n595), .A2(new_n582), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n352), .B1(new_n249), .B2(new_n254), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n271), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n580), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n598), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n578), .A2(new_n363), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n571), .A2(new_n577), .A3(new_n365), .A4(new_n477), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n600), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(G250), .B(new_n283), .C1(new_n250), .C2(new_n251), .ZN(new_n610));
  OAI211_X1 g0410(.A(G257), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n611));
  INV_X1    g0411(.A(G294), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n610), .B(new_n611), .C1(new_n540), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n355), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT89), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT89), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n613), .A2(new_n616), .A3(new_n355), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n291), .A2(new_n480), .A3(G264), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n477), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n615), .A2(new_n369), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n614), .A2(new_n477), .A3(new_n618), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n371), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT24), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n253), .B(G87), .C1(new_n250), .C2(new_n251), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT22), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT22), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n248), .A2(new_n627), .A3(new_n253), .A4(G87), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT23), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n253), .B2(G107), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n352), .A2(KEYINPUT23), .A3(G20), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n541), .A2(new_n253), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(KEYINPUT88), .B(new_n624), .C1(new_n629), .C2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n635), .B1(new_n626), .B2(new_n628), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT88), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT24), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI211_X1 g0439(.A(KEYINPUT88), .B(new_n635), .C1(new_n626), .C2(new_n628), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n636), .B(new_n271), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n303), .A2(new_n352), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n642), .B(KEYINPUT25), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n375), .A2(new_n302), .A3(new_n518), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n644), .B2(G107), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n623), .A2(new_n641), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n619), .A2(new_n617), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n616), .B1(new_n613), .B2(new_n355), .ZN(new_n648));
  OAI21_X1  g0448(.A(G169), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n614), .A2(G179), .A3(new_n477), .A4(new_n618), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n641), .A2(new_n645), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n609), .A2(new_n646), .A3(new_n651), .ZN(new_n652));
  AND4_X1   g0452(.A1(new_n458), .A2(new_n516), .A3(new_n566), .A4(new_n652), .ZN(G372));
  INV_X1    g0453(.A(KEYINPUT90), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n655), .B1(new_n566), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n553), .A2(new_n545), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n531), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n530), .A2(new_n556), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n563), .A2(new_n555), .A3(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n656), .A2(new_n655), .A3(new_n659), .A4(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n659), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n654), .B1(new_n657), .B2(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n662), .A2(new_n659), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n563), .A2(new_n558), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n555), .A2(new_n530), .A3(new_n556), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n565), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(new_n659), .A3(new_n656), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT26), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n665), .A2(KEYINPUT90), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n515), .A2(new_n651), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n667), .A2(new_n563), .B1(new_n658), .B2(new_n531), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n623), .A2(new_n641), .A3(new_n645), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n673), .A2(new_n674), .A3(new_n608), .A4(new_n600), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n664), .A2(new_n671), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n458), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g0479(.A(new_n679), .B(KEYINPUT91), .Z(new_n680));
  AND3_X1   g0480(.A1(new_n322), .A2(new_n325), .A3(new_n321), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n326), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n419), .A2(new_n415), .A3(new_n414), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n347), .A2(new_n364), .A3(new_n366), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n412), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n318), .B(KEYINPUT17), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n683), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n456), .B1(new_n689), .B2(new_n453), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n680), .A2(new_n691), .ZN(G369));
  OR3_X1    g0492(.A1(new_n463), .A2(KEYINPUT27), .A3(G20), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT27), .B1(new_n463), .B2(G20), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G213), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n516), .B1(new_n498), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n498), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n515), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n641), .A2(new_n645), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n649), .A2(new_n650), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n697), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n707), .A3(new_n674), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n651), .A2(new_n697), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n708), .A2(KEYINPUT92), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT92), .B1(new_n708), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n703), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n706), .A2(new_n697), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n708), .A2(new_n709), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT92), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n708), .A2(KEYINPUT92), .A3(new_n709), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n515), .A2(new_n698), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n715), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n714), .A2(new_n723), .ZN(G399));
  INV_X1    g0524(.A(new_n224), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G41), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n218), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n726), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G1), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n521), .A2(new_n460), .A3(new_n522), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n727), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n678), .A2(new_n698), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n733), .A2(KEYINPUT29), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n614), .A2(new_n618), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n552), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(G179), .A3(new_n493), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n735), .B1(new_n738), .B2(new_n578), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n512), .A2(new_n365), .A3(new_n552), .A4(new_n621), .ZN(new_n740));
  INV_X1    g0540(.A(new_n578), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT93), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n552), .A2(new_n365), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n493), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT93), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n744), .A2(new_n745), .A3(new_n621), .A4(new_n578), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n513), .A2(KEYINPUT30), .A3(new_n741), .A4(new_n737), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n739), .A2(new_n742), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n697), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT31), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n739), .B(new_n747), .C1(new_n741), .C2(new_n740), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n698), .A2(new_n750), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n749), .A2(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n516), .A2(new_n652), .A3(new_n566), .A4(new_n698), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n673), .A2(new_n656), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n554), .B1(new_n757), .B2(KEYINPUT26), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n758), .B1(KEYINPUT26), .B2(new_n669), .C1(new_n672), .C2(new_n675), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n698), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT29), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n734), .A2(new_n756), .A3(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n732), .B1(new_n763), .B2(G1), .ZN(G364));
  INV_X1    g0564(.A(G330), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n699), .B2(new_n701), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n300), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n312), .B1(new_n767), .B2(G45), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n726), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(G330), .B2(new_n702), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n725), .A2(new_n252), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G355), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(G116), .B2(new_n224), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n219), .A2(new_n293), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n252), .A2(new_n224), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n241), .B2(G45), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n775), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n220), .B1(G20), .B2(new_n363), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n770), .B1(new_n779), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n365), .A2(new_n371), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT95), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n369), .A2(G20), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT94), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(KEYINPUT96), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(KEYINPUT96), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(KEYINPUT98), .B1(new_n371), .B2(G179), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR3_X1   g0598(.A1(new_n371), .A2(KEYINPUT98), .A3(G179), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n791), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT99), .Z(new_n802));
  AOI22_X1  g0602(.A1(new_n796), .A2(G329), .B1(new_n802), .B2(G283), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n253), .A2(new_n365), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n804), .A2(new_n369), .A3(new_n371), .ZN(new_n805));
  INV_X1    g0605(.A(G311), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n789), .A2(new_n365), .A3(new_n371), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(KEYINPUT33), .B(G317), .Z(new_n809));
  OAI221_X1 g0609(.A(new_n252), .B1(new_n805), .B2(new_n806), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n804), .A2(G190), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n371), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G326), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n811), .A2(G200), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G322), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n813), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n800), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n253), .A2(new_n369), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n810), .B(new_n817), .C1(G303), .C2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(G20), .B1(new_n788), .B2(new_n369), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n803), .B(new_n822), .C1(new_n612), .C2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G159), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n795), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(KEYINPUT97), .B(KEYINPUT32), .Z(new_n828));
  XOR2_X1   g0628(.A(new_n827), .B(new_n828), .Z(new_n829));
  NOR2_X1   g0629(.A1(new_n824), .A2(new_n467), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n820), .A2(new_n521), .ZN(new_n831));
  INV_X1    g0631(.A(new_n812), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n815), .A2(new_n256), .B1(new_n832), .B2(new_n217), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n248), .B1(new_n805), .B2(new_n345), .C1(new_n808), .C2(new_n244), .ZN(new_n834));
  NOR4_X1   g0634(.A1(new_n830), .A2(new_n831), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n802), .A2(G107), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n825), .B1(new_n829), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n786), .B1(new_n838), .B2(new_n783), .ZN(new_n839));
  INV_X1    g0639(.A(new_n782), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n702), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n772), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G396));
  NAND2_X1  g0643(.A1(new_n367), .A2(new_n698), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n698), .B1(new_n336), .B2(new_n346), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n373), .B2(new_n368), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n844), .B1(new_n846), .B2(new_n367), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n733), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n686), .A2(new_n697), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n373), .A2(new_n368), .ZN(new_n850));
  INV_X1    g0650(.A(new_n845), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n849), .B1(new_n852), .B2(new_n686), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n678), .A2(new_n698), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n848), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n770), .B1(new_n855), .B2(new_n756), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n756), .B2(new_n855), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n796), .A2(G311), .ZN(new_n858));
  INV_X1    g0658(.A(G283), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n252), .B1(new_n805), .B2(new_n460), .C1(new_n808), .C2(new_n859), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n815), .A2(new_n612), .B1(new_n832), .B2(new_n489), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n860), .B(new_n861), .C1(G107), .C2(new_n821), .ZN(new_n862));
  INV_X1    g0662(.A(new_n830), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n802), .A2(G87), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n858), .A2(new_n862), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n802), .A2(G68), .ZN(new_n866));
  INV_X1    g0666(.A(new_n805), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n867), .A2(G159), .B1(new_n807), .B2(G150), .ZN(new_n868));
  INV_X1    g0668(.A(G143), .ZN(new_n869));
  INV_X1    g0669(.A(G137), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n868), .B1(new_n815), .B2(new_n869), .C1(new_n870), .C2(new_n832), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT34), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n866), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n252), .B1(new_n821), .B2(G50), .ZN(new_n876));
  INV_X1    g0676(.A(G132), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n876), .B1(new_n256), .B2(new_n824), .C1(new_n795), .C2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n865), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n783), .ZN(new_n880));
  INV_X1    g0680(.A(new_n770), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n783), .A2(new_n780), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n881), .B1(new_n345), .B2(new_n882), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n880), .B(new_n883), .C1(new_n853), .C2(new_n781), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n857), .A2(new_n884), .ZN(G384));
  NOR3_X1   g0685(.A1(new_n220), .A2(new_n253), .A3(new_n460), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n589), .A2(new_n594), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT35), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n888), .B2(new_n887), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT36), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n218), .B(G77), .C1(new_n256), .C2(new_n244), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n217), .A2(G68), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n312), .B(G13), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n262), .A2(new_n266), .A3(new_n376), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n314), .ZN(new_n898));
  INV_X1    g0698(.A(new_n695), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n325), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(new_n318), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n322), .A2(new_n325), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n322), .A2(new_n899), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n904), .A2(new_n905), .A3(new_n906), .A4(new_n318), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n900), .B1(new_n688), .B2(new_n682), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n896), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  INV_X1    g0711(.A(new_n900), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n330), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n903), .A2(new_n907), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(KEYINPUT38), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n910), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n749), .A2(new_n750), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n748), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n754), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n410), .A2(new_n411), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n421), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n415), .A2(new_n698), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n922), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n412), .A2(new_n684), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n847), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(KEYINPUT101), .A2(KEYINPUT40), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n916), .A2(new_n919), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n905), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n330), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n904), .A2(new_n905), .A3(new_n318), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT37), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n907), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n330), .A2(new_n912), .B1(new_n903), .B2(new_n907), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n934), .A2(new_n935), .B1(new_n936), .B2(KEYINPUT38), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n406), .A2(G169), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT14), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(new_n409), .A3(new_n408), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n418), .B2(new_n420), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n925), .B1(new_n941), .B2(new_n924), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n919), .A2(new_n853), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n937), .B1(new_n943), .B2(KEYINPUT101), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n928), .B1(new_n944), .B2(new_n911), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n458), .A2(new_n919), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT102), .ZN(new_n948));
  OAI21_X1  g0748(.A(G330), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n948), .B2(new_n946), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n910), .A2(KEYINPUT39), .A3(new_n915), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n940), .A2(new_n387), .A3(new_n698), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n951), .B(new_n953), .C1(new_n937), .C2(KEYINPUT39), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n683), .A2(new_n695), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n910), .A2(new_n915), .ZN(new_n957));
  INV_X1    g0757(.A(new_n942), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n854), .B2(new_n844), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n956), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n761), .B1(KEYINPUT29), .B2(new_n733), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n458), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n691), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n960), .B(new_n963), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n950), .A2(new_n964), .B1(new_n312), .B2(new_n767), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n950), .A2(new_n964), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n895), .B1(new_n965), .B2(new_n966), .ZN(G367));
  NAND2_X1  g0767(.A1(new_n605), .A2(new_n697), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n600), .A2(new_n608), .A3(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT105), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n656), .A2(new_n697), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n600), .A2(new_n608), .A3(KEYINPUT105), .A4(new_n968), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT106), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT106), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n971), .A2(new_n976), .A3(new_n972), .A4(new_n973), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n722), .B1(new_n710), .B2(new_n711), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n979), .A2(KEYINPUT42), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n706), .B1(new_n975), .B2(new_n977), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n698), .B1(new_n982), .B2(new_n656), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT42), .B1(new_n979), .B2(new_n980), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n659), .B(new_n661), .C1(new_n660), .C2(new_n698), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(KEYINPUT103), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(KEYINPUT103), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n659), .A2(new_n660), .A3(new_n698), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT104), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n994));
  AND3_X1   g0794(.A1(new_n985), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n993), .B1(new_n985), .B2(new_n994), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n995), .A2(new_n996), .B1(new_n714), .B2(new_n979), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n985), .A2(new_n994), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n992), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n714), .A2(new_n979), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n985), .A2(new_n993), .A3(new_n994), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n726), .B(KEYINPUT41), .Z(new_n1004));
  NAND2_X1  g0804(.A1(new_n712), .A2(new_n721), .ZN(new_n1005));
  AND3_X1   g0805(.A1(new_n1005), .A2(new_n766), .A3(new_n980), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n766), .B1(new_n1005), .B2(new_n980), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1008), .A2(new_n756), .A3(new_n734), .A4(new_n761), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n723), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n715), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n980), .A2(new_n978), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1011), .A2(new_n1015), .B1(KEYINPUT107), .B2(new_n713), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n713), .A2(KEYINPUT107), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT44), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n723), .B2(new_n978), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n980), .A2(new_n1012), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1021), .A2(KEYINPUT44), .A3(new_n979), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  AND3_X1   g0823(.A1(new_n1016), .A2(new_n1018), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1018), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1010), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1004), .B1(new_n1026), .B2(new_n763), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1003), .B1(new_n1027), .B2(new_n769), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n784), .B1(new_n224), .B2(new_n339), .C1(new_n234), .C2(new_n777), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n770), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n796), .A2(G137), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n248), .B1(new_n808), .B2(new_n826), .ZN(new_n1032));
  INV_X1    g0832(.A(G150), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n815), .A2(new_n1033), .B1(new_n832), .B2(new_n869), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1032), .B(new_n1034), .C1(G50), .C2(new_n867), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n823), .A2(G68), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n821), .A2(G58), .B1(G77), .B2(new_n801), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1031), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n821), .A2(G116), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT46), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n248), .B1(new_n807), .B2(G294), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n815), .B2(new_n489), .C1(new_n806), .C2(new_n832), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G97), .B2(new_n801), .ZN(new_n1043));
  INV_X1    g0843(.A(G317), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1040), .B(new_n1043), .C1(new_n1044), .C2(new_n795), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n823), .A2(G107), .B1(G283), .B2(new_n867), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT108), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1038), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g0848(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n1049));
  XNOR2_X1  g0849(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1030), .B1(new_n1050), .B2(new_n783), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n990), .A2(new_n840), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1028), .A2(new_n1053), .ZN(G387));
  NAND2_X1  g0854(.A1(new_n1008), .A2(new_n769), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n801), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n252), .B1(new_n1056), .B2(new_n460), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n867), .A2(G303), .B1(new_n807), .B2(G311), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n815), .B2(new_n1044), .C1(new_n816), .C2(new_n832), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT48), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n859), .B2(new_n824), .C1(new_n612), .C2(new_n820), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT49), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1057), .B(new_n1065), .C1(G326), .C2(new_n796), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n795), .A2(new_n1033), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n808), .A2(new_n311), .B1(new_n805), .B2(new_n244), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n820), .A2(new_n345), .B1(new_n1068), .B2(KEYINPUT111), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(KEYINPUT111), .B2(new_n1068), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n823), .A2(new_n517), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n248), .B1(new_n815), .B2(new_n217), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G159), .B2(new_n812), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1067), .B(new_n1074), .C1(G97), .C2(new_n802), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n783), .B1(new_n1066), .B2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n773), .A2(new_n730), .B1(new_n352), .B2(new_n725), .ZN(new_n1077));
  AOI211_X1 g0877(.A(G45), .B(new_n730), .C1(G68), .C2(G77), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n311), .A2(G50), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT50), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n777), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT110), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n1081), .A2(new_n1082), .B1(new_n293), .B2(new_n231), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1077), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n881), .B1(new_n1085), .B2(new_n784), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1076), .B(new_n1086), .C1(new_n720), .C2(new_n840), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n763), .A2(new_n1008), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1009), .A2(new_n726), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1055), .B(new_n1087), .C1(new_n1088), .C2(new_n1089), .ZN(G393));
  INV_X1    g0890(.A(KEYINPUT107), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1091), .B(new_n714), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1016), .A2(new_n1018), .A3(new_n1023), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n1009), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1026), .A2(new_n1096), .A3(new_n726), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n979), .A2(new_n782), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n238), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n784), .B1(new_n467), .B2(new_n224), .C1(new_n1100), .C2(new_n777), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n770), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n796), .A2(G322), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n252), .B1(new_n805), .B2(new_n612), .C1(new_n808), .C2(new_n489), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n820), .A2(new_n859), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(G116), .C2(new_n823), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n814), .A2(G311), .B1(new_n812), .B2(G317), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT52), .Z(new_n1108));
  NAND4_X1  g0908(.A1(new_n1103), .A2(new_n1106), .A3(new_n836), .A4(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n252), .B1(new_n821), .B2(G68), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n864), .B(new_n1110), .C1(new_n869), .C2(new_n795), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT112), .Z(new_n1112));
  NAND2_X1  g0912(.A1(new_n823), .A2(G77), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n217), .B2(new_n808), .C1(new_n311), .C2(new_n805), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1114), .A2(KEYINPUT113), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(KEYINPUT113), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n814), .A2(G159), .B1(new_n812), .B2(G150), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT51), .Z(new_n1118));
  NAND3_X1  g0918(.A1(new_n1115), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1109), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1102), .B1(new_n1120), .B2(new_n783), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1098), .A2(new_n769), .B1(new_n1099), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1097), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(KEYINPUT114), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT114), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1097), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(G390));
  OAI21_X1  g0927(.A(new_n951), .B1(new_n937), .B2(KEYINPUT39), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n959), .B2(new_n953), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n846), .A2(new_n367), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n844), .B1(new_n760), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n942), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n935), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n930), .B2(new_n933), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n915), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n952), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1132), .A2(new_n1138), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n756), .A2(new_n847), .A3(new_n958), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1129), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n919), .A2(new_n942), .A3(G330), .A4(new_n853), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1129), .B2(new_n1139), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1128), .A2(new_n780), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n882), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1147), .A2(new_n337), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n866), .B1(new_n612), .B2(new_n795), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n821), .A2(G87), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n252), .B1(new_n808), .B2(new_n352), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G97), .B2(new_n867), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n814), .A2(G116), .B1(new_n812), .B2(G283), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1150), .A2(new_n1152), .A3(new_n1113), .A4(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1149), .A2(new_n1154), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1155), .A2(KEYINPUT118), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(KEYINPUT118), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT54), .B(G143), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n808), .A2(new_n870), .B1(new_n805), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n823), .B2(G159), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT117), .Z(new_n1161));
  NOR2_X1   g0961(.A1(new_n820), .A2(new_n1033), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT53), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n796), .A2(G125), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n812), .A2(G128), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1165), .B(new_n248), .C1(new_n815), .C2(new_n877), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G50), .B2(new_n801), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .A4(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1156), .A2(new_n1157), .A3(new_n1168), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n881), .B(new_n1148), .C1(new_n1169), .C2(new_n783), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1145), .A2(new_n769), .B1(new_n1146), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT116), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1129), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1137), .B1(new_n1131), .B2(new_n942), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n665), .A2(new_n670), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n676), .B1(new_n1175), .B2(new_n654), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n697), .B1(new_n1176), .B2(new_n671), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n849), .B1(new_n1177), .B2(new_n853), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n952), .B1(new_n1178), .B2(new_n958), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1174), .B1(new_n1179), .B2(new_n1128), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1173), .B1(new_n1180), .B2(new_n1143), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1140), .A2(new_n1131), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n919), .A2(G330), .A3(new_n853), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n958), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n765), .B(new_n847), .C1(new_n753), .C2(new_n754), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1143), .B1(new_n1186), .B2(new_n942), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n854), .A2(new_n844), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n1188), .A3(KEYINPUT115), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(KEYINPUT115), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1185), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n458), .A2(G330), .A3(new_n919), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n962), .A2(new_n691), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1172), .B(new_n726), .C1(new_n1181), .C2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1181), .A2(new_n1195), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n962), .A2(new_n691), .A3(new_n1193), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT115), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1189), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1199), .B1(new_n1203), .B2(new_n1185), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1144), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n1173), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1172), .B1(new_n1206), .B2(new_n726), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1171), .B1(new_n1198), .B2(new_n1207), .ZN(G378));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1199), .B1(new_n1145), .B2(new_n1192), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n441), .A2(new_n899), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT120), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n453), .B2(new_n457), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n445), .A2(new_n452), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n449), .B1(new_n445), .B2(new_n431), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n456), .B(new_n1212), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1217));
  XOR2_X1   g1017(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1218));
  AND3_X1   g1018(.A1(new_n1214), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1218), .B1(new_n1214), .B2(new_n1217), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT101), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n926), .B2(new_n919), .ZN(new_n1223));
  OAI21_X1  g1023(.A(KEYINPUT40), .B1(new_n1223), .B2(new_n937), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n765), .B(new_n1221), .C1(new_n1224), .C2(new_n928), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1221), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n945), .B2(G330), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n959), .A2(new_n957), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(new_n955), .A3(new_n954), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1225), .A2(new_n1227), .A3(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n754), .A2(new_n917), .A3(new_n918), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n924), .B1(new_n421), .B2(new_n920), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n684), .A2(new_n924), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n940), .B2(new_n387), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n853), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(KEYINPUT101), .B1(new_n1231), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n911), .B1(new_n1236), .B2(new_n1136), .ZN(new_n1237));
  AND4_X1   g1037(.A1(new_n919), .A2(new_n916), .A3(new_n926), .A4(new_n927), .ZN(new_n1238));
  OAI21_X1  g1038(.A(G330), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1221), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n945), .A2(G330), .A3(new_n1226), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n960), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1230), .A2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1209), .B1(new_n1210), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1194), .B1(new_n1181), .B2(new_n1195), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1229), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1240), .A2(new_n960), .A3(new_n1241), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1209), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n728), .B1(new_n1245), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1244), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1221), .A2(new_n780), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n770), .B1(G50), .B2(new_n1147), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n867), .A2(new_n517), .B1(new_n807), .B2(G97), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n460), .B2(new_n832), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G107), .B2(new_n814), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1056), .A2(new_n256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(new_n1036), .A3(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n292), .B(new_n252), .C1(new_n820), .C2(new_n345), .ZN(new_n1260));
  XOR2_X1   g1060(.A(new_n1260), .B(KEYINPUT119), .Z(new_n1261));
  AOI211_X1 g1061(.A(new_n1259), .B(new_n1261), .C1(G283), .C2(new_n796), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1262), .A2(KEYINPUT58), .ZN(new_n1263));
  AOI21_X1  g1063(.A(G50), .B1(new_n540), .B2(new_n292), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n248), .B2(G41), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1262), .A2(KEYINPUT58), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n808), .A2(new_n877), .B1(new_n805), .B2(new_n870), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n812), .A2(G125), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1267), .B(new_n1268), .C1(G128), .C2(new_n814), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n1269), .B1(new_n1033), .B2(new_n824), .C1(new_n820), .C2(new_n1158), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1270), .A2(KEYINPUT59), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(KEYINPUT59), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n796), .A2(G124), .ZN(new_n1273));
  AOI211_X1 g1073(.A(G33), .B(G41), .C1(new_n801), .C2(G159), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1263), .A2(new_n1265), .A3(new_n1266), .A4(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1253), .B1(new_n1276), .B2(new_n783), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1251), .A2(new_n769), .B1(new_n1252), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1250), .A2(new_n1278), .ZN(G375));
  INV_X1    g1079(.A(new_n1004), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1203), .A2(new_n1199), .A3(new_n1185), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1195), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n796), .A2(G128), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n248), .B1(new_n808), .B2(new_n1158), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n815), .A2(new_n870), .B1(new_n832), .B2(new_n877), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n1284), .B(new_n1285), .C1(G150), .C2(new_n867), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n823), .A2(G50), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1257), .B1(G159), .B2(new_n821), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1283), .A2(new_n1286), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n796), .A2(G303), .ZN(new_n1290));
  OAI221_X1 g1090(.A(new_n252), .B1(new_n805), .B2(new_n352), .C1(new_n808), .C2(new_n460), .ZN(new_n1291));
  OAI22_X1  g1091(.A1(new_n815), .A2(new_n859), .B1(new_n832), .B2(new_n612), .ZN(new_n1292));
  AOI211_X1 g1092(.A(new_n1291), .B(new_n1292), .C1(G97), .C2(new_n821), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n802), .A2(G77), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1290), .A2(new_n1293), .A3(new_n1071), .A4(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1289), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n783), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1297), .B(new_n770), .C1(G68), .C2(new_n1147), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1298), .B1(new_n958), .B2(new_n780), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1299), .B1(new_n1192), .B2(new_n769), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1282), .A2(new_n1300), .ZN(G381));
  OR3_X1    g1101(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1302));
  NOR4_X1   g1102(.A1(G390), .A2(G387), .A3(G381), .A4(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(G378), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1303), .A2(new_n1304), .A3(new_n1250), .A4(new_n1278), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1305), .B(KEYINPUT121), .ZN(G407));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n696), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G407), .B(G213), .C1(G375), .C2(new_n1307), .ZN(G409));
  INV_X1    g1108(.A(new_n1126), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1125), .B1(new_n1097), .B2(new_n1122), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n997), .A2(new_n1002), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1009), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1280), .B1(new_n1312), .B2(new_n762), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1311), .B1(new_n1313), .B2(new_n768), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1053), .ZN(new_n1315));
  OAI22_X1  g1115(.A1(new_n1309), .A2(new_n1310), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1124), .A2(new_n1028), .A3(new_n1053), .A4(new_n1126), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1317), .A3(KEYINPUT124), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(G393), .B(new_n842), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1319), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1316), .A2(new_n1317), .A3(KEYINPUT124), .A4(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT61), .ZN(new_n1325));
  INV_X1    g1125(.A(G213), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1326), .A2(G343), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(G2897), .ZN(new_n1328));
  XOR2_X1   g1128(.A(new_n1328), .B(KEYINPUT123), .Z(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT60), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1281), .A2(new_n1331), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1203), .A2(new_n1199), .A3(KEYINPUT60), .A4(new_n1185), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1332), .A2(new_n1333), .A3(new_n726), .A4(new_n1195), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1334), .A2(G384), .A3(new_n1300), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(G384), .B1(new_n1334), .B2(new_n1300), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1330), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1334), .A2(new_n1300), .ZN(new_n1339));
  INV_X1    g1139(.A(G384), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1341), .A2(new_n1335), .A3(new_n1329), .ZN(new_n1342));
  AND2_X1   g1142(.A1(new_n1338), .A2(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(G378), .A2(new_n1250), .A3(new_n1278), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n726), .B1(new_n1181), .B2(new_n1195), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(KEYINPUT116), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1346), .A2(new_n1197), .A3(new_n1196), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1245), .A2(new_n1280), .A3(new_n1251), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(new_n1278), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1347), .A2(new_n1349), .A3(new_n1171), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1327), .B1(new_n1344), .B2(new_n1350), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1325), .B1(new_n1343), .B2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT62), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1353), .B1(new_n1351), .B2(new_n1354), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1352), .A2(new_n1355), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1351), .A2(new_n1353), .A3(new_n1354), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1324), .B1(new_n1356), .B2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1344), .A2(new_n1350), .ZN(new_n1359));
  INV_X1    g1159(.A(new_n1327), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1359), .A2(new_n1360), .A3(new_n1354), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT63), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  AND3_X1   g1163(.A1(new_n1320), .A2(new_n1325), .A3(new_n1322), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1351), .A2(KEYINPUT63), .A3(new_n1354), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1363), .A2(new_n1364), .A3(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT122), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1367), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1368));
  AOI211_X1 g1168(.A(KEYINPUT122), .B(new_n1327), .C1(new_n1344), .C2(new_n1350), .ZN(new_n1369));
  NOR3_X1   g1169(.A1(new_n1368), .A2(new_n1369), .A3(new_n1343), .ZN(new_n1370));
  NOR2_X1   g1170(.A1(new_n1366), .A2(new_n1370), .ZN(new_n1371));
  OAI21_X1  g1171(.A(KEYINPUT125), .B1(new_n1358), .B2(new_n1371), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1320), .A2(new_n1325), .A3(new_n1322), .ZN(new_n1373));
  AOI21_X1  g1173(.A(new_n1373), .B1(new_n1362), .B2(new_n1361), .ZN(new_n1374));
  OR2_X1    g1174(.A1(new_n1369), .A2(new_n1343), .ZN(new_n1375));
  OAI211_X1 g1175(.A(new_n1374), .B(new_n1365), .C1(new_n1375), .C2(new_n1368), .ZN(new_n1376));
  OR2_X1    g1176(.A1(new_n1343), .A2(new_n1351), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1361), .A2(KEYINPUT62), .ZN(new_n1378));
  NAND4_X1  g1178(.A1(new_n1377), .A2(new_n1378), .A3(new_n1325), .A4(new_n1357), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1379), .A2(new_n1323), .ZN(new_n1380));
  INV_X1    g1180(.A(KEYINPUT125), .ZN(new_n1381));
  NAND3_X1  g1181(.A1(new_n1376), .A2(new_n1380), .A3(new_n1381), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1372), .A2(new_n1382), .ZN(G405));
  NAND2_X1  g1183(.A1(G375), .A2(new_n1304), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1384), .A2(new_n1344), .ZN(new_n1385));
  OR2_X1    g1185(.A1(new_n1385), .A2(new_n1354), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1385), .A2(new_n1354), .ZN(new_n1387));
  OAI211_X1 g1187(.A(new_n1386), .B(new_n1387), .C1(KEYINPUT126), .C2(new_n1323), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1323), .A2(KEYINPUT126), .ZN(new_n1389));
  XOR2_X1   g1189(.A(new_n1388), .B(new_n1389), .Z(G402));
endmodule


