//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G58), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(KEYINPUT64), .B(KEYINPUT2), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT65), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n215), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT70), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n206), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n251), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n206), .A2(G20), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(G68), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n219), .A2(G20), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n207), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI221_X1 g0063(.A(new_n259), .B1(new_n260), .B2(new_n261), .C1(new_n263), .C2(new_n202), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT11), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n264), .A2(new_n265), .A3(new_n251), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n265), .B1(new_n264), .B2(new_n251), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n258), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n254), .A2(new_n255), .ZN(new_n269));
  OAI21_X1  g0069(.A(KEYINPUT12), .B1(new_n269), .B2(G68), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT74), .ZN(new_n271));
  INV_X1    g0071(.A(G13), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G1), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OR3_X1    g0074(.A1(new_n274), .A2(KEYINPUT12), .A3(new_n259), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n268), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT14), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  INV_X1    g0078(.A(G226), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n226), .A2(G1698), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n281), .B(new_n282), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G97), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G1), .A3(G13), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G41), .ZN(new_n292));
  INV_X1    g0092(.A(G45), .ZN(new_n293));
  AOI21_X1  g0093(.A(G1), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n294), .A2(new_n289), .A3(G274), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n289), .A2(G238), .A3(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n278), .B1(new_n291), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n289), .B1(new_n285), .B2(new_n286), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n295), .A2(new_n297), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT13), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n277), .B(G169), .C1(new_n299), .C2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n291), .A2(new_n298), .A3(new_n278), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT13), .B1(new_n300), .B2(new_n301), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(G179), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n305), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n277), .B1(new_n308), .B2(G169), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT75), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n299), .A2(new_n302), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT14), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT75), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n313), .A2(new_n314), .A3(new_n306), .A4(new_n303), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n276), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n311), .A2(G190), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n308), .A2(G200), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n276), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT66), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT3), .ZN(new_n323));
  INV_X1    g0123(.A(G33), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(KEYINPUT3), .A2(G33), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n322), .B1(new_n327), .B2(G1698), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n322), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(G238), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n283), .A2(new_n284), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(G1698), .ZN(new_n333));
  INV_X1    g0133(.A(G107), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT67), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT67), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G107), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n333), .A2(G232), .B1(new_n338), .B2(new_n332), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n289), .B1(new_n331), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n295), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n290), .A2(new_n294), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(G244), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT68), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(G1698), .B1(new_n283), .B2(new_n284), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT66), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n220), .B1(new_n347), .B2(new_n329), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n327), .A2(new_n280), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT67), .B(G107), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n349), .A2(new_n226), .B1(new_n327), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n290), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT68), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(new_n353), .A3(new_n343), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n345), .A2(new_n354), .A3(new_n312), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT8), .B(G58), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(new_n262), .B1(G20), .B2(G77), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n260), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n251), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n256), .A2(G77), .A3(new_n257), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n361), .B(new_n362), .C1(G77), .C2(new_n269), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n355), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT71), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT71), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n355), .A2(new_n366), .A3(new_n363), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n345), .A2(new_n354), .ZN(new_n368));
  INV_X1    g0168(.A(G179), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n365), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n356), .B1(new_n206), .B2(G20), .ZN(new_n372));
  INV_X1    g0172(.A(new_n252), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n373), .A2(new_n251), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n372), .A2(new_n374), .B1(new_n356), .B2(new_n373), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n325), .A2(new_n207), .A3(new_n326), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT78), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n332), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n377), .B1(new_n376), .B2(new_n378), .ZN(new_n382));
  OAI21_X1  g0182(.A(G68), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(G58), .A2(G68), .ZN(new_n384));
  OAI21_X1  g0184(.A(G20), .B1(new_n384), .B2(new_n201), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT77), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n262), .A2(G159), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT77), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n388), .B(G20), .C1(new_n384), .C2(new_n201), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT16), .B1(new_n383), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n219), .B1(new_n376), .B2(KEYINPUT7), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n283), .A2(new_n284), .A3(G20), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n378), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n390), .A2(KEYINPUT16), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n251), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n375), .B1(new_n391), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G223), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n280), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n279), .A2(G1698), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n400), .B(new_n401), .C1(new_n283), .C2(new_n284), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G87), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n290), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n289), .A2(G232), .A3(new_n296), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n295), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n405), .A2(new_n407), .A3(new_n369), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n289), .B1(new_n402), .B2(new_n403), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n295), .A2(new_n406), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n312), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT79), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT79), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n408), .A2(new_n414), .A3(new_n411), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n398), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT18), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT18), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n398), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT80), .ZN(new_n422));
  INV_X1    g0222(.A(G190), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n405), .A2(new_n407), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G200), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n409), .B2(new_n410), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n409), .A2(new_n410), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n422), .B1(new_n428), .B2(new_n423), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT81), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n405), .A2(new_n407), .A3(new_n423), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT80), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT81), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n426), .A4(new_n424), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n375), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n383), .A2(new_n390), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT16), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n396), .A2(new_n251), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n435), .A2(new_n441), .A3(KEYINPUT17), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT17), .B1(new_n435), .B2(new_n441), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n321), .A2(new_n371), .A3(new_n421), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n251), .ZN(new_n446));
  INV_X1    g0246(.A(new_n260), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n357), .A2(new_n447), .B1(G150), .B2(new_n262), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n203), .A2(G20), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n374), .A2(G50), .A3(new_n257), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(G50), .B2(new_n252), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  OR3_X1    g0253(.A1(new_n453), .A2(KEYINPUT72), .A3(KEYINPUT9), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(KEYINPUT9), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT72), .B1(new_n453), .B2(KEYINPUT9), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n399), .B1(new_n347), .B2(new_n329), .ZN(new_n458));
  INV_X1    g0258(.A(G222), .ZN(new_n459));
  OAI22_X1  g0259(.A1(new_n349), .A2(new_n459), .B1(new_n261), .B2(new_n327), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n290), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n341), .B1(G226), .B2(new_n342), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G190), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(new_n425), .B2(new_n463), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n457), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT73), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT10), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(KEYINPUT10), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n467), .A2(KEYINPUT10), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n469), .B(new_n470), .C1(new_n457), .C2(new_n465), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n463), .A2(new_n369), .ZN(new_n472));
  OAI221_X1 g0272(.A(new_n472), .B1(G169), .B2(new_n463), .C1(new_n450), .C2(new_n452), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n340), .A2(new_n344), .A3(KEYINPUT68), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n353), .B1(new_n352), .B2(new_n343), .ZN(new_n475));
  OAI21_X1  g0275(.A(G190), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT69), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n368), .A2(KEYINPUT69), .A3(G190), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n368), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n363), .B1(new_n481), .B2(G200), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n468), .A2(new_n471), .A3(new_n473), .A4(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n445), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G303), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n289), .B1(new_n332), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(G257), .A2(G1698), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n280), .A2(G264), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n327), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT5), .B(G41), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n293), .A2(G1), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n492), .A2(G274), .A3(new_n289), .A4(new_n493), .ZN(new_n494));
  AND2_X1   g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  NOR2_X1   g0295(.A1(KEYINPUT5), .A2(G41), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(G270), .A3(new_n289), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n491), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(new_n312), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT20), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n207), .B1(new_n227), .B2(G33), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT84), .B1(G33), .B2(G283), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(KEYINPUT84), .A2(G33), .A3(G283), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G116), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G20), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n251), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n501), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(G20), .B1(new_n324), .B2(G97), .ZN(new_n511));
  INV_X1    g0311(.A(new_n505), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(new_n512), .B2(new_n503), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n513), .A2(KEYINPUT20), .A3(new_n251), .A4(new_n508), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n507), .B1(new_n206), .B2(G33), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n510), .A2(new_n514), .B1(new_n256), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT90), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT89), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n269), .B2(G116), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n254), .A2(KEYINPUT89), .A3(new_n507), .A4(new_n255), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n516), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n517), .B1(new_n516), .B2(new_n521), .ZN(new_n523));
  OAI211_X1 g0323(.A(KEYINPUT21), .B(new_n500), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n491), .A2(G179), .A3(new_n494), .A4(new_n498), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n522), .B2(new_n523), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n510), .A2(new_n514), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n256), .A2(new_n515), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n521), .ZN(new_n532));
  OAI21_X1  g0332(.A(KEYINPUT90), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n516), .A2(new_n517), .A3(new_n521), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT21), .B1(new_n535), .B2(new_n500), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n491), .A2(new_n494), .A3(new_n498), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(new_n423), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(G200), .B2(new_n537), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n539), .A2(new_n534), .A3(new_n533), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n528), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n497), .A2(G264), .A3(new_n289), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n222), .A2(new_n280), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n228), .A2(G1698), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n543), .B(new_n544), .C1(new_n283), .C2(new_n284), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G294), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT92), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n289), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(KEYINPUT92), .A3(new_n546), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n542), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(new_n369), .A3(new_n494), .ZN(new_n552));
  INV_X1    g0352(.A(new_n494), .ZN(new_n553));
  AOI211_X1 g0353(.A(new_n553), .B(new_n542), .C1(new_n549), .C2(new_n550), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n552), .B1(new_n554), .B2(G169), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n350), .A2(G20), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT23), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT22), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(KEYINPUT91), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n327), .A2(new_n207), .A3(G87), .A4(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n207), .B(G87), .C1(new_n283), .C2(new_n284), .ZN(new_n561));
  XNOR2_X1  g0361(.A(KEYINPUT91), .B(KEYINPUT22), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n334), .A2(G20), .ZN(new_n564));
  OAI22_X1  g0364(.A1(KEYINPUT23), .A2(new_n564), .B1(new_n260), .B2(new_n507), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n557), .A2(new_n560), .A3(new_n563), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT24), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n565), .B1(new_n556), .B2(KEYINPUT23), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT24), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n560), .A4(new_n563), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n446), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n274), .A2(new_n564), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n573), .B(KEYINPUT25), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n206), .A2(G33), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n252), .A2(new_n575), .A3(new_n215), .A4(new_n250), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n574), .B1(new_n334), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n555), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT93), .B1(new_n554), .B2(G200), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n551), .A2(new_n494), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT93), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n425), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n551), .A2(new_n423), .A3(new_n494), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n580), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n579), .B1(new_n578), .B2(new_n585), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n289), .A2(G274), .A3(new_n493), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G116), .ZN(new_n588));
  INV_X1    g0388(.A(G244), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G1698), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(G238), .B2(G1698), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n588), .B1(new_n591), .B2(new_n332), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n587), .B1(new_n592), .B2(new_n290), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT86), .B1(new_n293), .B2(G1), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT86), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(new_n206), .A3(G45), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n289), .A2(new_n594), .A3(new_n596), .A4(G250), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT87), .ZN(new_n598));
  AND2_X1   g0398(.A1(G1), .A2(G13), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n222), .B1(new_n599), .B2(new_n288), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT87), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n600), .A2(new_n601), .A3(new_n596), .A4(new_n594), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n593), .A2(new_n603), .A3(G190), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT88), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n598), .A2(new_n602), .ZN(new_n607));
  INV_X1    g0407(.A(new_n587), .ZN(new_n608));
  NOR2_X1   g0408(.A1(G238), .A2(G1698), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n589), .B2(G1698), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n610), .A2(new_n327), .B1(G33), .B2(G116), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n608), .B1(new_n611), .B2(new_n289), .ZN(new_n612));
  OAI21_X1  g0412(.A(G200), .B1(new_n607), .B2(new_n612), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n254), .A2(new_n255), .A3(new_n359), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n576), .A2(new_n221), .ZN(new_n615));
  NOR2_X1   g0415(.A1(G87), .A2(G97), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n335), .A2(new_n337), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT19), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n207), .B1(new_n286), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n327), .A2(new_n207), .A3(G68), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n618), .B1(new_n260), .B2(new_n227), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AOI211_X1 g0423(.A(new_n614), .B(new_n615), .C1(new_n623), .C2(new_n251), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n593), .A2(new_n603), .A3(KEYINPUT88), .A4(G190), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n606), .A2(new_n613), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n312), .B1(new_n607), .B2(new_n612), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n623), .A2(new_n251), .ZN(new_n628));
  INV_X1    g0428(.A(new_n614), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n576), .A2(new_n359), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n593), .A2(new_n603), .A3(new_n369), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n627), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n626), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n373), .A2(new_n227), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n576), .B2(new_n227), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n334), .A2(KEYINPUT6), .A3(G97), .ZN(new_n638));
  XNOR2_X1  g0438(.A(G97), .B(G107), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT6), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI22_X1  g0441(.A1(new_n641), .A2(new_n207), .B1(new_n261), .B2(new_n263), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT7), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT76), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT76), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT7), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT78), .B1(new_n393), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n380), .A3(new_n379), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n642), .B1(new_n649), .B2(new_n338), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n637), .B1(new_n650), .B2(new_n446), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n280), .B1(new_n325), .B2(new_n326), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n653), .A2(G250), .B1(new_n504), .B2(new_n505), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT83), .ZN(new_n655));
  OAI211_X1 g0455(.A(G244), .B(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT4), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XOR2_X1   g0458(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n659));
  NAND2_X1  g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n654), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n656), .A2(new_n655), .A3(new_n657), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n290), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n497), .A2(G257), .A3(new_n289), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n664), .A2(KEYINPUT85), .A3(new_n494), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT85), .B1(new_n664), .B2(new_n494), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n663), .A2(new_n667), .A3(new_n423), .ZN(new_n668));
  AOI21_X1  g0468(.A(G200), .B1(new_n663), .B2(new_n667), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n652), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n663), .A2(new_n667), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n312), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n663), .A2(new_n667), .A3(new_n369), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n651), .A3(new_n673), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n634), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  AND4_X1   g0475(.A1(new_n485), .A2(new_n541), .A3(new_n586), .A4(new_n675), .ZN(G372));
  NAND2_X1  g0476(.A1(new_n626), .A2(new_n633), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT26), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n613), .A2(new_n624), .A3(new_n604), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n633), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n651), .A2(new_n673), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n680), .A2(new_n681), .A3(new_n682), .A4(new_n672), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n678), .A2(new_n683), .A3(new_n633), .ZN(new_n684));
  AOI21_X1  g0484(.A(G200), .B1(new_n551), .B2(new_n494), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n584), .B1(new_n685), .B2(new_n582), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n554), .A2(KEYINPUT93), .A3(G200), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n578), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AND4_X1   g0488(.A1(new_n688), .A2(new_n674), .A3(new_n670), .A4(new_n680), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n500), .B1(new_n522), .B2(new_n523), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT21), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI221_X1 g0492(.A(new_n552), .B1(new_n554), .B2(G169), .C1(new_n572), .C2(new_n577), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n692), .A2(new_n693), .A3(new_n527), .A4(new_n524), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n684), .B1(new_n689), .B2(new_n694), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n695), .A2(new_n445), .A3(new_n484), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT94), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT95), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n365), .A2(new_n367), .A3(new_n370), .A4(new_n319), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n310), .A2(new_n315), .ZN(new_n700));
  INV_X1    g0500(.A(new_n276), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n435), .A2(new_n441), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT17), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n435), .A2(new_n441), .A3(KEYINPUT17), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n698), .B(new_n421), .C1(new_n703), .C2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n708), .B1(new_n699), .B2(new_n702), .ZN(new_n710));
  INV_X1    g0510(.A(new_n421), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT95), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n468), .A2(new_n471), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n709), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n714), .A2(new_n473), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n697), .A2(new_n715), .ZN(G369));
  NOR2_X1   g0516(.A1(new_n528), .A2(new_n536), .ZN(new_n717));
  OR3_X1    g0517(.A1(new_n274), .A2(KEYINPUT27), .A3(G20), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT27), .B1(new_n274), .B2(G20), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G213), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(G343), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n535), .A2(new_n722), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n541), .A2(new_n723), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  INV_X1    g0527(.A(new_n722), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n586), .B1(new_n578), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n579), .A2(new_n722), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n728), .B1(new_n528), .B2(new_n536), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n586), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n579), .A2(new_n728), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n732), .A2(new_n737), .ZN(G399));
  INV_X1    g0538(.A(new_n210), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G41), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n617), .A2(G116), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(G1), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(new_n213), .B2(new_n741), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT28), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n678), .A2(new_n683), .A3(new_n633), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n670), .A2(new_n674), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n633), .A2(new_n679), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n585), .B2(new_n578), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n694), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n722), .B1(new_n746), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(KEYINPUT96), .B1(new_n751), .B2(KEYINPUT29), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT96), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT29), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n753), .B(new_n754), .C1(new_n695), .C2(new_n722), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n634), .A2(new_n682), .A3(new_n672), .A4(new_n681), .ZN(new_n756));
  OAI21_X1  g0556(.A(KEYINPUT26), .B1(new_n674), .B2(new_n748), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n756), .A2(new_n633), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n722), .B1(new_n758), .B2(new_n750), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(KEYINPUT29), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n752), .A2(new_n755), .A3(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G330), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n607), .A2(new_n612), .ZN(new_n763));
  AND3_X1   g0563(.A1(new_n763), .A2(new_n526), .A3(new_n551), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n663), .A2(new_n667), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n764), .A2(new_n765), .A3(KEYINPUT30), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n763), .A2(G179), .A3(new_n499), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(new_n671), .A3(new_n581), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT30), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n763), .A2(new_n526), .A3(new_n551), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n769), .B1(new_n770), .B2(new_n671), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n766), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  AND3_X1   g0572(.A1(new_n772), .A2(KEYINPUT31), .A3(new_n722), .ZN(new_n773));
  AOI21_X1  g0573(.A(KEYINPUT31), .B1(new_n772), .B2(new_n722), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n541), .A2(new_n586), .A3(new_n675), .A4(new_n728), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n762), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n761), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n745), .B1(new_n780), .B2(G1), .ZN(G364));
  INV_X1    g0581(.A(new_n727), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n272), .A2(G20), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n206), .B1(new_n783), .B2(G45), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n740), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(G330), .B2(new_n726), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n210), .A2(new_n327), .ZN(new_n789));
  INV_X1    g0589(.A(G355), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n790), .B1(G116), .B2(new_n210), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n739), .A2(new_n327), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(new_n293), .B2(new_n214), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n245), .A2(new_n293), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n272), .A2(new_n324), .A3(KEYINPUT97), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT97), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(G13), .B2(G33), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n215), .B1(G20), .B2(new_n312), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n786), .B1(new_n796), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT99), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n207), .A2(new_n369), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G200), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n807), .B1(new_n809), .B2(G190), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n809), .A2(new_n807), .A3(G190), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(KEYINPUT33), .B(G317), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n808), .A2(G190), .A3(new_n425), .ZN(new_n817));
  INV_X1    g0617(.A(G322), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G190), .A2(G200), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n808), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n332), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n207), .A2(G179), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n820), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n819), .B(new_n823), .C1(G329), .C2(new_n826), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n423), .A2(G179), .A3(G200), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n207), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n824), .A2(G190), .A3(G200), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n830), .A2(G294), .B1(new_n832), .B2(G303), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n809), .A2(new_n423), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n824), .A2(new_n423), .A3(G200), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n834), .A2(G326), .B1(new_n836), .B2(G283), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n816), .A2(new_n827), .A3(new_n833), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n814), .A2(G68), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n817), .A2(new_n225), .B1(new_n821), .B2(new_n261), .ZN(new_n840));
  INV_X1    g0640(.A(G159), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n825), .A2(KEYINPUT32), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT32), .B1(new_n825), .B2(new_n841), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G97), .A2(new_n830), .B1(new_n834), .B2(G50), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n839), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n832), .A2(G87), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n847), .B(new_n327), .C1(new_n334), .C2(new_n835), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT98), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n838), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n806), .B1(new_n850), .B2(new_n803), .ZN(new_n851));
  INV_X1    g0651(.A(new_n802), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n726), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n788), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G396));
  NAND2_X1  g0655(.A1(new_n363), .A2(new_n722), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n364), .A2(KEYINPUT71), .B1(new_n369), .B2(new_n368), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(new_n367), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n483), .A2(new_n371), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n858), .B1(new_n859), .B2(new_n856), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n751), .ZN(new_n861));
  INV_X1    g0661(.A(new_n856), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n483), .B2(new_n371), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT101), .B1(new_n863), .B2(new_n858), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT101), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n371), .A2(new_n862), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n857), .A2(new_n367), .B1(new_n480), .B2(new_n482), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n865), .B(new_n866), .C1(new_n867), .C2(new_n862), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n861), .B1(new_n869), .B2(new_n751), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n786), .B1(new_n870), .B2(new_n778), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n778), .B2(new_n870), .ZN(new_n872));
  INV_X1    g0672(.A(new_n817), .ZN(new_n873));
  INV_X1    g0673(.A(new_n821), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n873), .A2(G143), .B1(new_n874), .B2(G159), .ZN(new_n875));
  INV_X1    g0675(.A(G137), .ZN(new_n876));
  INV_X1    g0676(.A(new_n834), .ZN(new_n877));
  INV_X1    g0677(.A(G150), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n875), .B1(new_n876), .B2(new_n877), .C1(new_n813), .C2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT34), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n836), .A2(G68), .ZN(new_n883));
  INV_X1    g0683(.A(G132), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n883), .B(new_n327), .C1(new_n884), .C2(new_n825), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n829), .A2(new_n225), .B1(new_n831), .B2(new_n202), .ZN(new_n886));
  NOR4_X1   g0686(.A1(new_n881), .A2(new_n882), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n327), .B1(new_n826), .B2(G311), .ZN(new_n888));
  INV_X1    g0688(.A(G294), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n888), .B1(new_n507), .B2(new_n821), .C1(new_n889), .C2(new_n817), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n832), .A2(G107), .B1(new_n836), .B2(G87), .ZN(new_n891));
  OAI221_X1 g0691(.A(new_n891), .B1(new_n227), .B2(new_n829), .C1(new_n486), .C2(new_n877), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n813), .A2(KEYINPUT100), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n813), .A2(KEYINPUT100), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n890), .B(new_n892), .C1(new_n897), .C2(G283), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n803), .B1(new_n887), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n786), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n800), .A2(new_n803), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n900), .B1(new_n261), .B2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n899), .B(new_n902), .C1(new_n860), .C2(new_n801), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n872), .A2(new_n903), .ZN(G384));
  INV_X1    g0704(.A(new_n641), .ZN(new_n905));
  OAI211_X1 g0705(.A(G116), .B(new_n216), .C1(new_n905), .C2(KEYINPUT35), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n906), .A2(KEYINPUT102), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(KEYINPUT35), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(KEYINPUT102), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT36), .Z(new_n911));
  OAI211_X1 g0711(.A(new_n214), .B(G77), .C1(new_n225), .C2(new_n219), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n202), .A2(G68), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n206), .B(G13), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n775), .A2(new_n776), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n276), .A2(new_n728), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n702), .A2(new_n319), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n917), .B1(new_n700), .B2(new_n320), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(KEYINPUT103), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT103), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n702), .A2(new_n922), .A3(new_n319), .A4(new_n918), .ZN(new_n923));
  AND4_X1   g0723(.A1(new_n916), .A2(new_n860), .A3(new_n921), .A4(new_n923), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n706), .A2(new_n418), .A3(new_n420), .A4(new_n707), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n390), .A2(new_n395), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n438), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n251), .A3(new_n396), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n720), .B1(new_n928), .B2(new_n375), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n398), .B1(new_n430), .B2(new_n434), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n408), .A2(new_n414), .A3(new_n411), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n414), .B1(new_n408), .B2(new_n411), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n934), .A2(new_n720), .B1(new_n375), .B2(new_n928), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT37), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT37), .ZN(new_n937));
  INV_X1    g0737(.A(new_n720), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n398), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n704), .A2(new_n937), .A3(new_n417), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n930), .A2(KEYINPUT38), .A3(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n939), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n704), .A2(new_n417), .A3(new_n939), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT37), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n925), .A2(new_n943), .B1(new_n945), .B2(new_n940), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n942), .B1(KEYINPUT38), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n924), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT38), .ZN(new_n949));
  INV_X1    g0749(.A(new_n929), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n444), .B2(new_n421), .ZN(new_n951));
  INV_X1    g0751(.A(new_n941), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT40), .B1(new_n953), .B2(new_n942), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n948), .A2(KEYINPUT40), .B1(new_n924), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n485), .A2(new_n916), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n958), .A2(new_n959), .A3(new_n762), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n752), .A2(new_n755), .A3(new_n485), .A4(new_n760), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n715), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT39), .ZN(new_n963));
  AOI221_X4 g0763(.A(new_n949), .B1(new_n936), .B2(new_n940), .C1(new_n925), .C2(new_n929), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n925), .A2(new_n943), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n945), .A2(new_n940), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT38), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n963), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n702), .A2(new_n722), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n953), .A2(KEYINPUT39), .A3(new_n942), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n371), .A2(new_n722), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n861), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n953), .A2(new_n942), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n920), .A2(KEYINPUT103), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n316), .A2(new_n320), .A3(new_n917), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n923), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n974), .A2(new_n975), .A3(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n421), .A2(new_n938), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n971), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n962), .B(new_n983), .Z(new_n984));
  OAI22_X1  g0784(.A1(new_n960), .A2(new_n984), .B1(new_n206), .B2(new_n783), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n960), .A2(new_n984), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n915), .B1(new_n985), .B2(new_n986), .ZN(G367));
  XNOR2_X1  g0787(.A(new_n784), .B(KEYINPUT106), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n651), .A2(new_n722), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n747), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n681), .A2(new_n672), .A3(new_n722), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n737), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT44), .Z(new_n994));
  NOR2_X1   g0794(.A1(new_n737), .A2(new_n992), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT45), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n732), .ZN(new_n998));
  INV_X1    g0798(.A(new_n732), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n994), .A2(new_n999), .A3(new_n996), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT105), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n731), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n735), .B1(new_n1003), .B2(new_n734), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(new_n782), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n780), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1001), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1005), .A2(KEYINPUT105), .A3(new_n780), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n779), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n740), .B(KEYINPUT41), .Z(new_n1010));
  OAI21_X1  g0810(.A(new_n988), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n728), .A2(new_n624), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n633), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n680), .B2(new_n1012), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT104), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT43), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n992), .A2(new_n735), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1018), .A2(KEYINPUT42), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n747), .A2(new_n579), .A3(new_n989), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n722), .B1(new_n1020), .B2(new_n674), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n1018), .B2(KEYINPUT42), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1017), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n999), .A2(new_n992), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1011), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n836), .A2(G97), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n877), .B2(new_n822), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n338), .B2(new_n830), .ZN(new_n1031));
  AND3_X1   g0831(.A1(new_n832), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1032));
  AOI21_X1  g0832(.A(KEYINPUT46), .B1(new_n832), .B2(G116), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n332), .B1(new_n817), .B2(new_n486), .ZN(new_n1034));
  INV_X1    g0834(.A(G283), .ZN(new_n1035));
  INV_X1    g0835(.A(G317), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n821), .A2(new_n1035), .B1(new_n825), .B2(new_n1036), .ZN(new_n1037));
  NOR4_X1   g0837(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .A4(new_n1037), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1031), .B(new_n1038), .C1(new_n896), .C2(new_n889), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n829), .A2(new_n219), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G58), .B2(new_n832), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n836), .A2(G77), .ZN(new_n1042));
  INV_X1    g0842(.A(G143), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1041), .B(new_n1042), .C1(new_n1043), .C2(new_n877), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n327), .B1(new_n817), .B2(new_n878), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n821), .A2(new_n202), .B1(new_n825), .B2(new_n876), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n896), .B2(new_n841), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1039), .A2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT47), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n803), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1015), .A2(new_n802), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n359), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n805), .B1(new_n739), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n792), .A2(new_n241), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n900), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AND3_X1   g0856(.A1(new_n1051), .A2(new_n1052), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1028), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(G387));
  INV_X1    g0859(.A(new_n988), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1005), .A2(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n789), .A2(new_n742), .B1(G107), .B2(new_n210), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n238), .A2(G45), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n742), .B(KEYINPUT107), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n202), .B2(new_n357), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n356), .A2(new_n1065), .A3(G50), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n293), .B1(new_n219), .B2(new_n261), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n793), .B1(new_n1064), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1062), .B1(new_n1063), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n786), .B1(new_n1072), .B2(new_n805), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT109), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n830), .A2(new_n1053), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n834), .A2(G159), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n832), .A2(G77), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1075), .A2(new_n1076), .A3(new_n1029), .A4(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n332), .B1(new_n826), .B2(G150), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(new_n202), .B2(new_n817), .C1(new_n219), .C2(new_n821), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(new_n357), .C2(new_n814), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n835), .A2(new_n507), .ZN(new_n1082));
  INV_X1    g0882(.A(G326), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n332), .B1(new_n825), .B2(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n873), .A2(G317), .B1(new_n874), .B2(G303), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n818), .B2(new_n877), .C1(new_n896), .C2(new_n822), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT48), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n829), .A2(new_n1035), .B1(new_n831), .B2(new_n889), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT110), .Z(new_n1091));
  NAND3_X1  g0891(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1082), .B(new_n1084), .C1(new_n1093), .C2(KEYINPUT49), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1093), .A2(KEYINPUT49), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1081), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n803), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1074), .B1(new_n1003), .B2(new_n852), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1006), .A2(new_n740), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1005), .A2(new_n780), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1061), .B(new_n1098), .C1(new_n1099), .C2(new_n1100), .ZN(G393));
  NAND2_X1  g0901(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n741), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT111), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n988), .B1(new_n1001), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n998), .A2(KEYINPUT111), .A3(new_n1000), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n992), .A2(new_n802), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n877), .A2(new_n1036), .B1(new_n822), .B2(new_n817), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT52), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n334), .A2(new_n835), .B1(new_n831), .B2(new_n1035), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n332), .B1(new_n825), .B2(new_n818), .C1(new_n889), .C2(new_n821), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1111), .B(new_n1112), .C1(G116), .C2(new_n830), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1110), .B(new_n1113), .C1(new_n896), .C2(new_n486), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n327), .B1(new_n825), .B2(new_n1043), .C1(new_n356), .C2(new_n821), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n830), .A2(G77), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n221), .B2(new_n835), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1115), .B(new_n1117), .C1(G68), .C2(new_n832), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n877), .A2(new_n878), .B1(new_n841), .B2(new_n817), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT51), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1118), .B(new_n1120), .C1(new_n896), .C2(new_n202), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1097), .B1(new_n1114), .B2(new_n1121), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n793), .A2(new_n248), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n805), .B1(G97), .B2(new_n739), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n900), .B(new_n1122), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1106), .A2(new_n1107), .B1(new_n1108), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1104), .A2(new_n1126), .ZN(G390));
  NAND2_X1  g0927(.A1(new_n968), .A2(new_n970), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n969), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n972), .B1(new_n860), .B2(new_n751), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1129), .B1(new_n1130), .B2(new_n978), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n866), .B1(new_n867), .B2(new_n862), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n978), .A2(new_n1133), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1134), .A2(KEYINPUT112), .A3(new_n777), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n972), .B1(new_n759), .B2(new_n860), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1129), .B(new_n947), .C1(new_n1136), .C2(new_n978), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1132), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1135), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1060), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT54), .B(G143), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n897), .A2(G137), .B1(new_n874), .B2(new_n1142), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1143), .A2(KEYINPUT114), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(KEYINPUT114), .ZN(new_n1145));
  INV_X1    g0945(.A(G128), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n877), .A2(new_n1146), .B1(new_n835), .B2(new_n202), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G159), .B2(new_n830), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n831), .A2(new_n878), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT53), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n817), .A2(new_n884), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n332), .B(new_n1151), .C1(G125), .C2(new_n826), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1148), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n1144), .A2(new_n1145), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT115), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n834), .A2(G283), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1116), .A2(new_n1157), .A3(new_n847), .A4(new_n883), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n332), .B1(new_n817), .B2(new_n507), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n821), .A2(new_n227), .B1(new_n825), .B2(new_n889), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n896), .B2(new_n350), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1156), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1155), .A2(KEYINPUT115), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n803), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1128), .A2(new_n800), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n900), .B1(new_n356), .B2(new_n901), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1140), .A2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n485), .A2(new_n777), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n961), .A2(new_n473), .A3(new_n714), .A4(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(KEYINPUT113), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT113), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n715), .A2(new_n1174), .A3(new_n961), .A4(new_n1171), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n916), .A2(new_n860), .A3(G330), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n777), .A2(new_n1134), .B1(new_n1176), .B2(new_n978), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n979), .B1(new_n869), .B2(new_n777), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n860), .A2(new_n921), .A3(new_n923), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1136), .B1(new_n778), .B2(new_n1179), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n1177), .A2(new_n1130), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1173), .A2(new_n1175), .A3(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1170), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n741), .B1(new_n1170), .B2(new_n1182), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1169), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(G378));
  NAND2_X1  g0986(.A1(new_n713), .A2(new_n473), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n453), .A2(new_n720), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT117), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n964), .A2(new_n967), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n916), .A2(new_n860), .A3(new_n921), .A4(new_n923), .ZN(new_n1198));
  OAI21_X1  g0998(.A(KEYINPUT40), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n924), .A2(new_n954), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n762), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1201), .A2(new_n983), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n983), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1196), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n980), .A2(new_n982), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n971), .B(new_n1205), .C1(new_n955), .C2(new_n762), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1201), .A2(new_n983), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n1195), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n988), .B1(new_n1204), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n901), .A2(new_n202), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n786), .A2(new_n1210), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1192), .A2(new_n1193), .A3(new_n801), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n877), .A2(new_n507), .B1(new_n835), .B2(new_n225), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1040), .B(new_n1213), .C1(G77), .C2(new_n832), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n332), .A2(new_n292), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n817), .A2(new_n334), .B1(new_n821), .B2(new_n359), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(G283), .C2(new_n826), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1214), .B(new_n1217), .C1(new_n227), .C2(new_n813), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT58), .ZN(new_n1219));
  AOI21_X1  g1019(.A(G50), .B1(new_n324), .B2(new_n292), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1218), .A2(new_n1219), .B1(new_n1215), .B2(new_n1220), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n817), .A2(new_n1146), .B1(new_n821), .B2(new_n876), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G150), .B2(new_n830), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n834), .A2(G125), .B1(new_n832), .B2(new_n1142), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n813), .C2(new_n884), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1227));
  OR2_X1    g1027(.A1(KEYINPUT116), .A2(G124), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(KEYINPUT116), .A2(G124), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n826), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1230), .A2(new_n324), .A3(new_n292), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1227), .B(new_n1231), .C1(new_n841), .C2(new_n835), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1221), .B1(new_n1219), .B2(new_n1218), .C1(new_n1226), .C2(new_n1232), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1211), .B(new_n1212), .C1(new_n803), .C2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1209), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1204), .A2(new_n1208), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1181), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1238), .B1(new_n1170), .B2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1236), .A2(KEYINPUT57), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n740), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT57), .B1(new_n1236), .B2(new_n1240), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1235), .B1(new_n1242), .B2(new_n1243), .ZN(G375));
  AOI21_X1  g1044(.A(new_n900), .B1(new_n219), .B2(new_n901), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n830), .A2(G50), .B1(new_n832), .B2(G159), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n834), .A2(G132), .B1(new_n836), .B2(G58), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n332), .B1(new_n873), .B2(G137), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G150), .A2(new_n874), .B1(new_n826), .B2(G128), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n897), .B2(new_n1142), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n332), .B1(new_n825), .B2(new_n486), .C1(new_n817), .C2(new_n1035), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n834), .A2(G294), .B1(new_n832), .B2(G97), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1253), .A2(new_n1042), .A3(new_n1075), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n897), .A2(G116), .B1(new_n338), .B2(new_n874), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1252), .B(new_n1254), .C1(new_n1256), .C2(KEYINPUT118), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1256), .A2(KEYINPUT118), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1251), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1245), .B1(new_n1259), .B2(new_n1097), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n978), .B2(new_n800), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n1181), .B2(new_n1060), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1010), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1182), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1181), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1262), .B1(new_n1264), .B2(new_n1265), .ZN(G381));
  XOR2_X1   g1066(.A(G375), .B(KEYINPUT119), .Z(new_n1267));
  OR2_X1    g1067(.A1(G393), .A2(G396), .ZN(new_n1268));
  NOR4_X1   g1068(.A1(G390), .A2(G384), .A3(new_n1268), .A4(G381), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1058), .A2(new_n1185), .A3(new_n1269), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1267), .A2(new_n1270), .ZN(G407));
  NAND2_X1  g1071(.A1(new_n721), .A2(G213), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1185), .A2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G407), .B(G213), .C1(new_n1267), .C2(new_n1274), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(KEYINPUT120), .ZN(G409));
  NAND3_X1  g1076(.A1(new_n1237), .A2(KEYINPUT60), .A3(new_n1239), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n740), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1265), .B1(KEYINPUT60), .B2(new_n1182), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1262), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(G384), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G384), .B(new_n1262), .C1(new_n1278), .C2(new_n1279), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G378), .B(new_n1235), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1209), .A2(new_n1234), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1236), .A2(new_n1263), .A3(new_n1240), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1185), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1273), .B(new_n1284), .C1(new_n1285), .C2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(KEYINPUT124), .B1(new_n1289), .B2(KEYINPUT62), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1284), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1291), .A2(KEYINPUT62), .A3(new_n1272), .A4(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT125), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1273), .B1(new_n1285), .B2(new_n1288), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1296), .A2(KEYINPUT125), .A3(KEYINPUT62), .A4(new_n1292), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1291), .A2(new_n1272), .A3(new_n1292), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT124), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT62), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1290), .A2(new_n1295), .A3(new_n1297), .A4(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT61), .ZN(new_n1303));
  OR2_X1    g1103(.A1(new_n1272), .A2(KEYINPUT121), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1282), .A2(new_n1283), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1273), .A2(G2897), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1282), .A2(new_n1306), .A3(new_n1283), .A4(new_n1304), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1303), .B1(new_n1310), .B2(new_n1296), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(KEYINPUT123), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT123), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1313), .B(new_n1303), .C1(new_n1310), .C2(new_n1296), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1302), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(KEYINPUT126), .ZN(new_n1317));
  OR2_X1    g1117(.A1(new_n1058), .A2(G390), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT122), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1058), .A2(G390), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(G393), .B(new_n854), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1318), .A2(new_n1319), .A3(new_n1320), .A4(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1319), .B1(new_n1058), .B2(G390), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  AOI22_X1  g1126(.A1(new_n1326), .A2(new_n1322), .B1(new_n1318), .B2(new_n1320), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1324), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT126), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1302), .A2(new_n1315), .A3(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1317), .A2(new_n1328), .A3(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1311), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1298), .B(KEYINPUT63), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1332), .B(new_n1333), .C1(new_n1324), .C2(new_n1327), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1331), .A2(new_n1334), .ZN(G405));
  XNOR2_X1  g1135(.A(G375), .B(G378), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1292), .A2(KEYINPUT127), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1320), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1058), .A2(G390), .ZN(new_n1340));
  OAI22_X1  g1140(.A1(new_n1339), .A2(new_n1340), .B1(new_n1325), .B2(new_n1321), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1292), .A2(KEYINPUT127), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1341), .A2(new_n1323), .A3(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1343), .B1(new_n1341), .B2(new_n1323), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1338), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1342), .B1(new_n1324), .B2(new_n1327), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1338), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1348), .A2(new_n1349), .A3(new_n1344), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1347), .A2(new_n1350), .ZN(G402));
endmodule


