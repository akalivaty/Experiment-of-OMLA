

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577;

  XOR2_X1 U322 ( .A(n469), .B(KEYINPUT28), .Z(n524) );
  XNOR2_X1 U323 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U324 ( .A(n405), .B(n313), .Z(n510) );
  XOR2_X1 U325 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n290) );
  XOR2_X1 U326 ( .A(KEYINPUT94), .B(n301), .Z(n291) );
  XOR2_X1 U327 ( .A(n303), .B(KEYINPUT95), .Z(n292) );
  AND2_X1 U328 ( .A1(G227GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U329 ( .A(n311), .B(n310), .Z(n294) );
  XNOR2_X1 U330 ( .A(KEYINPUT25), .B(KEYINPUT101), .ZN(n413) );
  XNOR2_X1 U331 ( .A(n414), .B(n413), .ZN(n418) );
  INV_X1 U332 ( .A(KEYINPUT48), .ZN(n463) );
  XNOR2_X1 U333 ( .A(n383), .B(n349), .ZN(n350) );
  XNOR2_X1 U334 ( .A(n463), .B(KEYINPUT114), .ZN(n464) );
  XNOR2_X1 U335 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U336 ( .A(n465), .B(n464), .ZN(n519) );
  INV_X1 U337 ( .A(G78GAT), .ZN(n357) );
  XNOR2_X1 U338 ( .A(n374), .B(n293), .ZN(n375) );
  NOR2_X1 U339 ( .A1(n426), .A2(n425), .ZN(n427) );
  XNOR2_X1 U340 ( .A(n358), .B(n357), .ZN(n359) );
  NOR2_X1 U341 ( .A1(n447), .A2(n575), .ZN(n448) );
  XNOR2_X1 U342 ( .A(KEYINPUT103), .B(n427), .ZN(n478) );
  XNOR2_X1 U343 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U344 ( .A(n392), .B(n379), .ZN(n522) );
  XNOR2_X1 U345 ( .A(n449), .B(KEYINPUT38), .ZN(n494) );
  XNOR2_X1 U346 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U347 ( .A(n450), .B(G29GAT), .ZN(n451) );
  XNOR2_X1 U348 ( .A(n475), .B(n474), .ZN(G1351GAT) );
  XNOR2_X1 U349 ( .A(n452), .B(n451), .ZN(G1328GAT) );
  XOR2_X1 U350 ( .A(KEYINPUT2), .B(KEYINPUT91), .Z(n296) );
  XNOR2_X1 U351 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n295) );
  XNOR2_X1 U352 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U353 ( .A(n297), .B(G162GAT), .Z(n299) );
  XNOR2_X1 U354 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n405) );
  XNOR2_X1 U356 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n290), .B(n300), .ZN(n301) );
  NAND2_X1 U358 ( .A1(G225GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n291), .B(n302), .ZN(n303) );
  XOR2_X1 U360 ( .A(G120GAT), .B(KEYINPUT82), .Z(n305) );
  XNOR2_X1 U361 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U363 ( .A(KEYINPUT81), .B(n306), .Z(n376) );
  XNOR2_X1 U364 ( .A(n376), .B(G57GAT), .ZN(n307) );
  XNOR2_X1 U365 ( .A(n292), .B(n307), .ZN(n311) );
  XOR2_X1 U366 ( .A(G127GAT), .B(G155GAT), .Z(n356) );
  XOR2_X1 U367 ( .A(G148GAT), .B(n356), .Z(n309) );
  XOR2_X1 U368 ( .A(G134GAT), .B(KEYINPUT76), .Z(n438) );
  XNOR2_X1 U369 ( .A(G1GAT), .B(n438), .ZN(n308) );
  XNOR2_X1 U370 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U371 ( .A(G29GAT), .B(G85GAT), .ZN(n312) );
  XNOR2_X1 U372 ( .A(n294), .B(n312), .ZN(n313) );
  XNOR2_X1 U373 ( .A(G169GAT), .B(G36GAT), .ZN(n314) );
  XNOR2_X1 U374 ( .A(n314), .B(G8GAT), .ZN(n380) );
  XOR2_X1 U375 ( .A(G197GAT), .B(n380), .Z(n316) );
  NAND2_X1 U376 ( .A1(G229GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U378 ( .A(n317), .B(KEYINPUT65), .Z(n327) );
  XOR2_X1 U379 ( .A(G50GAT), .B(G29GAT), .Z(n319) );
  XNOR2_X1 U380 ( .A(KEYINPUT67), .B(KEYINPUT7), .ZN(n318) );
  XNOR2_X1 U381 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U382 ( .A(n320), .B(KEYINPUT8), .Z(n322) );
  XNOR2_X1 U383 ( .A(G43GAT), .B(KEYINPUT68), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n322), .B(n321), .ZN(n444) );
  XOR2_X1 U385 ( .A(KEYINPUT70), .B(KEYINPUT29), .Z(n324) );
  XNOR2_X1 U386 ( .A(G141GAT), .B(G113GAT), .ZN(n323) );
  XNOR2_X1 U387 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U388 ( .A(n444), .B(n325), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U390 ( .A(n328), .B(KEYINPUT30), .Z(n332) );
  XOR2_X1 U391 ( .A(G1GAT), .B(G15GAT), .Z(n330) );
  XNOR2_X1 U392 ( .A(KEYINPUT69), .B(G22GAT), .ZN(n329) );
  XNOR2_X1 U393 ( .A(n330), .B(n329), .ZN(n353) );
  XNOR2_X1 U394 ( .A(n353), .B(KEYINPUT66), .ZN(n331) );
  XNOR2_X1 U395 ( .A(n332), .B(n331), .ZN(n563) );
  XNOR2_X1 U396 ( .A(n563), .B(KEYINPUT71), .ZN(n551) );
  XOR2_X1 U397 ( .A(KEYINPUT72), .B(KEYINPUT13), .Z(n334) );
  XNOR2_X1 U398 ( .A(G71GAT), .B(G57GAT), .ZN(n333) );
  XNOR2_X1 U399 ( .A(n334), .B(n333), .ZN(n351) );
  XOR2_X1 U400 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n336) );
  NAND2_X1 U401 ( .A1(G230GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U402 ( .A(n336), .B(n335), .ZN(n339) );
  XOR2_X1 U403 ( .A(G64GAT), .B(G204GAT), .Z(n338) );
  XNOR2_X1 U404 ( .A(G176GAT), .B(G92GAT), .ZN(n337) );
  XNOR2_X1 U405 ( .A(n338), .B(n337), .ZN(n389) );
  XOR2_X1 U406 ( .A(n339), .B(n389), .Z(n342) );
  XNOR2_X1 U407 ( .A(G148GAT), .B(G106GAT), .ZN(n340) );
  XNOR2_X1 U408 ( .A(n340), .B(G78GAT), .ZN(n404) );
  XNOR2_X1 U409 ( .A(G120GAT), .B(n404), .ZN(n341) );
  XNOR2_X1 U410 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U411 ( .A(n343), .B(KEYINPUT31), .Z(n345) );
  XOR2_X1 U412 ( .A(G99GAT), .B(G85GAT), .Z(n434) );
  XNOR2_X1 U413 ( .A(n434), .B(KEYINPUT32), .ZN(n344) );
  XNOR2_X1 U414 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U415 ( .A(n351), .B(n346), .ZN(n453) );
  NAND2_X1 U416 ( .A1(n551), .A2(n453), .ZN(n480) );
  XOR2_X1 U417 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n348) );
  XNOR2_X1 U418 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n347) );
  XNOR2_X1 U419 ( .A(n348), .B(n347), .ZN(n362) );
  XOR2_X1 U420 ( .A(G183GAT), .B(G211GAT), .Z(n383) );
  AND2_X1 U421 ( .A1(G231GAT), .A2(G233GAT), .ZN(n349) );
  XOR2_X1 U422 ( .A(n352), .B(KEYINPUT78), .Z(n355) );
  XNOR2_X1 U423 ( .A(n353), .B(KEYINPUT12), .ZN(n354) );
  XNOR2_X1 U424 ( .A(n355), .B(n354), .ZN(n360) );
  XNOR2_X1 U425 ( .A(G8GAT), .B(n356), .ZN(n358) );
  XNOR2_X1 U426 ( .A(n362), .B(n361), .ZN(n571) );
  XOR2_X1 U427 ( .A(KEYINPUT17), .B(G190GAT), .Z(n364) );
  XNOR2_X1 U428 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n363) );
  XNOR2_X1 U429 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U430 ( .A(KEYINPUT83), .B(n365), .Z(n392) );
  XOR2_X1 U431 ( .A(KEYINPUT84), .B(G127GAT), .Z(n367) );
  XNOR2_X1 U432 ( .A(G71GAT), .B(G183GAT), .ZN(n366) );
  XNOR2_X1 U433 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U434 ( .A(G176GAT), .B(G15GAT), .Z(n369) );
  XNOR2_X1 U435 ( .A(G169GAT), .B(G43GAT), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U437 ( .A(n371), .B(n370), .ZN(n378) );
  XOR2_X1 U438 ( .A(G99GAT), .B(G134GAT), .Z(n373) );
  XNOR2_X1 U439 ( .A(KEYINPUT85), .B(KEYINPUT20), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U442 ( .A(n380), .B(KEYINPUT97), .Z(n382) );
  NAND2_X1 U443 ( .A1(G226GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n382), .B(n381), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n383), .B(KEYINPUT96), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n384), .B(KEYINPUT98), .ZN(n385) );
  XOR2_X1 U447 ( .A(n386), .B(n385), .Z(n391) );
  XOR2_X1 U448 ( .A(KEYINPUT88), .B(KEYINPUT21), .Z(n388) );
  XNOR2_X1 U449 ( .A(G197GAT), .B(G218GAT), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n389), .B(n394), .ZN(n390) );
  XOR2_X1 U452 ( .A(n391), .B(n390), .Z(n393) );
  XNOR2_X1 U453 ( .A(n393), .B(n392), .ZN(n512) );
  NAND2_X1 U454 ( .A1(n522), .A2(n512), .ZN(n412) );
  XOR2_X1 U455 ( .A(n394), .B(G22GAT), .Z(n396) );
  NAND2_X1 U456 ( .A1(G228GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U457 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U458 ( .A(G50GAT), .B(n397), .ZN(n411) );
  XOR2_X1 U459 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n399) );
  XNOR2_X1 U460 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n398) );
  XNOR2_X1 U461 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U462 ( .A(KEYINPUT86), .B(G211GAT), .Z(n401) );
  XNOR2_X1 U463 ( .A(G155GAT), .B(G204GAT), .ZN(n400) );
  XNOR2_X1 U464 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n403), .B(n402), .ZN(n409) );
  XOR2_X1 U466 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n407) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n469) );
  NAND2_X1 U471 ( .A1(n412), .A2(n469), .ZN(n414) );
  NOR2_X1 U472 ( .A1(n469), .A2(n522), .ZN(n416) );
  XNOR2_X1 U473 ( .A(KEYINPUT26), .B(KEYINPUT100), .ZN(n415) );
  XNOR2_X1 U474 ( .A(n416), .B(n415), .ZN(n561) );
  XNOR2_X1 U475 ( .A(n512), .B(KEYINPUT27), .ZN(n421) );
  NAND2_X1 U476 ( .A1(n561), .A2(n421), .ZN(n417) );
  NAND2_X1 U477 ( .A1(n418), .A2(n417), .ZN(n419) );
  XOR2_X1 U478 ( .A(KEYINPUT102), .B(n419), .Z(n420) );
  NOR2_X1 U479 ( .A1(n510), .A2(n420), .ZN(n426) );
  NAND2_X1 U480 ( .A1(n421), .A2(n510), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n422), .B(KEYINPUT99), .ZN(n520) );
  INV_X1 U482 ( .A(n524), .ZN(n423) );
  NAND2_X1 U483 ( .A1(n520), .A2(n423), .ZN(n424) );
  NOR2_X1 U484 ( .A1(n424), .A2(n522), .ZN(n425) );
  NAND2_X1 U485 ( .A1(n571), .A2(n478), .ZN(n447) );
  XOR2_X1 U486 ( .A(KEYINPUT10), .B(KEYINPUT75), .Z(n429) );
  XNOR2_X1 U487 ( .A(G218GAT), .B(KEYINPUT64), .ZN(n428) );
  XNOR2_X1 U488 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U489 ( .A(G92GAT), .B(G162GAT), .Z(n431) );
  XNOR2_X1 U490 ( .A(G36GAT), .B(G190GAT), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U492 ( .A(n433), .B(n432), .Z(n440) );
  XOR2_X1 U493 ( .A(n434), .B(G106GAT), .Z(n436) );
  NAND2_X1 U494 ( .A1(G232GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U497 ( .A(n440), .B(n439), .ZN(n446) );
  XOR2_X1 U498 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n442) );
  XNOR2_X1 U499 ( .A(KEYINPUT9), .B(KEYINPUT77), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U501 ( .A(n444), .B(n443), .Z(n445) );
  XOR2_X1 U502 ( .A(n446), .B(n445), .Z(n534) );
  XOR2_X1 U503 ( .A(KEYINPUT36), .B(n534), .Z(n575) );
  XNOR2_X1 U504 ( .A(n448), .B(KEYINPUT37), .ZN(n508) );
  NOR2_X1 U505 ( .A1(n480), .A2(n508), .ZN(n449) );
  NAND2_X1 U506 ( .A1(n510), .A2(n494), .ZN(n452) );
  XOR2_X1 U507 ( .A(KEYINPUT106), .B(KEYINPUT39), .Z(n450) );
  INV_X1 U508 ( .A(n534), .ZN(n548) );
  XNOR2_X1 U509 ( .A(KEYINPUT113), .B(n571), .ZN(n530) );
  XOR2_X1 U510 ( .A(n453), .B(KEYINPUT41), .Z(n553) );
  NOR2_X1 U511 ( .A1(n563), .A2(n553), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n454), .B(KEYINPUT46), .ZN(n455) );
  NOR2_X1 U513 ( .A1(n530), .A2(n455), .ZN(n456) );
  NAND2_X1 U514 ( .A1(n456), .A2(n548), .ZN(n457) );
  XNOR2_X1 U515 ( .A(n457), .B(KEYINPUT47), .ZN(n462) );
  NOR2_X1 U516 ( .A1(n575), .A2(n571), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n458), .B(KEYINPUT45), .ZN(n459) );
  NAND2_X1 U518 ( .A1(n459), .A2(n453), .ZN(n460) );
  NOR2_X1 U519 ( .A1(n551), .A2(n460), .ZN(n461) );
  NOR2_X1 U520 ( .A1(n462), .A2(n461), .ZN(n465) );
  XNOR2_X1 U521 ( .A(KEYINPUT122), .B(n512), .ZN(n466) );
  AND2_X1 U522 ( .A1(n519), .A2(n466), .ZN(n467) );
  XOR2_X1 U523 ( .A(KEYINPUT54), .B(n467), .Z(n468) );
  NOR2_X1 U524 ( .A1(n510), .A2(n468), .ZN(n562) );
  NAND2_X1 U525 ( .A1(n562), .A2(n469), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n470), .B(KEYINPUT55), .ZN(n471) );
  NAND2_X1 U527 ( .A1(n471), .A2(n522), .ZN(n554) );
  NOR2_X1 U528 ( .A1(n548), .A2(n554), .ZN(n475) );
  XNOR2_X1 U529 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n473) );
  INV_X1 U530 ( .A(G190GAT), .ZN(n472) );
  NOR2_X1 U531 ( .A1(n534), .A2(n571), .ZN(n477) );
  XNOR2_X1 U532 ( .A(KEYINPUT16), .B(KEYINPUT80), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n477), .B(n476), .ZN(n479) );
  NAND2_X1 U534 ( .A1(n479), .A2(n478), .ZN(n498) );
  NOR2_X1 U535 ( .A1(n480), .A2(n498), .ZN(n487) );
  NAND2_X1 U536 ( .A1(n487), .A2(n510), .ZN(n481) );
  XNOR2_X1 U537 ( .A(n481), .B(KEYINPUT34), .ZN(n482) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(n482), .ZN(G1324GAT) );
  NAND2_X1 U539 ( .A1(n487), .A2(n512), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n483), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n485) );
  NAND2_X1 U542 ( .A1(n487), .A2(n522), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U544 ( .A(G15GAT), .B(n486), .ZN(G1326GAT) );
  XOR2_X1 U545 ( .A(G22GAT), .B(KEYINPUT105), .Z(n489) );
  NAND2_X1 U546 ( .A1(n487), .A2(n524), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(G1327GAT) );
  NAND2_X1 U548 ( .A1(n494), .A2(n512), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n490), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n492) );
  NAND2_X1 U551 ( .A1(n494), .A2(n522), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U553 ( .A(G43GAT), .B(n493), .ZN(G1330GAT) );
  XNOR2_X1 U554 ( .A(G50GAT), .B(KEYINPUT108), .ZN(n496) );
  NAND2_X1 U555 ( .A1(n524), .A2(n494), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(G1331GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n500) );
  INV_X1 U558 ( .A(n553), .ZN(n526) );
  NAND2_X1 U559 ( .A1(n526), .A2(n563), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(KEYINPUT110), .ZN(n509) );
  NOR2_X1 U561 ( .A1(n509), .A2(n498), .ZN(n504) );
  NAND2_X1 U562 ( .A1(n504), .A2(n510), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(n501), .ZN(G1332GAT) );
  NAND2_X1 U565 ( .A1(n504), .A2(n512), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n502), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U567 ( .A1(n522), .A2(n504), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n503), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n506) );
  NAND2_X1 U570 ( .A1(n504), .A2(n524), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U572 ( .A(G78GAT), .B(n507), .Z(G1335GAT) );
  NOR2_X1 U573 ( .A1(n509), .A2(n508), .ZN(n516) );
  NAND2_X1 U574 ( .A1(n510), .A2(n516), .ZN(n511) );
  XNOR2_X1 U575 ( .A(G85GAT), .B(n511), .ZN(G1336GAT) );
  NAND2_X1 U576 ( .A1(n516), .A2(n512), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n513), .B(KEYINPUT112), .ZN(n514) );
  XNOR2_X1 U578 ( .A(G92GAT), .B(n514), .ZN(G1337GAT) );
  NAND2_X1 U579 ( .A1(n522), .A2(n516), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U581 ( .A1(n516), .A2(n524), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(KEYINPUT44), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G106GAT), .B(n518), .ZN(G1339GAT) );
  NAND2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U585 ( .A(KEYINPUT115), .B(n521), .ZN(n538) );
  NAND2_X1 U586 ( .A1(n538), .A2(n522), .ZN(n523) );
  NOR2_X1 U587 ( .A1(n524), .A2(n523), .ZN(n535) );
  NAND2_X1 U588 ( .A1(n551), .A2(n535), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n525), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n528) );
  NAND2_X1 U591 ( .A1(n535), .A2(n526), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U593 ( .A(G120GAT), .B(n529), .ZN(G1341GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n532) );
  NAND2_X1 U595 ( .A1(n535), .A2(n530), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U598 ( .A(G134GAT), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(G1343GAT) );
  NAND2_X1 U601 ( .A1(n561), .A2(n538), .ZN(n539) );
  XNOR2_X1 U602 ( .A(KEYINPUT118), .B(n539), .ZN(n549) );
  NOR2_X1 U603 ( .A1(n549), .A2(n563), .ZN(n542) );
  XNOR2_X1 U604 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n540), .B(KEYINPUT120), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(G1344GAT) );
  NOR2_X1 U607 ( .A1(n553), .A2(n549), .ZN(n546) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n544) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NOR2_X1 U612 ( .A1(n549), .A2(n571), .ZN(n547) );
  XOR2_X1 U613 ( .A(G155GAT), .B(n547), .Z(G1346GAT) );
  NOR2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U615 ( .A(G162GAT), .B(n550), .Z(G1347GAT) );
  INV_X1 U616 ( .A(n554), .ZN(n558) );
  AND2_X1 U617 ( .A1(n551), .A2(n558), .ZN(n552) );
  XOR2_X1 U618 ( .A(G169GAT), .B(n552), .Z(G1348GAT) );
  NOR2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n556) );
  XNOR2_X1 U620 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(n557), .ZN(G1349GAT) );
  XOR2_X1 U623 ( .A(G183GAT), .B(KEYINPUT123), .Z(n560) );
  NAND2_X1 U624 ( .A1(n558), .A2(n530), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1350GAT) );
  NAND2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n574) );
  NOR2_X1 U627 ( .A1(n574), .A2(n563), .ZN(n567) );
  XOR2_X1 U628 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n565) );
  XNOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n567), .B(n566), .ZN(G1352GAT) );
  NOR2_X1 U632 ( .A1(n453), .A2(n574), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT61), .B(KEYINPUT126), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G204GAT), .B(n570), .ZN(G1353GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n574), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1354GAT) );
  NOR2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U640 ( .A(KEYINPUT62), .B(n576), .Z(n577) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(n577), .ZN(G1355GAT) );
endmodule

