//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942;
  XNOR2_X1  g000(.A(KEYINPUT99), .B(G8gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G1gat), .ZN(new_n204));
  AND2_X1   g003(.A1(KEYINPUT97), .A2(G1gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT16), .B1(KEYINPUT97), .B2(G1gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  AOI211_X1 g006(.A(new_n202), .B(new_n204), .C1(KEYINPUT98), .C2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(KEYINPUT98), .B2(new_n207), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(G1gat), .B2(new_n203), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G8gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT100), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(KEYINPUT100), .ZN(new_n214));
  NOR2_X1   g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT14), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G29gat), .A2(G36gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n218), .B(KEYINPUT96), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT15), .ZN(new_n221));
  XNOR2_X1  g020(.A(G43gat), .B(G50gat), .ZN(new_n222));
  NOR3_X1   g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n220), .A2(new_n221), .ZN(new_n224));
  INV_X1    g023(.A(new_n222), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n220), .A2(new_n221), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n223), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT17), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n229), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n213), .B(new_n214), .C1(new_n230), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT101), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n209), .A2(new_n211), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(new_n228), .ZN(new_n237));
  INV_X1    g036(.A(new_n228), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(new_n212), .A3(KEYINPUT101), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n233), .A2(new_n234), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n233), .A2(KEYINPUT18), .A3(new_n240), .A4(new_n234), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n240), .B1(new_n212), .B2(new_n238), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n234), .B(KEYINPUT13), .Z(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G141gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT95), .B(G197gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT11), .B(G169gat), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT12), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n243), .A2(new_n247), .A3(new_n244), .A4(new_n254), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G85gat), .A2(G92gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT7), .ZN(new_n260));
  NAND2_X1  g059(.A1(G99gat), .A2(G106gat), .ZN(new_n261));
  INV_X1    g060(.A(G85gat), .ZN(new_n262));
  INV_X1    g061(.A(G92gat), .ZN(new_n263));
  AOI22_X1  g062(.A1(KEYINPUT8), .A2(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(G99gat), .B(G106gat), .Z(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n267), .B1(new_n232), .B2(new_n230), .ZN(new_n268));
  INV_X1    g067(.A(new_n267), .ZN(new_n269));
  AND2_X1   g068(.A1(G232gat), .A2(G233gat), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n238), .A2(new_n269), .B1(KEYINPUT41), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(G190gat), .B(G218gat), .Z(new_n273));
  XOR2_X1   g072(.A(new_n272), .B(new_n273), .Z(new_n274));
  NOR2_X1   g073(.A1(new_n270), .A2(KEYINPUT41), .ZN(new_n275));
  XNOR2_X1  g074(.A(G134gat), .B(G162gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n274), .A2(new_n277), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT21), .ZN(new_n282));
  XOR2_X1   g081(.A(G71gat), .B(G78gat), .Z(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT9), .ZN(new_n285));
  INV_X1    g084(.A(G71gat), .ZN(new_n286));
  INV_X1    g085(.A(G78gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(G57gat), .B(G64gat), .Z(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n288), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n283), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n236), .B1(new_n282), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT104), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n282), .ZN(new_n296));
  XOR2_X1   g095(.A(KEYINPUT103), .B(KEYINPUT19), .Z(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n295), .B(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G127gat), .B(G155gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(KEYINPUT20), .ZN(new_n301));
  NAND2_X1  g100(.A1(G231gat), .A2(G233gat), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n302), .B(KEYINPUT102), .Z(new_n303));
  XNOR2_X1  g102(.A(new_n301), .B(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G183gat), .B(G211gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n299), .A2(new_n306), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n293), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n265), .A2(KEYINPUT105), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n269), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n267), .A2(new_n310), .A3(new_n311), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT10), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n293), .A2(new_n316), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n315), .A2(new_n316), .B1(new_n269), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(G230gat), .A2(G233gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n313), .A2(new_n319), .A3(new_n314), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G120gat), .B(G148gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(G176gat), .B(G204gat), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n324), .B(new_n325), .Z(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n321), .A2(new_n322), .A3(new_n326), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n281), .A2(new_n309), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT87), .ZN(new_n333));
  XOR2_X1   g132(.A(G155gat), .B(G162gat), .Z(new_n334));
  INV_X1    g133(.A(G141gat), .ZN(new_n335));
  INV_X1    g134(.A(G148gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n334), .B1(KEYINPUT2), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT81), .ZN(new_n342));
  INV_X1    g141(.A(G155gat), .ZN(new_n343));
  INV_X1    g142(.A(G162gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT80), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT80), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G162gat), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n343), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT2), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n342), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT80), .B(G162gat), .ZN(new_n351));
  OAI211_X1 g150(.A(KEYINPUT81), .B(KEYINPUT2), .C1(new_n351), .C2(new_n343), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n334), .A2(new_n339), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT82), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n350), .A2(KEYINPUT82), .A3(new_n352), .A4(new_n353), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n341), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT29), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n361));
  OR2_X1    g160(.A1(G197gat), .A2(G204gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(G197gat), .A2(G204gat), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G211gat), .B(G218gat), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT75), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n365), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n362), .A2(new_n363), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n367), .B(new_n368), .C1(new_n369), .C2(new_n361), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n364), .A2(KEYINPUT76), .A3(new_n365), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT76), .B1(new_n364), .B2(new_n365), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n366), .B(new_n370), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n333), .B1(new_n360), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375));
  XNOR2_X1  g174(.A(G155gat), .B(G162gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(new_n337), .A3(new_n338), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT2), .B1(new_n351), .B2(new_n343), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n377), .B1(new_n378), .B2(new_n342), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT82), .B1(new_n379), .B2(new_n352), .ZN(new_n380));
  AND4_X1   g179(.A1(KEYINPUT82), .A2(new_n350), .A3(new_n352), .A4(new_n353), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n340), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n375), .B1(new_n382), .B2(KEYINPUT3), .ZN(new_n383));
  INV_X1    g182(.A(new_n373), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(KEYINPUT87), .A3(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n371), .A2(new_n372), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n364), .A2(new_n365), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n375), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n358), .B1(new_n359), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G228gat), .A2(G233gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT77), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n373), .B(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT89), .B1(new_n360), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n373), .B(KEYINPUT77), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT89), .ZN(new_n397));
  AOI211_X1 g196(.A(KEYINPUT3), .B(new_n341), .C1(new_n356), .C2(new_n357), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n396), .B(new_n397), .C1(new_n398), .C2(KEYINPUT29), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT3), .B1(new_n373), .B2(new_n375), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(KEYINPUT88), .A3(new_n382), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT88), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n404), .B1(new_n358), .B2(new_n401), .ZN(new_n405));
  INV_X1    g204(.A(new_n392), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n391), .A2(new_n392), .B1(new_n400), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(G22gat), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT91), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT86), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT31), .B(G50gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT90), .B(G22gat), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n414), .B1(new_n408), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT91), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n383), .A2(new_n384), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n389), .B1(new_n418), .B2(new_n333), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n406), .B1(new_n419), .B2(new_n385), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n406), .A3(new_n405), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n395), .B2(new_n399), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n417), .B(G22gat), .C1(new_n420), .C2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n410), .A2(new_n416), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n391), .A2(new_n392), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n400), .A2(new_n407), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n425), .A2(new_n415), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n415), .B1(new_n425), .B2(new_n426), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n414), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G71gat), .B(G99gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(KEYINPUT73), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(G15gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(G43gat), .ZN(new_n434));
  XOR2_X1   g233(.A(G113gat), .B(G120gat), .Z(new_n435));
  INV_X1    g234(.A(KEYINPUT1), .ZN(new_n436));
  INV_X1    g235(.A(G127gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G134gat), .ZN(new_n438));
  INV_X1    g237(.A(G134gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(G127gat), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n435), .A2(new_n436), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT71), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n439), .A2(KEYINPUT70), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT70), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(G134gat), .ZN(new_n446));
  AND4_X1   g245(.A1(new_n443), .A2(new_n444), .A3(new_n446), .A4(G127gat), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n444), .A2(new_n446), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(G127gat), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n443), .B1(new_n437), .B2(G134gat), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G113gat), .B(G120gat), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT1), .B1(new_n452), .B2(KEYINPUT72), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(KEYINPUT72), .B2(new_n452), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n442), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT25), .ZN(new_n456));
  NAND2_X1  g255(.A1(G183gat), .A2(G190gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n457), .B(KEYINPUT67), .ZN(new_n458));
  XOR2_X1   g257(.A(KEYINPUT68), .B(KEYINPUT24), .Z(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT69), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(KEYINPUT69), .A3(new_n459), .ZN(new_n463));
  NOR2_X1   g262(.A1(G183gat), .A2(G190gat), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT24), .ZN(new_n465));
  INV_X1    g264(.A(G183gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n464), .B1(new_n467), .B2(G190gat), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n462), .A2(new_n463), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(G169gat), .A2(G176gat), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT66), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT23), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(G169gat), .B2(G176gat), .ZN(new_n474));
  NOR2_X1   g273(.A1(G169gat), .A2(G176gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT23), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n456), .B1(new_n469), .B2(new_n478), .ZN(new_n479));
  OR2_X1    g278(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n480));
  INV_X1    g279(.A(G169gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n480), .A2(KEYINPUT23), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  AND4_X1   g282(.A1(new_n456), .A2(new_n472), .A3(new_n474), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n457), .A2(KEYINPUT64), .A3(new_n465), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT64), .ZN(new_n486));
  INV_X1    g285(.A(new_n457), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n486), .B1(new_n487), .B2(KEYINPUT24), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n468), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G183gat), .ZN(new_n491));
  INV_X1    g290(.A(G190gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT28), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n491), .A2(KEYINPUT28), .A3(new_n492), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n475), .B(KEYINPUT26), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n487), .B1(new_n498), .B2(new_n472), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n490), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n455), .B1(new_n479), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G227gat), .ZN(new_n503));
  INV_X1    g302(.A(G233gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n451), .A2(new_n454), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n441), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n489), .A2(new_n484), .B1(new_n497), .B2(new_n499), .ZN(new_n508));
  INV_X1    g307(.A(new_n468), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n460), .B2(new_n461), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n477), .B1(new_n510), .B2(new_n463), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n507), .B(new_n508), .C1(new_n511), .C2(new_n456), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n502), .A2(new_n505), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT33), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n434), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(KEYINPUT32), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n513), .B(KEYINPUT32), .C1(new_n514), .C2(new_n434), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT34), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n512), .ZN(new_n521));
  INV_X1    g320(.A(new_n505), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI211_X1 g322(.A(KEYINPUT34), .B(new_n505), .C1(new_n502), .C2(new_n512), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n519), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n517), .A3(new_n518), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(KEYINPUT74), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n525), .B1(new_n517), .B2(new_n518), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT74), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n430), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n455), .B1(new_n382), .B2(KEYINPUT3), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(KEYINPUT3), .B2(new_n382), .ZN(new_n536));
  NAND2_X1  g335(.A1(G225gat), .A2(G233gat), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n340), .B(new_n455), .C1(new_n380), .C2(new_n381), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT4), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT4), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n358), .A2(new_n540), .A3(new_n455), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n536), .A2(new_n537), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT5), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n382), .A2(new_n507), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n538), .ZN(new_n546));
  INV_X1    g345(.A(new_n537), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT84), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(new_n538), .B2(KEYINPUT4), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n358), .A2(KEYINPUT84), .A3(new_n540), .A4(new_n455), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT85), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n538), .A2(new_n553), .A3(KEYINPUT4), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n538), .B2(KEYINPUT4), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n551), .B(new_n552), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n507), .B1(new_n358), .B2(new_n359), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n544), .B(new_n537), .C1(new_n557), .C2(new_n398), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n549), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G1gat), .B(G29gat), .Z(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G57gat), .B(G85gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n561), .A2(KEYINPUT6), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT6), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n543), .A2(new_n548), .B1(new_n556), .B2(new_n559), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n569), .B1(new_n570), .B2(new_n566), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n561), .A2(new_n567), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n568), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G226gat), .A2(G233gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n574), .B(KEYINPUT78), .Z(new_n575));
  OAI22_X1  g374(.A1(new_n479), .A2(new_n501), .B1(KEYINPUT29), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n508), .B(new_n577), .C1(new_n511), .C2(new_n456), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n396), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n384), .A3(new_n578), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G8gat), .B(G36gat), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT79), .ZN(new_n584));
  XNOR2_X1  g383(.A(G64gat), .B(G92gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n580), .A2(new_n588), .A3(new_n581), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n587), .A2(KEYINPUT30), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT30), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n582), .A2(new_n591), .A3(new_n586), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n573), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT35), .B1(new_n534), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT94), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT35), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n424), .A2(new_n429), .B1(new_n532), .B2(new_n529), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n590), .A2(new_n592), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n561), .A2(new_n567), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n570), .A2(new_n566), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(new_n601), .A3(new_n569), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n599), .B1(new_n602), .B2(new_n568), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n597), .B1(new_n598), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT94), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT93), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(new_n571), .B2(new_n572), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n600), .A2(new_n601), .A3(KEYINPUT93), .A4(new_n569), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(new_n568), .A3(new_n609), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n525), .A2(new_n517), .A3(new_n518), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(new_n530), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n599), .A2(KEYINPUT35), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n610), .A2(new_n430), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n596), .A2(new_n606), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n430), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n533), .A2(KEYINPUT36), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n612), .A2(KEYINPUT36), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n616), .A2(new_n594), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n556), .A2(new_n536), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT92), .B1(new_n621), .B2(new_n547), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT92), .ZN(new_n623));
  AOI211_X1 g422(.A(new_n623), .B(new_n537), .C1(new_n556), .C2(new_n536), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n620), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n557), .A2(new_n398), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n551), .A2(new_n552), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n539), .A2(KEYINPUT85), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n538), .A2(new_n553), .A3(KEYINPUT4), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n626), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n623), .B1(new_n631), .B2(new_n537), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n621), .A2(KEYINPUT92), .A3(new_n547), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n546), .A2(new_n547), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n634), .A2(new_n620), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n625), .A2(new_n566), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n625), .A2(new_n636), .A3(KEYINPUT40), .A4(new_n566), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n593), .B1(new_n567), .B2(new_n561), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT37), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n576), .A2(new_n578), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(new_n373), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n645), .B1(new_n394), .B2(new_n644), .ZN(new_n646));
  INV_X1    g445(.A(new_n581), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n643), .B1(new_n647), .B2(new_n579), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n646), .A2(new_n648), .A3(new_n649), .A4(new_n588), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n587), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n586), .B1(new_n582), .B2(new_n643), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n580), .A2(KEYINPUT37), .A3(new_n581), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n608), .A2(new_n655), .A3(new_n568), .A4(new_n609), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n430), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n619), .B1(new_n642), .B2(new_n657), .ZN(new_n658));
  AOI211_X1 g457(.A(new_n258), .B(new_n332), .C1(new_n615), .C2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n573), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT106), .B(G1gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1324gat));
  AND2_X1   g462(.A1(new_n659), .A2(new_n599), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT16), .B(G8gat), .Z(new_n665));
  AND2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(G8gat), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT42), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n669), .B1(KEYINPUT42), .B2(new_n666), .ZN(G1325gat));
  INV_X1    g469(.A(G15gat), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n659), .A2(new_n671), .A3(new_n612), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n617), .A2(new_n618), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n659), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n672), .B1(new_n674), .B2(new_n671), .ZN(G1326gat));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n616), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  INV_X1    g477(.A(G29gat), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n614), .B1(new_n604), .B2(new_n605), .ZN(new_n680));
  AOI211_X1 g479(.A(KEYINPUT94), .B(new_n597), .C1(new_n598), .C2(new_n603), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n658), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT109), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n615), .A2(KEYINPUT109), .A3(new_n658), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .A4(new_n280), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n682), .A2(new_n280), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n689), .B2(KEYINPUT44), .ZN(new_n690));
  AOI211_X1 g489(.A(KEYINPUT108), .B(new_n686), .C1(new_n682), .C2(new_n280), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n309), .A2(new_n258), .A3(new_n330), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(new_n660), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT110), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n679), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n695), .B2(new_n694), .ZN(new_n697));
  INV_X1    g496(.A(new_n693), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n689), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(new_n679), .A3(new_n660), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n697), .A2(new_n702), .ZN(G1328gat));
  INV_X1    g502(.A(G36gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n689), .A2(KEYINPUT44), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT108), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n689), .A2(new_n688), .A3(KEYINPUT44), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n698), .B1(new_n708), .B2(new_n687), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n704), .B1(new_n709), .B2(new_n599), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n699), .A2(new_n704), .A3(new_n599), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT112), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n711), .B(new_n712), .Z(new_n715));
  INV_X1    g514(.A(KEYINPUT112), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n692), .A2(new_n599), .A3(new_n693), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(new_n704), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n714), .A2(new_n718), .ZN(G1329gat));
  NAND3_X1  g518(.A1(new_n692), .A2(new_n673), .A3(new_n693), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n692), .A2(KEYINPUT113), .A3(new_n673), .A4(new_n693), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n722), .A2(G43gat), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n612), .ZN(new_n725));
  NOR4_X1   g524(.A1(new_n689), .A2(G43gat), .A3(new_n725), .A4(new_n698), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT47), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n720), .A2(G43gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n727), .B1(new_n730), .B2(new_n726), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(G1330gat));
  AOI21_X1  g531(.A(G50gat), .B1(new_n699), .B2(new_n616), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n616), .A2(G50gat), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n709), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1331gat));
  INV_X1    g536(.A(new_n309), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(new_n280), .ZN(new_n739));
  INV_X1    g538(.A(new_n258), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(new_n331), .ZN(new_n741));
  AND4_X1   g540(.A1(new_n739), .A2(new_n684), .A3(new_n685), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n660), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g543(.A(new_n593), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT114), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1333gat));
  NAND3_X1  g548(.A1(new_n742), .A2(new_n286), .A3(new_n612), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n742), .A2(new_n673), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(new_n286), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g552(.A1(new_n742), .A2(new_n616), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g554(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n740), .A2(new_n309), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n682), .A2(new_n280), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n760), .A2(new_n330), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(new_n262), .A3(new_n660), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n741), .A2(new_n738), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n708), .B2(new_n687), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n764), .A2(new_n660), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n765), .B2(new_n262), .ZN(G1336gat));
  INV_X1    g565(.A(new_n763), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n692), .A2(new_n599), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G92gat), .ZN(new_n769));
  OR2_X1    g568(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n331), .A2(new_n593), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(G92gat), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n760), .A2(new_n773), .B1(KEYINPUT116), .B2(KEYINPUT52), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n769), .A2(new_n770), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n770), .B1(new_n769), .B2(new_n774), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(G1337gat));
  INV_X1    g576(.A(G99gat), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n692), .A2(new_n673), .A3(new_n767), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n780), .B2(new_n779), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n761), .A2(new_n778), .A3(new_n612), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1338gat));
  INV_X1    g583(.A(G106gat), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n764), .B2(new_n616), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n430), .A2(G106gat), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n760), .A2(new_n330), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT53), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n788), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n692), .A2(new_n616), .A3(new_n767), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n790), .B(new_n791), .C1(new_n785), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n789), .A2(new_n793), .ZN(G1339gat));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n245), .A2(new_n246), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n234), .B1(new_n233), .B2(new_n240), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n253), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n330), .A2(new_n257), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n318), .A2(new_n319), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n321), .A2(new_n800), .A3(KEYINPUT54), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n326), .B1(new_n320), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n801), .A2(KEYINPUT55), .A3(new_n803), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(new_n329), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n799), .B1(new_n258), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT118), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n811), .B(new_n799), .C1(new_n258), .C2(new_n808), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n281), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n808), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n257), .A2(new_n798), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n280), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n309), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n332), .A2(new_n740), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n795), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n818), .ZN(new_n820));
  INV_X1    g619(.A(new_n816), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n280), .B1(new_n809), .B2(KEYINPUT118), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(new_n822), .B2(new_n812), .ZN(new_n823));
  OAI211_X1 g622(.A(KEYINPUT119), .B(new_n820), .C1(new_n823), .C2(new_n309), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n616), .A2(new_n725), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n660), .A2(new_n593), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n819), .A2(new_n824), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(G113gat), .B1(new_n828), .B2(new_n258), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT120), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n534), .A2(new_n599), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n819), .A2(new_n824), .A3(new_n660), .A4(new_n831), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n832), .A2(G113gat), .A3(new_n258), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n830), .A2(new_n833), .ZN(G1340gat));
  INV_X1    g633(.A(G120gat), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n828), .A2(new_n835), .A3(new_n331), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n832), .A2(new_n331), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n835), .ZN(G1341gat));
  OAI21_X1  g637(.A(G127gat), .B1(new_n828), .B2(new_n738), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n309), .A2(new_n437), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n832), .B2(new_n840), .ZN(G1342gat));
  OAI21_X1  g640(.A(G134gat), .B1(new_n828), .B2(new_n281), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n280), .A2(new_n448), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n832), .A2(new_n844), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n845), .A2(KEYINPUT121), .A3(new_n843), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT121), .B1(new_n845), .B2(new_n843), .ZN(new_n847));
  OAI221_X1 g646(.A(new_n842), .B1(new_n843), .B2(new_n845), .C1(new_n846), .C2(new_n847), .ZN(G1343gat));
  OR2_X1    g647(.A1(new_n673), .A2(new_n826), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n819), .A2(new_n824), .A3(new_n616), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n809), .A2(new_n281), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n738), .B1(new_n853), .B2(new_n821), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n818), .B1(new_n854), .B2(KEYINPUT122), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(KEYINPUT122), .B2(new_n854), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n430), .A2(new_n851), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n849), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n335), .B1(new_n859), .B2(new_n740), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n819), .A2(new_n824), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n573), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n673), .A2(new_n599), .A3(new_n430), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n862), .A2(new_n335), .A3(new_n740), .A4(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT58), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867));
  AOI211_X1 g666(.A(new_n258), .B(new_n849), .C1(new_n852), .C2(new_n858), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n864), .B(new_n867), .C1(new_n868), .C2(new_n335), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n869), .ZN(G1344gat));
  AOI211_X1 g669(.A(KEYINPUT59), .B(new_n336), .C1(new_n859), .C2(new_n330), .ZN(new_n871));
  XOR2_X1   g670(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n872));
  NAND3_X1  g671(.A1(new_n819), .A2(new_n824), .A3(new_n857), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n854), .A2(new_n820), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n851), .B1(new_n874), .B2(new_n430), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n849), .A2(new_n331), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n872), .B1(new_n878), .B2(G148gat), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n863), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n330), .A2(new_n336), .ZN(new_n881));
  OAI22_X1  g680(.A1(new_n871), .A2(new_n879), .B1(new_n880), .B2(new_n881), .ZN(G1345gat));
  INV_X1    g681(.A(new_n859), .ZN(new_n883));
  OAI21_X1  g682(.A(G155gat), .B1(new_n883), .B2(new_n738), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n309), .A2(new_n343), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n880), .B2(new_n885), .ZN(G1346gat));
  NOR2_X1   g685(.A1(new_n883), .A2(new_n281), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n280), .A2(new_n351), .ZN(new_n888));
  OAI22_X1  g687(.A1(new_n887), .A2(new_n351), .B1(new_n880), .B2(new_n888), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n660), .A2(new_n593), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n819), .A2(new_n824), .A3(new_n825), .A4(new_n890), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n891), .A2(new_n481), .A3(new_n258), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n861), .A2(new_n660), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n534), .A2(new_n593), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n740), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n892), .B1(new_n897), .B2(new_n481), .ZN(G1348gat));
  AOI21_X1  g697(.A(G176gat), .B1(new_n896), .B2(new_n330), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n331), .B(new_n891), .C1(new_n480), .C2(new_n482), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(G1349gat));
  NAND2_X1  g700(.A1(new_n309), .A2(new_n491), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n905));
  OAI21_X1  g704(.A(G183gat), .B1(new_n891), .B2(new_n738), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n903), .A2(new_n904), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n904), .B1(new_n895), .B2(new_n902), .ZN(new_n908));
  INV_X1    g707(.A(new_n906), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT60), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n907), .A2(new_n910), .ZN(G1350gat));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n913));
  OAI221_X1 g712(.A(G190gat), .B1(new_n912), .B2(new_n913), .C1(new_n891), .C2(new_n281), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n914), .B(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n896), .A2(new_n492), .A3(new_n280), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1351gat));
  NOR3_X1   g717(.A1(new_n673), .A2(new_n660), .A3(new_n593), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n876), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT126), .B1(new_n920), .B2(new_n258), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G197gat), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n920), .A2(KEYINPUT126), .A3(new_n258), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n673), .A2(new_n430), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n893), .A2(new_n599), .A3(new_n924), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n258), .A2(G197gat), .ZN(new_n926));
  OAI22_X1  g725(.A1(new_n922), .A2(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1352gat));
  NOR2_X1   g726(.A1(new_n772), .A2(G204gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n893), .A2(new_n924), .A3(new_n928), .ZN(new_n929));
  XOR2_X1   g728(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(G204gat), .B1(new_n920), .B2(new_n331), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n929), .A2(new_n931), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(G1353gat));
  NAND3_X1  g734(.A1(new_n876), .A2(new_n309), .A3(new_n919), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n738), .A2(G211gat), .ZN(new_n939));
  OAI22_X1  g738(.A1(new_n937), .A2(new_n938), .B1(new_n925), .B2(new_n939), .ZN(G1354gat));
  OAI21_X1  g739(.A(G218gat), .B1(new_n920), .B2(new_n281), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n281), .A2(G218gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n925), .B2(new_n942), .ZN(G1355gat));
endmodule


