//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930;
  NAND3_X1  g000(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT64), .ZN(new_n203));
  AOI21_X1  g002(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n204));
  INV_X1    g003(.A(G183gat), .ZN(new_n205));
  INV_X1    g004(.A(G190gat), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(new_n208), .B(KEYINPUT65), .Z(new_n209));
  NOR2_X1   g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n210), .A2(KEYINPUT23), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(KEYINPUT23), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT25), .B1(new_n209), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT25), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n217), .B1(new_n207), .B2(new_n202), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT70), .ZN(new_n222));
  AND2_X1   g021(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n206), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT28), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(KEYINPUT66), .B(new_n206), .C1(new_n223), .C2(new_n224), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n228), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n233), .ZN(new_n235));
  AOI211_X1 g034(.A(KEYINPUT68), .B(new_n235), .C1(new_n230), .C2(new_n231), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n227), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT69), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n239), .B(new_n227), .C1(new_n234), .C2(new_n236), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n210), .A2(KEYINPUT26), .ZN(new_n242));
  NAND2_X1  g041(.A1(G183gat), .A2(G190gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT26), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n212), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n242), .B(new_n243), .C1(new_n245), .C2(new_n210), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n222), .B1(new_n241), .B2(new_n247), .ZN(new_n248));
  AOI211_X1 g047(.A(KEYINPUT70), .B(new_n246), .C1(new_n238), .C2(new_n240), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n221), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G127gat), .B(G134gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT71), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(KEYINPUT72), .B(KEYINPUT1), .Z(new_n255));
  NAND3_X1  g054(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n257));
  OR2_X1    g056(.A1(new_n257), .A2(new_n251), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n250), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G227gat), .A2(G233gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n259), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n262), .B(new_n221), .C1(new_n248), .C2(new_n249), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT34), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n260), .A2(KEYINPUT34), .A3(new_n261), .A4(new_n263), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n260), .A2(new_n263), .ZN(new_n270));
  INV_X1    g069(.A(new_n261), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT32), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n270), .A2(new_n271), .B1(new_n272), .B2(KEYINPUT33), .ZN(new_n273));
  XNOR2_X1  g072(.A(G15gat), .B(G43gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(G99gat), .ZN(new_n275));
  XOR2_X1   g074(.A(KEYINPUT73), .B(G71gat), .Z(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(KEYINPUT74), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n277), .A2(KEYINPUT74), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT33), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  AOI211_X1 g082(.A(new_n272), .B(new_n283), .C1(new_n270), .C2(new_n271), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n269), .B1(new_n278), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT75), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n287));
  INV_X1    g086(.A(new_n283), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n287), .A2(KEYINPUT32), .A3(new_n288), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n268), .B(new_n289), .C1(new_n277), .C2(new_n273), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n285), .A2(new_n286), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT36), .ZN(new_n292));
  OAI211_X1 g091(.A(KEYINPUT75), .B(new_n269), .C1(new_n278), .C2(new_n284), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n285), .A2(KEYINPUT36), .A3(new_n290), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G78gat), .B(G106gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT82), .ZN(new_n298));
  XOR2_X1   g097(.A(KEYINPUT31), .B(G50gat), .Z(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301));
  OR2_X1    g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(G141gat), .B(G148gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT79), .B(KEYINPUT2), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n301), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n303), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n301), .B1(new_n302), .B2(KEYINPUT2), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G197gat), .B(G204gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT22), .ZN(new_n311));
  INV_X1    g110(.A(G211gat), .ZN(new_n312));
  INV_X1    g111(.A(G218gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT76), .ZN(new_n317));
  XOR2_X1   g116(.A(G211gat), .B(G218gat), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n319), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n316), .A2(new_n322), .A3(new_n319), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT77), .B1(new_n315), .B2(new_n318), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n317), .A2(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(KEYINPUT29), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT83), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n326), .A2(KEYINPUT83), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n309), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n325), .A2(KEYINPUT78), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n325), .A2(KEYINPUT78), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n309), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT29), .B1(new_n335), .B2(new_n328), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n336), .A2(KEYINPUT84), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(KEYINPUT84), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n334), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G228gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n331), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G22gat), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n323), .A2(new_n324), .B1(new_n318), .B2(new_n315), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n328), .B1(new_n344), .B2(KEYINPUT29), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n309), .B(KEYINPUT81), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n333), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n348), .B2(new_n336), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n340), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n342), .A2(new_n343), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n343), .B1(new_n342), .B2(new_n350), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n300), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n342), .A2(new_n350), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G22gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n342), .A2(new_n343), .A3(new_n350), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n300), .A2(KEYINPUT85), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n352), .A2(KEYINPUT85), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n353), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n361), .B(new_n221), .C1(new_n248), .C2(new_n249), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(KEYINPUT29), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n246), .B1(new_n238), .B2(new_n240), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n363), .B1(new_n220), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n334), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n220), .A2(new_n364), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n250), .A2(new_n363), .B1(new_n361), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n366), .B1(new_n334), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G8gat), .B(G36gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n369), .A2(KEYINPUT30), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT30), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n362), .A2(new_n365), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n348), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n367), .A2(new_n361), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT27), .B(G183gat), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT66), .B1(new_n379), .B2(new_n206), .ZN(new_n380));
  INV_X1    g179(.A(new_n231), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n233), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT68), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n232), .A2(new_n228), .A3(new_n233), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n239), .B1(new_n385), .B2(new_n227), .ZN(new_n386));
  INV_X1    g185(.A(new_n240), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n247), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT70), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n364), .A2(new_n222), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n220), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n363), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n334), .B(new_n378), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n375), .B1(new_n394), .B2(new_n372), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n372), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n374), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n259), .B(new_n309), .ZN(new_n398));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n259), .A2(KEYINPUT4), .A3(new_n309), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n346), .A2(new_n259), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n309), .B(new_n328), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n259), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n399), .ZN(new_n408));
  OAI211_X1 g207(.A(KEYINPUT5), .B(new_n401), .C1(new_n405), .C2(new_n408), .ZN(new_n409));
  OR3_X1    g208(.A1(new_n346), .A2(new_n259), .A3(new_n404), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT4), .B1(new_n259), .B2(new_n309), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n410), .A2(new_n411), .B1(new_n259), .B2(new_n406), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n400), .A2(KEYINPUT5), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G1gat), .B(G29gat), .ZN(new_n416));
  INV_X1    g215(.A(G85gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT0), .B(G57gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  NAND2_X1  g219(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n415), .A2(KEYINPUT86), .A3(new_n420), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OR3_X1    g224(.A1(new_n412), .A2(KEYINPUT39), .A3(new_n399), .ZN(new_n426));
  INV_X1    g225(.A(new_n420), .ZN(new_n427));
  OR2_X1    g226(.A1(new_n398), .A2(new_n400), .ZN(new_n428));
  OAI211_X1 g227(.A(KEYINPUT39), .B(new_n428), .C1(new_n412), .C2(new_n399), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT40), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n426), .A2(KEYINPUT40), .A3(new_n427), .A4(new_n429), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n425), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n360), .B1(new_n397), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n348), .B1(new_n362), .B2(new_n365), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n348), .B2(new_n368), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT38), .B1(new_n438), .B2(KEYINPUT37), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT37), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT87), .B1(new_n369), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n377), .A2(KEYINPUT87), .A3(new_n393), .A4(new_n440), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n372), .B(new_n439), .C1(new_n441), .C2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n445), .B1(new_n415), .B2(new_n420), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n446), .B1(new_n423), .B2(new_n424), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n394), .A2(new_n372), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n421), .A2(new_n445), .ZN(new_n449));
  NOR3_X1   g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT38), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n377), .A2(new_n440), .A3(new_n393), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT87), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n373), .B1(new_n455), .B2(new_n442), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n394), .A2(KEYINPUT37), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n452), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n436), .B1(new_n451), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n446), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n449), .B1(new_n421), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n360), .B1(new_n397), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT35), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n447), .B2(new_n449), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n353), .A2(new_n358), .A3(new_n359), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n466), .A2(new_n396), .A3(new_n374), .A4(new_n395), .ZN(new_n467));
  AOI211_X1 g266(.A(new_n465), .B(new_n467), .C1(new_n291), .C2(new_n293), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n285), .A2(new_n290), .A3(new_n466), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n397), .A2(new_n461), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI22_X1  g270(.A1(new_n296), .A2(new_n463), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  OR3_X1    g272(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n474), .A2(new_n475), .B1(G29gat), .B2(G36gat), .ZN(new_n476));
  INV_X1    g275(.A(G43gat), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n477), .A2(G50gat), .ZN(new_n478));
  XOR2_X1   g277(.A(KEYINPUT89), .B(G50gat), .Z(new_n479));
  AOI21_X1  g278(.A(new_n478), .B1(new_n479), .B2(new_n477), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n476), .B1(new_n480), .B2(KEYINPUT15), .ZN(new_n481));
  INV_X1    g280(.A(new_n478), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n477), .A2(G50gat), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(KEYINPUT15), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n476), .A2(KEYINPUT15), .A3(new_n483), .A4(new_n482), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT90), .B(KEYINPUT17), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT91), .ZN(new_n490));
  XOR2_X1   g289(.A(G15gat), .B(G22gat), .Z(new_n491));
  INV_X1    g290(.A(G1gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(KEYINPUT16), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT92), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n493), .B1(new_n496), .B2(new_n491), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT93), .ZN(new_n498));
  AOI21_X1  g297(.A(G8gat), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n497), .B(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n487), .A2(new_n501), .A3(new_n488), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n486), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT17), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n490), .A2(new_n500), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n500), .B(KEYINPUT94), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n487), .ZN(new_n507));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT18), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n510), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT94), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n500), .B(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n503), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n508), .B(KEYINPUT13), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n511), .A2(new_n512), .A3(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n521));
  XNOR2_X1  g320(.A(G113gat), .B(G141gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(G169gat), .B(G197gat), .Z(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT12), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n526), .B1(new_n512), .B2(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n520), .B(new_n528), .Z(new_n529));
  NOR2_X1   g328(.A1(new_n473), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n490), .A2(new_n502), .A3(new_n504), .ZN(new_n531));
  NAND2_X1  g330(.A1(G85gat), .A2(G92gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT100), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g333(.A1(G99gat), .A2(G106gat), .ZN(new_n535));
  INV_X1    g334(.A(G92gat), .ZN(new_n536));
  AOI22_X1  g335(.A1(KEYINPUT8), .A2(new_n535), .B1(new_n417), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G99gat), .B(G106gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  OR3_X1    g339(.A1(new_n531), .A2(KEYINPUT101), .A3(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n540), .A2(new_n487), .B1(KEYINPUT41), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT101), .B1(new_n531), .B2(new_n540), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G190gat), .B(G218gat), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n546), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n542), .A2(KEYINPUT41), .ZN(new_n550));
  XNOR2_X1  g349(.A(G134gat), .B(G162gat), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n550), .B(new_n551), .Z(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n552), .B1(new_n547), .B2(new_n548), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G127gat), .B(G155gat), .Z(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT97), .ZN(new_n559));
  XOR2_X1   g358(.A(KEYINPUT99), .B(G211gat), .Z(new_n560));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n559), .B(new_n562), .Z(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G57gat), .B(G64gat), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G71gat), .B(G78gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT96), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT98), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n574), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT98), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n506), .B1(new_n580), .B2(KEYINPUT21), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n205), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n581), .A2(new_n205), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n566), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n577), .A2(KEYINPUT21), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n581), .A2(new_n205), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(new_n565), .A3(new_n582), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n585), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n587), .B1(new_n585), .B2(new_n589), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n564), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n589), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n565), .B1(new_n588), .B2(new_n582), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n586), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(new_n590), .A3(new_n563), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G230gat), .ZN(new_n599));
  INV_X1    g398(.A(G233gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n580), .A2(KEYINPUT10), .A3(new_n540), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n540), .A2(new_n571), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n575), .A2(new_n540), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n601), .B1(new_n602), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n601), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n605), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G120gat), .B(G148gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(G176gat), .B(G204gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  OR3_X1    g412(.A1(new_n608), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n613), .B1(new_n608), .B2(new_n610), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(KEYINPUT102), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT102), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n617), .B(new_n613), .C1(new_n608), .C2(new_n610), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n557), .A2(new_n598), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT103), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n530), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n461), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(new_n492), .ZN(G1324gat));
  INV_X1    g424(.A(new_n397), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT16), .B(G8gat), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT42), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n627), .A2(KEYINPUT42), .A3(new_n628), .ZN(new_n632));
  INV_X1    g431(.A(G8gat), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n627), .ZN(G1325gat));
  INV_X1    g433(.A(new_n622), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n635), .A2(G15gat), .A3(new_n296), .ZN(new_n636));
  INV_X1    g435(.A(new_n291), .ZN(new_n637));
  INV_X1    g436(.A(new_n293), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(G15gat), .B1(new_n635), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n636), .B1(new_n643), .B2(new_n644), .ZN(G1326gat));
  NOR2_X1   g444(.A1(new_n622), .A2(new_n466), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT43), .B(G22gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1327gat));
  INV_X1    g447(.A(new_n619), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n473), .A2(new_n529), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n557), .A2(new_n598), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n652), .A2(G29gat), .A3(new_n623), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT45), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n591), .A2(new_n592), .A3(new_n564), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n563), .B1(new_n596), .B2(new_n590), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(KEYINPUT105), .B1(new_n593), .B2(new_n597), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n529), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(new_n662), .A3(new_n619), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT106), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n472), .A2(new_n556), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n472), .B2(new_n556), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n664), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n461), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(G29gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n655), .A2(new_n673), .ZN(G1328gat));
  NOR3_X1   g473(.A1(new_n652), .A2(G36gat), .A3(new_n626), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT46), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n397), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(G36gat), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(G1329gat));
  OAI21_X1  g478(.A(new_n477), .B1(new_n652), .B2(new_n639), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n671), .A2(G43gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n296), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT47), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n685), .B(new_n680), .C1(new_n681), .C2(new_n682), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(G1330gat));
  NAND2_X1  g486(.A1(new_n652), .A2(KEYINPUT107), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n650), .A2(new_n689), .A3(new_n651), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n479), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n360), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT108), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n671), .A2(new_n360), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n479), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n695), .A2(new_n697), .A3(KEYINPUT48), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT48), .ZN(new_n699));
  INV_X1    g498(.A(new_n694), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n688), .B2(new_n690), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n692), .B1(new_n671), .B2(new_n360), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n698), .A2(new_n703), .ZN(G1331gat));
  NAND4_X1  g503(.A1(new_n557), .A2(new_n529), .A3(new_n598), .A4(new_n649), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT109), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n473), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n461), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g508(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n707), .A2(new_n397), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n711), .B(new_n712), .Z(G1333gat));
  NOR3_X1   g512(.A1(new_n473), .A2(new_n639), .A3(new_n706), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n714), .A2(G71gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n707), .A2(G71gat), .A3(new_n296), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n715), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT50), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT50), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n722), .B(new_n715), .C1(new_n718), .C2(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(G1334gat));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n360), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT111), .B(G78gat), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1335gat));
  NOR2_X1   g526(.A1(new_n598), .A2(new_n662), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n649), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT112), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n665), .A2(KEYINPUT44), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n731), .B2(new_n669), .ZN(new_n732));
  OAI21_X1  g531(.A(G85gat), .B1(new_n732), .B2(new_n623), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n472), .A2(new_n556), .A3(new_n728), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n472), .A2(KEYINPUT51), .A3(new_n556), .A4(new_n728), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n736), .A2(KEYINPUT113), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n666), .A2(new_n739), .A3(KEYINPUT51), .A4(new_n728), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n619), .A2(new_n623), .A3(G85gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT114), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n738), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n733), .A2(new_n743), .ZN(G1336gat));
  OAI21_X1  g543(.A(G92gat), .B1(new_n732), .B2(new_n626), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n626), .A2(G92gat), .A3(new_n619), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n738), .A2(new_n740), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT116), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n736), .A2(new_n750), .A3(new_n737), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n746), .A2(KEYINPUT115), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n734), .A2(KEYINPUT116), .A3(new_n735), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n746), .A2(KEYINPUT115), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n751), .A2(new_n752), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n745), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n749), .B1(new_n756), .B2(new_n748), .ZN(G1337gat));
  NOR2_X1   g556(.A1(new_n639), .A2(G99gat), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n738), .A2(new_n740), .A3(new_n649), .A4(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n296), .B(new_n730), .C1(new_n731), .C2(new_n669), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G99gat), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT117), .ZN(G1338gat));
  NOR2_X1   g562(.A1(new_n466), .A2(G106gat), .ZN(new_n764));
  AND4_X1   g563(.A1(new_n649), .A2(new_n751), .A3(new_n753), .A4(new_n764), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n360), .B(new_n730), .C1(new_n731), .C2(new_n669), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n766), .A2(G106gat), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT53), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  AND4_X1   g568(.A1(new_n649), .A2(new_n738), .A3(new_n740), .A4(new_n764), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT118), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n766), .B2(G106gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n738), .A2(new_n740), .A3(new_n649), .A4(new_n764), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n771), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n768), .B1(new_n773), .B2(new_n775), .ZN(G1339gat));
  NOR2_X1   g575(.A1(new_n659), .A2(new_n660), .ZN(new_n777));
  INV_X1    g576(.A(new_n613), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n608), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n538), .B(new_n539), .Z(new_n781));
  AOI211_X1 g580(.A(new_n603), .B(new_n781), .C1(new_n576), .C2(new_n579), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n577), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT10), .B1(new_n783), .B2(new_n604), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n609), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n602), .A2(new_n607), .A3(new_n601), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(KEYINPUT54), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n780), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n780), .A2(new_n787), .A3(KEYINPUT55), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n790), .A2(new_n614), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n516), .A2(new_n518), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n508), .B1(new_n505), .B2(new_n507), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n525), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n795), .A2(KEYINPUT119), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n511), .A2(new_n512), .A3(new_n526), .A4(new_n519), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(KEYINPUT119), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n529), .A2(new_n792), .B1(new_n619), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT120), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT120), .ZN(new_n802));
  OAI221_X1 g601(.A(new_n802), .B1(new_n619), .B2(new_n799), .C1(new_n529), .C2(new_n792), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(new_n557), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n792), .ZN(new_n805));
  INV_X1    g604(.A(new_n799), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n556), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n777), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n557), .A2(new_n529), .A3(new_n598), .A4(new_n619), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n639), .A2(new_n467), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n461), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(G113gat), .B1(new_n813), .B2(new_n529), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n397), .A2(new_n623), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n469), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n817), .A2(G113gat), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n814), .B1(new_n818), .B2(new_n529), .ZN(G1340gat));
  OAI21_X1  g618(.A(G120gat), .B1(new_n813), .B2(new_n619), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n817), .A2(G120gat), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n821), .B2(new_n619), .ZN(G1341gat));
  INV_X1    g621(.A(G127gat), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n813), .A2(new_n823), .A3(new_n661), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n811), .A2(new_n598), .A3(new_n816), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n823), .B2(new_n825), .ZN(G1342gat));
  NOR2_X1   g625(.A1(new_n557), .A2(G134gat), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n816), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n811), .A2(new_n461), .A3(new_n812), .A4(new_n556), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT121), .B1(new_n831), .B2(G134gat), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n831), .A2(KEYINPUT121), .A3(G134gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n830), .B(KEYINPUT122), .C1(new_n832), .C2(new_n833), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1343gat));
  INV_X1    g637(.A(G141gat), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  INV_X1    g639(.A(new_n810), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n840), .B(new_n360), .C1(new_n808), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n557), .A2(new_n800), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n598), .B1(new_n843), .B2(new_n807), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n360), .B1(new_n844), .B2(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT57), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n296), .A2(new_n623), .A3(new_n397), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n842), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT123), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT123), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n842), .A2(new_n846), .A3(new_n850), .A4(new_n847), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n839), .B1(new_n852), .B2(new_n662), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n466), .B1(new_n809), .B2(new_n810), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(new_n847), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n855), .A2(new_n839), .A3(new_n662), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT58), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n856), .A2(KEYINPUT58), .ZN(new_n858));
  OAI21_X1  g657(.A(G141gat), .B1(new_n848), .B2(new_n529), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n857), .A2(new_n860), .ZN(G1344gat));
  AOI21_X1  g660(.A(new_n619), .B1(new_n849), .B2(new_n851), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n854), .A2(new_n840), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n621), .A2(new_n529), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n840), .B(new_n360), .C1(new_n864), .C2(new_n844), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n649), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n847), .A2(KEYINPUT59), .ZN(new_n867));
  OAI22_X1  g666(.A1(new_n862), .A2(KEYINPUT59), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(G148gat), .B1(new_n855), .B2(new_n649), .ZN(new_n869));
  AOI22_X1  g668(.A1(new_n868), .A2(G148gat), .B1(KEYINPUT59), .B2(new_n869), .ZN(G1345gat));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n598), .A3(new_n847), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(KEYINPUT124), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(KEYINPUT124), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n872), .A2(new_n873), .A3(G155gat), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n661), .B1(new_n849), .B2(new_n851), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(G155gat), .B2(new_n875), .ZN(G1346gat));
  AOI21_X1  g675(.A(G162gat), .B1(new_n855), .B2(new_n556), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n557), .B1(new_n849), .B2(new_n851), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(G162gat), .ZN(G1347gat));
  AOI21_X1  g678(.A(new_n461), .B1(new_n809), .B2(new_n810), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n626), .A2(new_n360), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n640), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G169gat), .B1(new_n882), .B2(new_n529), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT126), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n881), .A2(new_n290), .A3(new_n285), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT125), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(G169gat), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n884), .B1(new_n888), .B2(new_n662), .ZN(new_n889));
  NOR4_X1   g688(.A1(new_n887), .A2(KEYINPUT126), .A3(G169gat), .A4(new_n529), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n883), .B1(new_n889), .B2(new_n890), .ZN(G1348gat));
  INV_X1    g690(.A(new_n887), .ZN(new_n892));
  AOI21_X1  g691(.A(G176gat), .B1(new_n892), .B2(new_n649), .ZN(new_n893));
  INV_X1    g692(.A(G176gat), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n882), .A2(new_n894), .A3(new_n619), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n893), .A2(new_n895), .ZN(G1349gat));
  NAND3_X1  g695(.A1(new_n892), .A2(new_n379), .A3(new_n598), .ZN(new_n897));
  OAI21_X1  g696(.A(G183gat), .B1(new_n882), .B2(new_n661), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g699(.A1(new_n892), .A2(new_n206), .A3(new_n556), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n882), .A2(new_n557), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n903), .A3(G190gat), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n903), .B1(new_n902), .B2(G190gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(G1351gat));
  NAND3_X1  g706(.A1(new_n682), .A2(new_n623), .A3(new_n397), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n863), .A2(new_n865), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G197gat), .B1(new_n910), .B2(new_n529), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n854), .A2(new_n909), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n912), .A2(G197gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n911), .B1(new_n529), .B2(new_n913), .ZN(G1352gat));
  NOR3_X1   g713(.A1(new_n912), .A2(G204gat), .A3(new_n619), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT62), .ZN(new_n916));
  OAI21_X1  g715(.A(G204gat), .B1(new_n866), .B2(new_n908), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1353gat));
  NAND4_X1  g717(.A1(new_n863), .A2(new_n598), .A3(new_n865), .A4(new_n909), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT63), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT127), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n919), .A2(G211gat), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n920), .A2(KEYINPUT127), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n854), .A2(new_n312), .A3(new_n598), .A4(new_n909), .ZN(new_n925));
  INV_X1    g724(.A(new_n923), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n919), .A2(G211gat), .A3(new_n926), .A4(new_n921), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(G1354gat));
  OAI21_X1  g727(.A(G218gat), .B1(new_n910), .B2(new_n557), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n556), .A2(new_n313), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n912), .B2(new_n930), .ZN(G1355gat));
endmodule


