

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776;

  XNOR2_X1 U371 ( .A(n510), .B(n509), .ZN(n579) );
  NOR2_X1 U372 ( .A1(n587), .A2(n586), .ZN(n448) );
  NOR2_X1 U373 ( .A1(G953), .A2(G237), .ZN(n519) );
  AND2_X1 U374 ( .A1(n720), .A2(n589), .ZN(n590) );
  BUF_X1 U375 ( .A(n668), .Z(n678) );
  XNOR2_X1 U376 ( .A(n585), .B(KEYINPUT104), .ZN(n598) );
  XNOR2_X2 U377 ( .A(n548), .B(n547), .ZN(n375) );
  AND2_X2 U378 ( .A1(n389), .A2(n419), .ZN(n548) );
  OR2_X2 U379 ( .A1(n665), .A2(KEYINPUT47), .ZN(n452) );
  NOR2_X2 U380 ( .A1(n608), .A2(n607), .ZN(n627) );
  OR2_X2 U381 ( .A1(n775), .A2(n634), .ZN(n636) );
  XNOR2_X2 U382 ( .A(n362), .B(n360), .ZN(n756) );
  NOR2_X2 U383 ( .A1(n697), .A2(n553), .ZN(n546) );
  XNOR2_X2 U384 ( .A(n605), .B(n552), .ZN(n588) );
  INV_X1 U385 ( .A(G146), .ZN(n366) );
  INV_X2 U386 ( .A(G953), .ZN(n768) );
  BUF_X1 U387 ( .A(n644), .Z(n767) );
  AND2_X1 U388 ( .A1(n380), .A2(n545), .ZN(n587) );
  NAND2_X1 U389 ( .A1(n385), .A2(n384), .ZN(n720) );
  INV_X2 U390 ( .A(G143), .ZN(n465) );
  AND2_X1 U391 ( .A1(n405), .A2(n401), .ZN(n400) );
  NOR2_X1 U392 ( .A1(n515), .A2(n514), .ZN(n736) );
  XNOR2_X1 U393 ( .A(n630), .B(KEYINPUT39), .ZN(n640) );
  INV_X1 U394 ( .A(n579), .ZN(n545) );
  INV_X1 U395 ( .A(n605), .ZN(n697) );
  AND2_X1 U396 ( .A1(n422), .A2(n436), .ZN(n392) );
  NAND2_X1 U397 ( .A1(n421), .A2(n440), .ZN(n420) );
  NAND2_X1 U398 ( .A1(n400), .A2(n399), .ZN(n644) );
  XNOR2_X1 U399 ( .A(n379), .B(n378), .ZN(n586) );
  OR2_X1 U400 ( .A1(n368), .A2(n601), .ZN(n597) );
  XNOR2_X1 U401 ( .A(n595), .B(KEYINPUT31), .ZN(n747) );
  XNOR2_X1 U402 ( .A(n505), .B(n504), .ZN(n530) );
  XNOR2_X2 U403 ( .A(n376), .B(n493), .ZN(n653) );
  AND2_X1 U404 ( .A1(n667), .A2(n597), .ZN(n445) );
  INV_X1 U405 ( .A(KEYINPUT48), .ZN(n449) );
  INV_X1 U406 ( .A(G237), .ZN(n469) );
  NOR2_X1 U407 ( .A1(n608), .A2(n563), .ZN(n544) );
  XNOR2_X1 U408 ( .A(n565), .B(KEYINPUT22), .ZN(n577) );
  BUF_X1 U409 ( .A(n698), .Z(n391) );
  NAND2_X1 U410 ( .A1(n653), .A2(n536), .ZN(n494) );
  XNOR2_X1 U411 ( .A(n432), .B(n453), .ZN(n489) );
  XNOR2_X1 U412 ( .A(n454), .B(G113), .ZN(n453) );
  XNOR2_X1 U413 ( .A(n460), .B(n455), .ZN(n432) );
  INV_X1 U414 ( .A(G116), .ZN(n454) );
  NAND2_X1 U415 ( .A1(n404), .A2(n403), .ZN(n402) );
  INV_X1 U416 ( .A(KEYINPUT85), .ZN(n403) );
  INV_X1 U417 ( .A(n639), .ZN(n404) );
  AND2_X1 U418 ( .A1(n639), .A2(KEYINPUT85), .ZN(n406) );
  INV_X1 U419 ( .A(KEYINPUT65), .ZN(n439) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n363) );
  INV_X1 U421 ( .A(KEYINPUT88), .ZN(n364) );
  NAND2_X1 U422 ( .A1(n599), .A2(n598), .ZN(n365) );
  INV_X1 U423 ( .A(G134), .ZN(n491) );
  XNOR2_X1 U424 ( .A(n502), .B(n501), .ZN(n521) );
  XNOR2_X1 U425 ( .A(n500), .B(KEYINPUT10), .ZN(n501) );
  INV_X1 U426 ( .A(G140), .ZN(n500) );
  XNOR2_X1 U427 ( .A(n518), .B(n516), .ZN(n417) );
  XNOR2_X1 U428 ( .A(KEYINPUT78), .B(KEYINPUT4), .ZN(n462) );
  XNOR2_X1 U429 ( .A(n464), .B(n428), .ZN(n427) );
  XNOR2_X1 U430 ( .A(KEYINPUT91), .B(KEYINPUT18), .ZN(n464) );
  XNOR2_X1 U431 ( .A(KEYINPUT92), .B(KEYINPUT17), .ZN(n428) );
  AND2_X1 U432 ( .A1(n699), .A2(n388), .ZN(n382) );
  AND2_X1 U433 ( .A1(n698), .A2(n588), .ZN(n383) );
  XNOR2_X1 U434 ( .A(n525), .B(n524), .ZN(n591) );
  XNOR2_X1 U435 ( .A(n523), .B(n522), .ZN(n524) );
  NOR2_X1 U436 ( .A1(n658), .A2(G902), .ZN(n525) );
  XNOR2_X1 U437 ( .A(n473), .B(n472), .ZN(n559) );
  NAND2_X1 U438 ( .A1(n474), .A2(G214), .ZN(n713) );
  NAND2_X1 U439 ( .A1(n669), .A2(n536), .ZN(n510) );
  INV_X1 U440 ( .A(KEYINPUT97), .ZN(n457) );
  XNOR2_X1 U441 ( .A(n486), .B(n488), .ZN(n458) );
  XNOR2_X1 U442 ( .A(n498), .B(n357), .ZN(n429) );
  XOR2_X1 U443 ( .A(G119), .B(KEYINPUT23), .Z(n507) );
  XNOR2_X1 U444 ( .A(n521), .B(n503), .ZN(n766) );
  INV_X1 U445 ( .A(KEYINPUT8), .ZN(n504) );
  NAND2_X1 U446 ( .A1(n768), .A2(G234), .ZN(n505) );
  XNOR2_X1 U447 ( .A(G107), .B(KEYINPUT102), .ZN(n526) );
  XOR2_X1 U448 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n527) );
  XNOR2_X1 U449 ( .A(G116), .B(G122), .ZN(n529) );
  XNOR2_X1 U450 ( .A(G101), .B(G140), .ZN(n495) );
  XOR2_X1 U451 ( .A(G137), .B(KEYINPUT68), .Z(n503) );
  NAND2_X1 U452 ( .A1(n434), .A2(n442), .ZN(n441) );
  NOR2_X1 U453 ( .A1(n767), .A2(n444), .ZN(n434) );
  NOR2_X1 U454 ( .A1(n397), .A2(n396), .ZN(n554) );
  NAND2_X1 U455 ( .A1(n588), .A2(n398), .ZN(n397) );
  NAND2_X1 U456 ( .A1(n412), .A2(KEYINPUT36), .ZN(n411) );
  INV_X1 U457 ( .A(n355), .ZN(n412) );
  NOR2_X1 U458 ( .A1(n581), .A2(n588), .ZN(n583) );
  NOR2_X1 U459 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U460 ( .A(n395), .B(n394), .ZN(n689) );
  INV_X1 U461 ( .A(n441), .ZN(n691) );
  NOR2_X1 U462 ( .A1(n736), .A2(n747), .ZN(n368) );
  NAND2_X1 U463 ( .A1(n597), .A2(n447), .ZN(n446) );
  INV_X1 U464 ( .A(KEYINPUT44), .ZN(n447) );
  AND2_X1 U465 ( .A1(n402), .A2(n641), .ZN(n401) );
  NAND2_X1 U466 ( .A1(n361), .A2(n437), .ZN(n436) );
  NAND2_X1 U467 ( .A1(n443), .A2(n438), .ZN(n437) );
  NAND2_X1 U468 ( .A1(KEYINPUT2), .A2(n439), .ZN(n438) );
  AND2_X1 U469 ( .A1(n444), .A2(KEYINPUT65), .ZN(n440) );
  NAND2_X1 U470 ( .A1(G234), .A2(G237), .ZN(n477) );
  XNOR2_X1 U471 ( .A(n591), .B(KEYINPUT100), .ZN(n549) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n521), .B(n350), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n520), .B(n517), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n753), .B(n468), .ZN(n646) );
  XNOR2_X1 U476 ( .A(n427), .B(n426), .ZN(n466) );
  INV_X1 U477 ( .A(KEYINPUT84), .ZN(n394) );
  NAND2_X1 U478 ( .A1(n593), .A2(KEYINPUT33), .ZN(n384) );
  AND2_X1 U479 ( .A1(n387), .A2(n386), .ZN(n385) );
  AND2_X1 U480 ( .A1(n555), .A2(n713), .ZN(n620) );
  XNOR2_X1 U481 ( .A(n476), .B(n349), .ZN(n377) );
  NAND2_X1 U482 ( .A1(n559), .A2(n713), .ZN(n476) );
  INV_X1 U483 ( .A(KEYINPUT95), .ZN(n390) );
  XNOR2_X1 U484 ( .A(n458), .B(n456), .ZN(n490) );
  XNOR2_X1 U485 ( .A(n487), .B(n457), .ZN(n456) );
  XNOR2_X1 U486 ( .A(n374), .B(n373), .ZN(n372) );
  XNOR2_X1 U487 ( .A(n507), .B(KEYINPUT24), .ZN(n373) );
  XNOR2_X1 U488 ( .A(n506), .B(n356), .ZN(n374) );
  XNOR2_X1 U489 ( .A(n535), .B(n534), .ZN(n674) );
  XNOR2_X1 U490 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n423) );
  XNOR2_X1 U492 ( .A(n503), .B(n497), .ZN(n424) );
  NOR2_X1 U493 ( .A1(n409), .A2(n408), .ZN(n750) );
  NAND2_X1 U494 ( .A1(n413), .A2(n410), .ZN(n409) );
  AND2_X1 U495 ( .A1(n622), .A2(n411), .ZN(n410) );
  INV_X1 U496 ( .A(n610), .ZN(n370) );
  INV_X1 U497 ( .A(KEYINPUT32), .ZN(n378) );
  NAND2_X1 U498 ( .A1(n570), .A2(n569), .ZN(n379) );
  AND2_X2 U499 ( .A1(n375), .A2(n377), .ZN(n665) );
  XNOR2_X1 U500 ( .A(n578), .B(n381), .ZN(n380) );
  INV_X1 U501 ( .A(KEYINPUT66), .ZN(n381) );
  INV_X1 U502 ( .A(KEYINPUT87), .ZN(n582) );
  NOR2_X1 U503 ( .A1(n734), .A2(n733), .ZN(n735) );
  INV_X1 U504 ( .A(n756), .ZN(n442) );
  XOR2_X1 U505 ( .A(n475), .B(KEYINPUT19), .Z(n349) );
  XNOR2_X1 U506 ( .A(G122), .B(G113), .ZN(n350) );
  XOR2_X1 U507 ( .A(n528), .B(KEYINPUT101), .Z(n351) );
  XNOR2_X1 U508 ( .A(KEYINPUT4), .B(G131), .ZN(n352) );
  XOR2_X1 U509 ( .A(n483), .B(KEYINPUT94), .Z(n353) );
  OR2_X1 U510 ( .A1(n600), .A2(KEYINPUT44), .ZN(n354) );
  AND2_X1 U511 ( .A1(n619), .A2(n713), .ZN(n355) );
  INV_X1 U512 ( .A(n396), .ZN(n743) );
  NAND2_X1 U513 ( .A1(n549), .A2(n562), .ZN(n396) );
  XOR2_X1 U514 ( .A(G128), .B(G110), .Z(n356) );
  XOR2_X1 U515 ( .A(KEYINPUT16), .B(G122), .Z(n357) );
  XNOR2_X1 U516 ( .A(n366), .B(G125), .ZN(n502) );
  XNOR2_X1 U517 ( .A(KEYINPUT79), .B(KEYINPUT35), .ZN(n358) );
  XOR2_X1 U518 ( .A(KEYINPUT71), .B(KEYINPUT34), .Z(n359) );
  XOR2_X1 U519 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n360) );
  XNOR2_X1 U520 ( .A(n372), .B(n766), .ZN(n669) );
  XNOR2_X1 U521 ( .A(n429), .B(n489), .ZN(n753) );
  XNOR2_X1 U522 ( .A(n418), .B(n415), .ZN(n658) );
  OR2_X1 U523 ( .A1(n443), .A2(KEYINPUT65), .ZN(n361) );
  INV_X1 U524 ( .A(n643), .ZN(n443) );
  XNOR2_X1 U525 ( .A(G902), .B(KEYINPUT15), .ZN(n643) );
  INV_X1 U526 ( .A(KEYINPUT2), .ZN(n444) );
  OR2_X1 U527 ( .A1(n407), .A2(KEYINPUT85), .ZN(n399) );
  NAND2_X1 U528 ( .A1(n363), .A2(n354), .ZN(n362) );
  XNOR2_X2 U529 ( .A(n367), .B(n366), .ZN(n376) );
  XNOR2_X1 U530 ( .A(n367), .B(KEYINPUT126), .ZN(n765) );
  XNOR2_X2 U531 ( .A(n531), .B(n352), .ZN(n367) );
  XNOR2_X2 U532 ( .A(n369), .B(n358), .ZN(n667) );
  NAND2_X1 U533 ( .A1(n371), .A2(n370), .ZN(n369) );
  XNOR2_X1 U534 ( .A(n590), .B(n359), .ZN(n371) );
  NAND2_X1 U535 ( .A1(n375), .A2(n729), .ZN(n576) );
  XNOR2_X1 U536 ( .A(n376), .B(n423), .ZN(n682) );
  NAND2_X1 U537 ( .A1(n377), .A2(n353), .ZN(n485) );
  NAND2_X1 U538 ( .A1(n383), .A2(n382), .ZN(n387) );
  NAND2_X1 U539 ( .A1(n698), .A2(n699), .ZN(n593) );
  OR2_X1 U540 ( .A1(n588), .A2(n388), .ZN(n386) );
  INV_X1 U541 ( .A(KEYINPUT33), .ZN(n388) );
  XNOR2_X2 U542 ( .A(n419), .B(KEYINPUT1), .ZN(n698) );
  XNOR2_X1 U543 ( .A(n546), .B(KEYINPUT28), .ZN(n389) );
  NOR2_X1 U544 ( .A1(n643), .A2(KEYINPUT65), .ZN(n435) );
  XNOR2_X1 U545 ( .A(n594), .B(n390), .ZN(n589) );
  XNOR2_X2 U546 ( .A(n485), .B(n484), .ZN(n594) );
  NAND2_X1 U547 ( .A1(n392), .A2(n420), .ZN(n433) );
  XNOR2_X1 U548 ( .A(n450), .B(n449), .ZN(n407) );
  NAND2_X1 U549 ( .A1(n393), .A2(n446), .ZN(n599) );
  NAND2_X1 U550 ( .A1(n445), .A2(n448), .ZN(n393) );
  NAND2_X1 U551 ( .A1(n756), .A2(n444), .ZN(n395) );
  INV_X1 U552 ( .A(n553), .ZN(n398) );
  NAND2_X1 U553 ( .A1(n407), .A2(n406), .ZN(n405) );
  NOR2_X1 U554 ( .A1(n555), .A2(n621), .ZN(n408) );
  NAND2_X1 U555 ( .A1(n555), .A2(n414), .ZN(n413) );
  AND2_X1 U556 ( .A1(n355), .A2(n621), .ZN(n414) );
  NAND2_X1 U557 ( .A1(n699), .A2(n419), .ZN(n612) );
  XNOR2_X2 U558 ( .A(n499), .B(G469), .ZN(n419) );
  INV_X1 U559 ( .A(n642), .ZN(n421) );
  NAND2_X1 U560 ( .A1(n642), .A2(n435), .ZN(n422) );
  XNOR2_X1 U561 ( .A(n498), .B(n496), .ZN(n425) );
  XNOR2_X2 U562 ( .A(n492), .B(n491), .ZN(n531) );
  INV_X1 U563 ( .A(n492), .ZN(n426) );
  NOR2_X2 U564 ( .A1(n577), .A2(n391), .ZN(n580) );
  INV_X1 U565 ( .A(n767), .ZN(n687) );
  NOR2_X2 U566 ( .A1(n756), .A2(n644), .ZN(n642) );
  XNOR2_X2 U567 ( .A(n431), .B(n430), .ZN(n498) );
  XNOR2_X2 U568 ( .A(KEYINPUT75), .B(G110), .ZN(n430) );
  XNOR2_X2 U569 ( .A(G107), .B(G104), .ZN(n431) );
  AND2_X2 U570 ( .A1(n433), .A2(n441), .ZN(n668) );
  NAND2_X1 U571 ( .A1(n448), .A2(n667), .ZN(n600) );
  NAND2_X1 U572 ( .A1(n638), .A2(n637), .ZN(n450) );
  NAND2_X1 U573 ( .A1(n452), .A2(n451), .ZN(n616) );
  NAND2_X1 U574 ( .A1(n665), .A2(n602), .ZN(n451) );
  XNOR2_X2 U575 ( .A(G101), .B(KEYINPUT70), .ZN(n455) );
  BUF_X1 U576 ( .A(n559), .Z(n619) );
  AND2_X1 U577 ( .A1(G217), .A2(n511), .ZN(n459) );
  INV_X1 U578 ( .A(n531), .ZN(n532) );
  XNOR2_X2 U579 ( .A(KEYINPUT3), .B(G119), .ZN(n460) );
  NAND2_X1 U580 ( .A1(n768), .A2(G224), .ZN(n461) );
  XNOR2_X1 U581 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U582 ( .A(n502), .B(n463), .ZN(n467) );
  XNOR2_X2 U583 ( .A(n465), .B(G128), .ZN(n492) );
  XNOR2_X1 U584 ( .A(n467), .B(n466), .ZN(n468) );
  NAND2_X1 U585 ( .A1(n646), .A2(n643), .ZN(n473) );
  INV_X1 U586 ( .A(G902), .ZN(n536) );
  NAND2_X1 U587 ( .A1(n536), .A2(n469), .ZN(n474) );
  NAND2_X1 U588 ( .A1(n474), .A2(G210), .ZN(n471) );
  INV_X1 U589 ( .A(KEYINPUT80), .ZN(n470) );
  XNOR2_X1 U590 ( .A(n471), .B(n470), .ZN(n472) );
  INV_X1 U591 ( .A(KEYINPUT76), .ZN(n475) );
  XOR2_X1 U592 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n478) );
  XNOR2_X1 U593 ( .A(n478), .B(n477), .ZN(n480) );
  NAND2_X1 U594 ( .A1(G952), .A2(n480), .ZN(n728) );
  NOR2_X1 U595 ( .A1(G953), .A2(n728), .ZN(n543) );
  AND2_X1 U596 ( .A1(G953), .A2(G902), .ZN(n479) );
  NAND2_X1 U597 ( .A1(n480), .A2(n479), .ZN(n540) );
  NOR2_X1 U598 ( .A1(G898), .A2(n540), .ZN(n481) );
  XOR2_X1 U599 ( .A(KEYINPUT93), .B(n481), .Z(n482) );
  NOR2_X1 U600 ( .A1(n543), .A2(n482), .ZN(n483) );
  XNOR2_X1 U601 ( .A(KEYINPUT67), .B(KEYINPUT0), .ZN(n484) );
  INV_X1 U602 ( .A(n589), .ZN(n515) );
  NAND2_X1 U603 ( .A1(n519), .A2(G210), .ZN(n487) );
  XOR2_X1 U604 ( .A(KEYINPUT74), .B(KEYINPUT96), .Z(n486) );
  XNOR2_X1 U605 ( .A(G137), .B(KEYINPUT5), .ZN(n488) );
  XNOR2_X1 U606 ( .A(n489), .B(n490), .ZN(n493) );
  XNOR2_X2 U607 ( .A(n494), .B(G472), .ZN(n605) );
  NAND2_X1 U608 ( .A1(G227), .A2(n768), .ZN(n497) );
  XNOR2_X1 U609 ( .A(KEYINPUT77), .B(n495), .ZN(n496) );
  NAND2_X1 U610 ( .A1(n682), .A2(n536), .ZN(n499) );
  NAND2_X1 U611 ( .A1(G221), .A2(n530), .ZN(n506) );
  NAND2_X1 U612 ( .A1(G234), .A2(n643), .ZN(n508) );
  XNOR2_X1 U613 ( .A(KEYINPUT20), .B(n508), .ZN(n511) );
  XNOR2_X1 U614 ( .A(KEYINPUT25), .B(n459), .ZN(n509) );
  AND2_X1 U615 ( .A1(n511), .A2(G221), .ZN(n512) );
  XNOR2_X1 U616 ( .A(n512), .B(KEYINPUT21), .ZN(n694) );
  AND2_X1 U617 ( .A1(n579), .A2(n694), .ZN(n699) );
  INV_X1 U618 ( .A(n612), .ZN(n513) );
  NAND2_X1 U619 ( .A1(n697), .A2(n513), .ZN(n514) );
  XNOR2_X1 U620 ( .A(G143), .B(G131), .ZN(n516) );
  XOR2_X1 U621 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n518) );
  XNOR2_X1 U622 ( .A(G104), .B(KEYINPUT98), .ZN(n517) );
  NAND2_X1 U623 ( .A1(G214), .A2(n519), .ZN(n520) );
  XNOR2_X1 U624 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n523) );
  INV_X1 U625 ( .A(G475), .ZN(n522) );
  XNOR2_X1 U626 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U627 ( .A(n351), .B(n529), .ZN(n535) );
  AND2_X1 U628 ( .A1(G217), .A2(n530), .ZN(n533) );
  AND2_X1 U629 ( .A1(n674), .A2(n536), .ZN(n538) );
  INV_X1 U630 ( .A(G478), .ZN(n537) );
  XNOR2_X1 U631 ( .A(n538), .B(n537), .ZN(n592) );
  INV_X1 U632 ( .A(n592), .ZN(n562) );
  NAND2_X1 U633 ( .A1(n736), .A2(n743), .ZN(n539) );
  XNOR2_X1 U634 ( .A(n539), .B(G104), .ZN(G6) );
  XOR2_X1 U635 ( .A(KEYINPUT105), .B(n540), .Z(n541) );
  NOR2_X1 U636 ( .A1(G900), .A2(n541), .ZN(n542) );
  NOR2_X1 U637 ( .A1(n543), .A2(n542), .ZN(n608) );
  NAND2_X1 U638 ( .A1(n545), .A2(n544), .ZN(n553) );
  INV_X1 U639 ( .A(KEYINPUT109), .ZN(n547) );
  OR2_X1 U640 ( .A1(n549), .A2(n562), .ZN(n596) );
  INV_X1 U641 ( .A(n596), .ZN(n746) );
  NAND2_X1 U642 ( .A1(n665), .A2(n746), .ZN(n551) );
  XOR2_X1 U643 ( .A(G128), .B(KEYINPUT29), .Z(n550) );
  XNOR2_X1 U644 ( .A(n551), .B(n550), .ZN(G30) );
  INV_X1 U645 ( .A(KEYINPUT6), .ZN(n552) );
  XNOR2_X1 U646 ( .A(n554), .B(KEYINPUT106), .ZN(n555) );
  INV_X1 U647 ( .A(n391), .ZN(n556) );
  NAND2_X1 U648 ( .A1(n620), .A2(n556), .ZN(n558) );
  XOR2_X1 U649 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n557) );
  XNOR2_X1 U650 ( .A(n558), .B(n557), .ZN(n560) );
  INV_X1 U651 ( .A(n619), .ZN(n609) );
  NAND2_X1 U652 ( .A1(n560), .A2(n609), .ZN(n639) );
  XNOR2_X1 U653 ( .A(n639), .B(G140), .ZN(G42) );
  INV_X1 U654 ( .A(n591), .ZN(n561) );
  NAND2_X1 U655 ( .A1(n562), .A2(n561), .ZN(n715) );
  INV_X1 U656 ( .A(n694), .ZN(n563) );
  NOR2_X1 U657 ( .A1(n715), .A2(n563), .ZN(n564) );
  NAND2_X1 U658 ( .A1(n594), .A2(n564), .ZN(n565) );
  INV_X1 U659 ( .A(n577), .ZN(n570) );
  INV_X1 U660 ( .A(KEYINPUT89), .ZN(n566) );
  XNOR2_X1 U661 ( .A(n698), .B(n566), .ZN(n622) );
  INV_X1 U662 ( .A(n622), .ZN(n568) );
  XOR2_X1 U663 ( .A(KEYINPUT103), .B(n579), .Z(n693) );
  OR2_X1 U664 ( .A1(n588), .A2(n693), .ZN(n567) );
  NOR2_X1 U665 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U666 ( .A(G119), .B(n586), .Z(G21) );
  INV_X1 U667 ( .A(n713), .ZN(n571) );
  NOR2_X1 U668 ( .A1(n715), .A2(n571), .ZN(n573) );
  INV_X1 U669 ( .A(KEYINPUT38), .ZN(n572) );
  XNOR2_X1 U670 ( .A(n619), .B(n572), .ZN(n714) );
  NAND2_X1 U671 ( .A1(n573), .A2(n714), .ZN(n574) );
  XNOR2_X1 U672 ( .A(n574), .B(KEYINPUT41), .ZN(n729) );
  INV_X1 U673 ( .A(KEYINPUT42), .ZN(n575) );
  XNOR2_X1 U674 ( .A(n576), .B(n575), .ZN(n634) );
  XOR2_X1 U675 ( .A(G137), .B(n634), .Z(G39) );
  NAND2_X1 U676 ( .A1(n580), .A2(n697), .ZN(n578) );
  XOR2_X1 U677 ( .A(G110), .B(n587), .Z(G12) );
  INV_X1 U678 ( .A(n580), .ZN(n581) );
  XNOR2_X1 U679 ( .A(n583), .B(n582), .ZN(n584) );
  NAND2_X1 U680 ( .A1(n584), .A2(n693), .ZN(n585) );
  XNOR2_X1 U681 ( .A(n598), .B(G101), .ZN(G3) );
  NAND2_X1 U682 ( .A1(n592), .A2(n591), .ZN(n610) );
  NOR2_X1 U683 ( .A1(n593), .A2(n697), .ZN(n705) );
  NAND2_X1 U684 ( .A1(n705), .A2(n594), .ZN(n595) );
  NAND2_X1 U685 ( .A1(n396), .A2(n596), .ZN(n710) );
  XNOR2_X1 U686 ( .A(n710), .B(KEYINPUT83), .ZN(n601) );
  OR2_X1 U687 ( .A1(n601), .A2(KEYINPUT47), .ZN(n602) );
  INV_X1 U688 ( .A(KEYINPUT47), .ZN(n603) );
  OR2_X1 U689 ( .A1(n710), .A2(n603), .ZN(n604) );
  XNOR2_X1 U690 ( .A(n604), .B(KEYINPUT82), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n605), .A2(n713), .ZN(n606) );
  XNOR2_X1 U692 ( .A(KEYINPUT30), .B(n606), .ZN(n607) );
  NOR2_X1 U693 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n627), .A2(n611), .ZN(n613) );
  XNOR2_X1 U695 ( .A(n612), .B(KEYINPUT108), .ZN(n628) );
  OR2_X1 U696 ( .A1(n613), .A2(n628), .ZN(n741) );
  AND2_X1 U697 ( .A1(n614), .A2(n741), .ZN(n615) );
  NAND2_X1 U698 ( .A1(n616), .A2(n615), .ZN(n618) );
  INV_X1 U699 ( .A(KEYINPUT72), .ZN(n617) );
  XNOR2_X1 U700 ( .A(n618), .B(n617), .ZN(n625) );
  INV_X1 U701 ( .A(KEYINPUT36), .ZN(n621) );
  INV_X1 U702 ( .A(KEYINPUT86), .ZN(n623) );
  XNOR2_X1 U703 ( .A(n750), .B(n623), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U705 ( .A(n626), .B(KEYINPUT69), .ZN(n638) );
  NAND2_X1 U706 ( .A1(n627), .A2(n714), .ZN(n629) );
  OR2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n640), .A2(n743), .ZN(n633) );
  INV_X1 U709 ( .A(KEYINPUT110), .ZN(n631) );
  XNOR2_X1 U710 ( .A(n631), .B(KEYINPUT40), .ZN(n632) );
  XNOR2_X1 U711 ( .A(n633), .B(n632), .ZN(n775) );
  INV_X1 U712 ( .A(KEYINPUT46), .ZN(n635) );
  XNOR2_X1 U713 ( .A(n636), .B(n635), .ZN(n637) );
  AND2_X1 U714 ( .A1(n640), .A2(n746), .ZN(n752) );
  INV_X1 U715 ( .A(n752), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n668), .A2(G210), .ZN(n648) );
  XOR2_X1 U717 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n645) );
  XNOR2_X1 U718 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n648), .B(n647), .ZN(n650) );
  INV_X1 U720 ( .A(G952), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n649), .A2(G953), .ZN(n672) );
  NAND2_X1 U722 ( .A1(n650), .A2(n672), .ZN(n652) );
  XOR2_X1 U723 ( .A(KEYINPUT118), .B(KEYINPUT56), .Z(n651) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(G51) );
  NAND2_X1 U725 ( .A1(n668), .A2(G472), .ZN(n655) );
  XNOR2_X1 U726 ( .A(n653), .B(KEYINPUT62), .ZN(n654) );
  XNOR2_X1 U727 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U728 ( .A1(n656), .A2(n672), .ZN(n657) );
  XNOR2_X1 U729 ( .A(n657), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U730 ( .A1(n668), .A2(G475), .ZN(n661) );
  XNOR2_X1 U731 ( .A(KEYINPUT90), .B(KEYINPUT59), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n658), .B(n659), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n661), .B(n660), .ZN(n662) );
  NAND2_X1 U734 ( .A1(n662), .A2(n672), .ZN(n664) );
  INV_X1 U735 ( .A(KEYINPUT60), .ZN(n663) );
  XNOR2_X1 U736 ( .A(n664), .B(n663), .ZN(G60) );
  NAND2_X1 U737 ( .A1(n665), .A2(n743), .ZN(n666) );
  XNOR2_X1 U738 ( .A(n666), .B(G146), .ZN(G48) );
  XNOR2_X1 U739 ( .A(n667), .B(G122), .ZN(G24) );
  NAND2_X1 U740 ( .A1(n678), .A2(G217), .ZN(n671) );
  XOR2_X1 U741 ( .A(n669), .B(KEYINPUT122), .Z(n670) );
  XNOR2_X1 U742 ( .A(n671), .B(n670), .ZN(n673) );
  INV_X1 U743 ( .A(n672), .ZN(n685) );
  NOR2_X1 U744 ( .A1(n673), .A2(n685), .ZN(G66) );
  NAND2_X1 U745 ( .A1(n678), .A2(G478), .ZN(n676) );
  XNOR2_X1 U746 ( .A(n674), .B(KEYINPUT121), .ZN(n675) );
  XNOR2_X1 U747 ( .A(n676), .B(n675), .ZN(n677) );
  NOR2_X1 U748 ( .A1(n677), .A2(n685), .ZN(G63) );
  NAND2_X1 U749 ( .A1(n678), .A2(G469), .ZN(n684) );
  XOR2_X1 U750 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n680) );
  XNOR2_X1 U751 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n679) );
  XNOR2_X1 U752 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U753 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U754 ( .A(n684), .B(n683), .ZN(n686) );
  NOR2_X1 U755 ( .A1(n686), .A2(n685), .ZN(G54) );
  NOR2_X1 U756 ( .A1(n687), .A2(KEYINPUT2), .ZN(n688) );
  XNOR2_X1 U757 ( .A(n690), .B(KEYINPUT81), .ZN(n692) );
  NOR2_X1 U758 ( .A1(n692), .A2(n691), .ZN(n734) );
  NOR2_X1 U759 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U760 ( .A(n695), .B(KEYINPUT49), .ZN(n696) );
  NAND2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n702) );
  NOR2_X1 U762 ( .A1(n699), .A2(n391), .ZN(n700) );
  XNOR2_X1 U763 ( .A(n700), .B(KEYINPUT50), .ZN(n701) );
  NOR2_X1 U764 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U765 ( .A(n703), .B(KEYINPUT114), .ZN(n704) );
  NOR2_X1 U766 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U767 ( .A(n706), .B(KEYINPUT51), .ZN(n707) );
  XNOR2_X1 U768 ( .A(KEYINPUT115), .B(n707), .ZN(n709) );
  INV_X1 U769 ( .A(n729), .ZN(n708) );
  NOR2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n724) );
  NAND2_X1 U771 ( .A1(n710), .A2(n713), .ZN(n712) );
  INV_X1 U772 ( .A(n714), .ZN(n711) );
  NOR2_X1 U773 ( .A1(n712), .A2(n711), .ZN(n718) );
  NOR2_X1 U774 ( .A1(n714), .A2(n713), .ZN(n716) );
  NOR2_X1 U775 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U776 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U777 ( .A(n719), .B(KEYINPUT116), .ZN(n722) );
  INV_X1 U778 ( .A(n720), .ZN(n721) );
  NOR2_X1 U779 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U780 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U781 ( .A(n725), .B(KEYINPUT52), .ZN(n726) );
  XOR2_X1 U782 ( .A(KEYINPUT117), .B(n726), .Z(n727) );
  NOR2_X1 U783 ( .A1(n728), .A2(n727), .ZN(n732) );
  NAND2_X1 U784 ( .A1(n720), .A2(n729), .ZN(n730) );
  NAND2_X1 U785 ( .A1(n730), .A2(n768), .ZN(n731) );
  OR2_X1 U786 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U787 ( .A(n735), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U788 ( .A1(n736), .A2(n746), .ZN(n738) );
  XOR2_X1 U789 ( .A(KEYINPUT111), .B(KEYINPUT27), .Z(n737) );
  XNOR2_X1 U790 ( .A(n738), .B(n737), .ZN(n740) );
  XOR2_X1 U791 ( .A(G107), .B(KEYINPUT26), .Z(n739) );
  XNOR2_X1 U792 ( .A(n740), .B(n739), .ZN(G9) );
  INV_X1 U793 ( .A(n741), .ZN(n742) );
  XOR2_X1 U794 ( .A(G143), .B(n742), .Z(G45) );
  NAND2_X1 U795 ( .A1(n747), .A2(n743), .ZN(n744) );
  XNOR2_X1 U796 ( .A(n744), .B(KEYINPUT112), .ZN(n745) );
  XNOR2_X1 U797 ( .A(G113), .B(n745), .ZN(G15) );
  XOR2_X1 U798 ( .A(G116), .B(KEYINPUT113), .Z(n749) );
  NAND2_X1 U799 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U800 ( .A(n749), .B(n748), .ZN(G18) );
  XNOR2_X1 U801 ( .A(n750), .B(G125), .ZN(n751) );
  XNOR2_X1 U802 ( .A(n751), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U803 ( .A(G134), .B(n752), .Z(G36) );
  XNOR2_X1 U804 ( .A(n753), .B(KEYINPUT125), .ZN(n755) );
  NOR2_X1 U805 ( .A1(G898), .A2(n768), .ZN(n754) );
  NOR2_X1 U806 ( .A1(n755), .A2(n754), .ZN(n764) );
  NAND2_X1 U807 ( .A1(n442), .A2(n768), .ZN(n762) );
  XOR2_X1 U808 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n758) );
  NAND2_X1 U809 ( .A1(G224), .A2(G953), .ZN(n757) );
  XNOR2_X1 U810 ( .A(n758), .B(n757), .ZN(n759) );
  NAND2_X1 U811 ( .A1(G898), .A2(n759), .ZN(n760) );
  XNOR2_X1 U812 ( .A(n760), .B(KEYINPUT124), .ZN(n761) );
  NAND2_X1 U813 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U814 ( .A(n764), .B(n763), .ZN(G69) );
  XNOR2_X1 U815 ( .A(n766), .B(n765), .ZN(n770) );
  XNOR2_X1 U816 ( .A(n767), .B(n770), .ZN(n769) );
  NAND2_X1 U817 ( .A1(n769), .A2(n768), .ZN(n774) );
  XNOR2_X1 U818 ( .A(G227), .B(n770), .ZN(n771) );
  NAND2_X1 U819 ( .A1(n771), .A2(G900), .ZN(n772) );
  NAND2_X1 U820 ( .A1(n772), .A2(G953), .ZN(n773) );
  NAND2_X1 U821 ( .A1(n774), .A2(n773), .ZN(G72) );
  XNOR2_X1 U822 ( .A(G131), .B(n775), .ZN(n776) );
  XNOR2_X1 U823 ( .A(n776), .B(KEYINPUT127), .ZN(G33) );
endmodule

