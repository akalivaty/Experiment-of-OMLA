//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT64), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT1), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT66), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n219));
  AND3_X1   g0019(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  AOI21_X1  g0022(.A(new_n208), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n207), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n201), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n214), .B1(new_n215), .B2(new_n223), .C1(new_n226), .C2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n223), .A2(new_n215), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT67), .Z(new_n231));
  NOR2_X1   g0031(.A1(new_n229), .A2(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT68), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT69), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(G222), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G223), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n256), .B1(new_n257), .B2(new_n254), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  AND2_X1   g0063(.A1(G1), .A2(G13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G226), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n261), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G179), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n224), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n206), .A2(G20), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G50), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(G50), .B2(new_n278), .ZN(new_n285));
  INV_X1    g0085(.A(new_n281), .ZN(new_n286));
  XOR2_X1   g0086(.A(KEYINPUT8), .B(G58), .Z(new_n287));
  NAND2_X1  g0087(.A1(new_n207), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT70), .ZN(new_n289));
  OR3_X1    g0089(.A1(new_n251), .A2(KEYINPUT70), .A3(G20), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n286), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n285), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n295), .B1(new_n274), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n277), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  XOR2_X1   g0099(.A(new_n295), .B(KEYINPUT9), .Z(new_n300));
  NAND2_X1  g0100(.A1(new_n275), .A2(G190), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n274), .A2(G200), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n300), .A2(new_n305), .A3(new_n301), .A4(new_n302), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n299), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT71), .ZN(new_n308));
  INV_X1    g0108(.A(G244), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n261), .A2(new_n268), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n254), .A2(G232), .A3(new_n255), .ZN(new_n311));
  INV_X1    g0111(.A(G107), .ZN(new_n312));
  INV_X1    g0112(.A(G238), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n311), .B1(new_n312), .B2(new_n254), .C1(new_n258), .C2(new_n313), .ZN(new_n314));
  AOI211_X1 g0114(.A(new_n270), .B(new_n310), .C1(new_n314), .C2(new_n261), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n315), .A2(new_n276), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n282), .A2(G77), .A3(new_n283), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(G77), .B2(new_n278), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n287), .A2(new_n292), .B1(G20), .B2(G77), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT15), .B(G87), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n320), .A2(new_n288), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n286), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n315), .B2(G169), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n316), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n324), .B1(G190), .B2(new_n315), .ZN(new_n327));
  INV_X1    g0127(.A(G200), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(new_n315), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n307), .A2(new_n308), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n264), .A2(new_n265), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n271), .A2(new_n255), .ZN(new_n333));
  AND2_X1   g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  NOR2_X1   g0134(.A1(KEYINPUT3), .A2(G33), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n333), .B1(G232), .B2(new_n255), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G33), .A2(G97), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n332), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n332), .A2(G238), .A3(new_n267), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n269), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n339), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT13), .B1(new_n338), .B2(new_n342), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G200), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT72), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n290), .A2(new_n289), .A3(G77), .ZN(new_n350));
  INV_X1    g0150(.A(G68), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n292), .A2(G50), .B1(G20), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n286), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT11), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT12), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n356), .A2(KEYINPUT73), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(KEYINPUT73), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n357), .B(new_n358), .C1(G68), .C2(new_n278), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n359), .A2(KEYINPUT74), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n278), .A2(KEYINPUT12), .A3(G68), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n359), .B2(KEYINPUT74), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n354), .A2(new_n355), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n351), .B1(new_n206), .B2(G20), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n353), .A2(KEYINPUT11), .B1(new_n282), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(KEYINPUT75), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT75), .B1(new_n363), .B2(new_n365), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n367), .A2(new_n368), .B1(new_n369), .B2(new_n346), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n349), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT77), .B1(new_n367), .B2(new_n368), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n354), .A2(new_n355), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n360), .A2(new_n362), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n365), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT75), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT77), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n366), .A3(new_n378), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n372), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n346), .A2(G169), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n381), .A2(KEYINPUT14), .B1(new_n276), .B2(new_n346), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT76), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n296), .B1(new_n344), .B2(new_n345), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT14), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n382), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n346), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(G179), .B1(new_n384), .B2(new_n385), .ZN(new_n389));
  INV_X1    g0189(.A(new_n386), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT76), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n380), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n331), .A2(new_n371), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT8), .B(G58), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(new_n206), .B2(G20), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(new_n282), .B1(new_n279), .B2(new_n394), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n334), .A2(new_n335), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT7), .B1(new_n398), .B2(new_n207), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n253), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  AND2_X1   g0202(.A1(G58), .A2(G68), .ZN(new_n403));
  OAI21_X1  g0203(.A(G20), .B1(new_n403), .B2(new_n201), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n292), .A2(G159), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT16), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n286), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n402), .A2(KEYINPUT16), .A3(new_n407), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n397), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n271), .A2(G1698), .ZN(new_n413));
  OAI221_X1 g0213(.A(new_n413), .B1(G223), .B2(G1698), .C1(new_n334), .C2(new_n335), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G87), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n261), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n332), .A2(G232), .A3(new_n267), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n269), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n276), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n332), .B1(new_n414), .B2(new_n415), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n269), .A2(new_n418), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n296), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT18), .B1(new_n412), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n252), .A2(new_n207), .A3(new_n253), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT7), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n351), .B1(new_n428), .B2(new_n400), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n409), .B1(new_n429), .B2(new_n406), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(new_n411), .A3(new_n281), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n424), .B1(new_n431), .B2(new_n396), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n425), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n417), .A2(new_n369), .A3(new_n419), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n328), .B1(new_n421), .B2(new_n422), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n431), .A2(new_n396), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT17), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n431), .A2(new_n438), .A3(KEYINPUT17), .A4(new_n396), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(KEYINPUT78), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT78), .B1(new_n441), .B2(new_n442), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n435), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n308), .B1(new_n307), .B2(new_n330), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n393), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n278), .A2(G107), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT25), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n251), .A2(G1), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n279), .A2(new_n281), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n450), .B1(new_n453), .B2(new_n312), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n207), .B(G87), .C1(new_n334), .C2(new_n335), .ZN(new_n455));
  AND2_X1   g0255(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n456));
  NOR2_X1   g0256(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n254), .A2(new_n207), .A3(G87), .A4(new_n456), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G116), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G20), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT23), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n207), .B2(G107), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n312), .A2(KEYINPUT23), .A3(G20), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n459), .A2(new_n460), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT24), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT24), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n459), .A2(new_n460), .A3(new_n466), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n454), .B1(new_n471), .B2(new_n281), .ZN(new_n472));
  XOR2_X1   g0272(.A(new_n472), .B(KEYINPUT86), .Z(new_n473));
  OAI211_X1 g0273(.A(G257), .B(G1698), .C1(new_n334), .C2(new_n335), .ZN(new_n474));
  OAI211_X1 g0274(.A(G250), .B(new_n255), .C1(new_n334), .C2(new_n335), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G294), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n261), .ZN(new_n478));
  INV_X1    g0278(.A(G45), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(G1), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n261), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G264), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT87), .ZN(new_n485));
  INV_X1    g0285(.A(new_n266), .ZN(new_n486));
  AND2_X1   g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n480), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT87), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n478), .A2(new_n483), .A3(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n485), .A2(G179), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(G169), .B1(new_n484), .B2(new_n490), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n473), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n485), .A2(new_n491), .A3(new_n493), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n328), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n484), .A2(new_n490), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n369), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT88), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(new_n503), .A3(new_n472), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n498), .A2(new_n328), .B1(new_n369), .B2(new_n500), .ZN(new_n505));
  INV_X1    g0305(.A(new_n472), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT88), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n497), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT81), .ZN(new_n510));
  NOR2_X1   g0310(.A1(G238), .A2(G1698), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n309), .B2(G1698), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n254), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n332), .B1(new_n513), .B2(new_n461), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n206), .A2(G45), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n515), .A2(G250), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n332), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n486), .B2(new_n515), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n296), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n332), .A2(new_n516), .B1(new_n266), .B2(new_n480), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n512), .A2(new_n254), .B1(G33), .B2(G116), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n520), .B(new_n276), .C1(new_n332), .C2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n519), .B1(new_n522), .B2(KEYINPUT80), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(KEYINPUT80), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n510), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n207), .B(G68), .C1(new_n334), .C2(new_n335), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  INV_X1    g0328(.A(G97), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n288), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT82), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n531), .A2(new_n532), .A3(new_n207), .ZN(new_n533));
  INV_X1    g0333(.A(G87), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(new_n529), .A3(new_n312), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n532), .B1(new_n531), .B2(new_n207), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n527), .B(new_n530), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT83), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n286), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n527), .A2(new_n530), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n541), .B(KEYINPUT83), .C1(new_n537), .C2(new_n536), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n320), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(new_n278), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n452), .A2(new_n544), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OR2_X1    g0348(.A1(new_n522), .A2(KEYINPUT80), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n549), .A2(KEYINPUT81), .A3(new_n524), .A4(new_n519), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n526), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n453), .A2(new_n534), .ZN(new_n552));
  AOI211_X1 g0352(.A(new_n545), .B(new_n552), .C1(new_n540), .C2(new_n542), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n520), .B1(new_n521), .B2(new_n332), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n328), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(G190), .B2(new_n554), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G244), .B(new_n255), .C1(new_n334), .C2(new_n335), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT4), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n254), .A2(KEYINPUT4), .A3(G244), .A4(new_n255), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G33), .A2(G283), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n254), .A2(G250), .A3(G1698), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n560), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n564), .A2(new_n261), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT79), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n482), .A2(new_n566), .A3(G257), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n489), .A2(G257), .A3(new_n332), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT79), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n491), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n296), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n292), .A2(G77), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT6), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n573), .A2(new_n529), .A3(G107), .ZN(new_n574));
  XNOR2_X1  g0374(.A(G97), .B(G107), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n574), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n572), .B1(new_n576), .B2(new_n207), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n312), .B1(new_n428), .B2(new_n400), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n281), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n279), .A2(new_n529), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n452), .A2(G97), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n564), .A2(new_n261), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n490), .B1(KEYINPUT79), .B2(new_n568), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n583), .A2(new_n584), .A3(new_n276), .A4(new_n567), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n571), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(G200), .B1(new_n565), .B2(new_n570), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n581), .A2(new_n580), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n575), .A2(new_n573), .ZN(new_n589));
  INV_X1    g0389(.A(new_n574), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n591), .A2(G20), .B1(G77), .B2(new_n292), .ZN(new_n592));
  INV_X1    g0392(.A(new_n578), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n588), .B1(new_n594), .B2(new_n281), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n583), .A2(new_n584), .A3(G190), .A4(new_n567), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n587), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n551), .A2(new_n557), .A3(new_n586), .A4(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(G264), .B(G1698), .C1(new_n334), .C2(new_n335), .ZN(new_n599));
  OAI211_X1 g0399(.A(G257), .B(new_n255), .C1(new_n334), .C2(new_n335), .ZN(new_n600));
  INV_X1    g0400(.A(G303), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n599), .B(new_n600), .C1(new_n601), .C2(new_n254), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n261), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT84), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n482), .B2(G270), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n489), .A2(G270), .A3(new_n332), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(KEYINPUT84), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n491), .B(new_n603), .C1(new_n605), .C2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n562), .B(new_n207), .C1(G33), .C2(new_n529), .ZN(new_n609));
  INV_X1    g0409(.A(G116), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(G20), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n281), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT20), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n609), .A2(KEYINPUT20), .A3(new_n281), .A4(new_n611), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n278), .A2(G116), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n452), .B2(G116), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n296), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n608), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT21), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n608), .A2(KEYINPUT21), .A3(new_n619), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n482), .A2(new_n604), .A3(G270), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n606), .A2(KEYINPUT84), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n490), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n616), .A2(new_n618), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n626), .A2(new_n627), .A3(G179), .A4(new_n603), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n622), .A2(new_n623), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n627), .B1(new_n608), .B2(G200), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n369), .B2(new_n608), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n598), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n448), .A2(new_n509), .A3(new_n633), .ZN(G372));
  NOR2_X1   g0434(.A1(new_n349), .A2(new_n370), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n392), .B1(new_n326), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT90), .ZN(new_n637));
  OAI22_X1  g0437(.A1(new_n636), .A2(new_n637), .B1(new_n445), .B2(new_n444), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n435), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n304), .A2(new_n306), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n299), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n448), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n586), .A2(KEYINPUT89), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n519), .A2(new_n522), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n553), .A2(new_n556), .B1(new_n548), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT89), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n571), .A2(new_n582), .A3(new_n647), .A4(new_n585), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n644), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n586), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n551), .A2(KEYINPUT26), .A3(new_n557), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n496), .A2(new_n506), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n629), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n548), .A2(new_n645), .ZN(new_n657));
  AND4_X1   g0457(.A1(new_n557), .A2(new_n597), .A3(new_n586), .A4(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n503), .B1(new_n502), .B2(new_n472), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n505), .A2(KEYINPUT88), .A3(new_n506), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n656), .B(new_n658), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n654), .A2(new_n661), .A3(new_n657), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n642), .B1(new_n643), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g0464(.A(new_n664), .B(KEYINPUT91), .Z(G369));
  NAND3_X1  g0465(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT92), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT27), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(G213), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G343), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n473), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n509), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n473), .A2(new_n496), .A3(new_n674), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT94), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n673), .B1(new_n616), .B2(new_n618), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n632), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n622), .A2(new_n623), .A3(new_n628), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT93), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT93), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n681), .A2(new_n686), .A3(new_n683), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n679), .B1(new_n688), .B2(G330), .ZN(new_n689));
  INV_X1    g0489(.A(G330), .ZN(new_n690));
  AOI211_X1 g0490(.A(KEYINPUT94), .B(new_n690), .C1(new_n685), .C2(new_n687), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n678), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n629), .A2(new_n674), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n472), .B1(new_n495), .B2(new_n494), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n509), .A2(new_n693), .B1(new_n694), .B2(new_n673), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(G399));
  NOR2_X1   g0496(.A1(new_n210), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n535), .A2(G116), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G1), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n228), .B2(new_n698), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT29), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n497), .A2(new_n629), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(new_n508), .A3(new_n658), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n551), .A2(new_n557), .A3(new_n652), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n650), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n707), .A2(KEYINPUT96), .B1(new_n650), .B2(new_n649), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n707), .A2(KEYINPUT96), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n657), .B(new_n705), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n703), .B1(new_n710), .B2(new_n673), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n662), .A2(new_n673), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n633), .A2(new_n497), .A3(new_n508), .A4(new_n673), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n583), .A2(new_n584), .A3(new_n567), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n554), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n485), .A2(new_n493), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT95), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n608), .B2(new_n276), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n626), .A2(KEYINPUT95), .A3(G179), .A4(new_n603), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n717), .A2(new_n718), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  AND4_X1   g0523(.A1(new_n276), .A2(new_n716), .A3(new_n608), .A4(new_n554), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n722), .A2(new_n723), .B1(new_n724), .B2(new_n498), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n717), .A2(new_n718), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(KEYINPUT30), .A3(new_n721), .A4(new_n720), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n673), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT31), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n715), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n728), .A2(KEYINPUT31), .ZN(new_n731));
  OAI21_X1  g0531(.A(G330), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n714), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n702), .B1(new_n734), .B2(G1), .ZN(G364));
  AOI21_X1  g0535(.A(new_n224), .B1(G20), .B2(new_n296), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n207), .A2(new_n276), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G200), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G190), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n207), .A2(G179), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(new_n369), .A3(G200), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n739), .A2(G68), .B1(new_n742), .B2(G107), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G190), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G159), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n738), .A2(new_n369), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n743), .B1(KEYINPUT32), .B2(new_n747), .C1(new_n202), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n737), .A2(new_n744), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n254), .B1(new_n751), .B2(new_n257), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(KEYINPUT32), .B2(new_n747), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n740), .A2(G190), .A3(G200), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n369), .A2(G179), .A3(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n207), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n753), .B1(new_n534), .B2(new_n754), .C1(new_n529), .C2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n737), .A2(G190), .A3(new_n328), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT99), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n750), .B(new_n757), .C1(G58), .C2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G317), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(KEYINPUT33), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n762), .A2(KEYINPUT33), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n739), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G283), .ZN(new_n766));
  INV_X1    g0566(.A(G326), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n765), .B1(new_n766), .B2(new_n741), .C1(new_n767), .C2(new_n749), .ZN(new_n768));
  INV_X1    g0568(.A(new_n751), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G311), .A2(new_n769), .B1(new_n746), .B2(G329), .ZN(new_n770));
  INV_X1    g0570(.A(G322), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n770), .B(new_n398), .C1(new_n771), .C2(new_n758), .ZN(new_n772));
  INV_X1    g0572(.A(G294), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n756), .A2(new_n773), .B1(new_n754), .B2(new_n601), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n768), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n736), .B1(new_n761), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n736), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n248), .A2(G45), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n210), .A2(new_n254), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n228), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n783), .B1(new_n479), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n781), .B1(new_n786), .B2(KEYINPUT98), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(KEYINPUT98), .B2(new_n786), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n210), .A2(new_n398), .ZN(new_n789));
  NAND2_X1  g0589(.A1(G355), .A2(KEYINPUT97), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G355), .A2(KEYINPUT97), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n791), .A2(new_n792), .B1(G116), .B2(new_n211), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n780), .B1(new_n788), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n209), .A2(G20), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n206), .B1(new_n795), .B2(G45), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n698), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n776), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n688), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(new_n800), .B2(new_n779), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n689), .A2(new_n691), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n798), .B1(new_n800), .B2(new_n690), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  NOR2_X1   g0605(.A1(new_n736), .A2(new_n777), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n797), .B1(new_n257), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n736), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n254), .B1(new_n746), .B2(G311), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n809), .B1(new_n610), .B2(new_n751), .C1(new_n773), .C2(new_n758), .ZN(new_n810));
  INV_X1    g0610(.A(new_n754), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n811), .A2(G107), .B1(new_n742), .B2(G87), .ZN(new_n812));
  INV_X1    g0612(.A(new_n739), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n766), .B2(new_n813), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n749), .A2(new_n601), .B1(new_n529), .B2(new_n756), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n810), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n748), .A2(G137), .B1(new_n769), .B2(G159), .ZN(new_n817));
  INV_X1    g0617(.A(G150), .ZN(new_n818));
  INV_X1    g0618(.A(G143), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(new_n818), .B2(new_n813), .C1(new_n759), .C2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT34), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n254), .B1(new_n745), .B2(new_n822), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n202), .A2(new_n754), .B1(new_n741), .B2(new_n351), .ZN(new_n824));
  INV_X1    g0624(.A(new_n756), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n823), .B(new_n824), .C1(G58), .C2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n816), .B1(new_n821), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n326), .A2(new_n674), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n329), .B1(new_n323), .B2(new_n673), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n326), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n807), .B1(new_n808), .B2(new_n827), .C1(new_n833), .C2(new_n778), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n712), .A2(new_n832), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT100), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n330), .A2(new_n673), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n682), .A2(new_n694), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n557), .A2(new_n597), .A3(new_n586), .A4(new_n657), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n840), .A2(new_n508), .B1(new_n548), .B2(new_n645), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n836), .B(new_n837), .C1(new_n841), .C2(new_n654), .ZN(new_n842));
  INV_X1    g0642(.A(new_n837), .ZN(new_n843));
  AOI21_X1  g0643(.A(KEYINPUT100), .B1(new_n662), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n835), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n798), .B1(new_n845), .B2(new_n732), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n845), .A2(new_n732), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n834), .B1(new_n847), .B2(new_n848), .ZN(G384));
  NOR2_X1   g0649(.A1(new_n795), .A2(new_n206), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n829), .B1(new_n842), .B2(new_n844), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n380), .A2(new_n674), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n392), .A2(new_n371), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n383), .B1(new_n382), .B2(new_n386), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT76), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n380), .B(new_n674), .C1(new_n856), .C2(new_n635), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n432), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n431), .A2(new_n396), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n672), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n859), .A2(new_n861), .A3(new_n439), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n859), .A2(new_n861), .A3(new_n864), .A4(new_n439), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n425), .A2(new_n434), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n441), .A2(new_n442), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT78), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n867), .B1(new_n870), .B2(new_n443), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n866), .B1(new_n871), .B2(new_n861), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(KEYINPUT38), .B(new_n866), .C1(new_n871), .C2(new_n861), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n851), .A2(new_n858), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n435), .A2(new_n672), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n875), .A2(KEYINPUT103), .ZN(new_n881));
  INV_X1    g0681(.A(new_n861), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n446), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT103), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT38), .A4(new_n866), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n425), .A2(new_n434), .A3(new_n441), .A4(new_n442), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n882), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n866), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT102), .B1(new_n889), .B2(new_n873), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT102), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n891), .B(KEYINPUT38), .C1(new_n866), .C2(new_n888), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT39), .B1(new_n886), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n392), .A2(new_n674), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n876), .A2(new_n897), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n894), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT104), .B1(new_n880), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n886), .A2(new_n893), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n897), .ZN(new_n902));
  INV_X1    g0702(.A(new_n898), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(new_n895), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT104), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n904), .A2(new_n905), .A3(new_n877), .A4(new_n879), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n448), .B1(new_n711), .B2(new_n713), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n642), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n907), .B(new_n909), .Z(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT31), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT105), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n912), .B1(new_n728), .B2(new_n913), .ZN(new_n914));
  AOI211_X1 g0714(.A(KEYINPUT105), .B(new_n673), .C1(new_n725), .C2(new_n727), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n729), .B(new_n715), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n832), .B1(new_n853), .B2(new_n857), .ZN(new_n917));
  AND4_X1   g0717(.A1(new_n911), .A2(new_n876), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n901), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n918), .B1(new_n920), .B2(KEYINPUT40), .ZN(new_n921));
  INV_X1    g0721(.A(new_n916), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n921), .B1(new_n643), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n911), .B1(new_n919), .B2(new_n901), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n448), .B(new_n916), .C1(new_n924), .C2(new_n918), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n923), .A2(G330), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n850), .B1(new_n910), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n926), .B2(new_n910), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT35), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n610), .B(new_n226), .C1(new_n576), .C2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n931), .A2(KEYINPUT101), .B1(KEYINPUT35), .B2(new_n591), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(KEYINPUT101), .B2(new_n931), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT36), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n228), .A2(new_n257), .A3(new_n403), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n351), .A2(G50), .ZN(new_n936));
  OAI211_X1 g0736(.A(G1), .B(new_n209), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n928), .A2(new_n934), .A3(new_n937), .ZN(G367));
  INV_X1    g0738(.A(G159), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n813), .A2(new_n939), .B1(new_n741), .B2(new_n257), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(G143), .B2(new_n748), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n254), .B1(new_n758), .B2(new_n818), .ZN(new_n942));
  INV_X1    g0742(.A(G137), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n751), .A2(new_n202), .B1(new_n745), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n756), .A2(new_n351), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(G58), .B2(new_n811), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n941), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n398), .B1(new_n745), .B2(new_n762), .C1(new_n766), .C2(new_n751), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n760), .B2(G303), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT46), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n754), .B2(new_n610), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n811), .A2(KEYINPUT46), .A3(G116), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n739), .A2(G294), .B1(new_n742), .B2(G97), .ZN(new_n955));
  INV_X1    g0755(.A(G311), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n955), .B1(new_n312), .B2(new_n756), .C1(new_n956), .C2(new_n749), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n948), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT107), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT47), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n736), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n646), .B1(new_n553), .B2(new_n673), .ZN(new_n962));
  OR3_X1    g0762(.A1(new_n657), .A2(new_n553), .A3(new_n673), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n962), .A2(new_n963), .A3(new_n779), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n236), .A2(new_n783), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n736), .B(new_n779), .C1(new_n210), .C2(new_n544), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n797), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n961), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n796), .B(KEYINPUT106), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n509), .A2(new_n693), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n678), .A2(new_n693), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n802), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n971), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n691), .B2(new_n689), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n678), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n688), .A2(G330), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT94), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n688), .A2(new_n679), .A3(G330), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT45), .ZN(new_n983));
  INV_X1    g0783(.A(new_n695), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n652), .A2(new_n674), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n597), .B(new_n586), .C1(new_n595), .C2(new_n673), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n983), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n695), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n984), .A2(KEYINPUT44), .A3(new_n988), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT44), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n695), .B2(new_n987), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n982), .A2(new_n996), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n990), .A2(new_n989), .B1(new_n992), .B2(new_n994), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n692), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n734), .B1(new_n977), .B2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n697), .B(KEYINPUT41), .Z(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n970), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n509), .A2(new_n693), .A3(new_n987), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n586), .B1(new_n497), .B2(new_n986), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n1005), .A2(KEYINPUT42), .B1(new_n673), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(KEYINPUT42), .B2(new_n1005), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n962), .A2(new_n963), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(KEYINPUT43), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1009), .A2(KEYINPUT43), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n1008), .A2(KEYINPUT43), .A3(new_n1009), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n692), .A2(new_n988), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n968), .B1(new_n1004), .B2(new_n1017), .ZN(G387));
  NAND2_X1  g0818(.A1(new_n977), .A2(new_n733), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n976), .A2(new_n734), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(new_n697), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n699), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n789), .A2(new_n1022), .B1(new_n312), .B2(new_n210), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n240), .A2(new_n479), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n287), .A2(new_n202), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT50), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n699), .B(new_n479), .C1(new_n351), .C2(new_n257), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n782), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1023), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n797), .B1(new_n1029), .B2(new_n780), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n811), .A2(G77), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n320), .B2(new_n756), .C1(new_n749), .C2(new_n939), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n398), .B1(new_n746), .B2(G150), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n202), .B2(new_n758), .C1(new_n351), .C2(new_n751), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n813), .A2(new_n394), .B1(new_n529), .B2(new_n741), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n741), .A2(new_n610), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n398), .B1(new_n745), .B2(new_n767), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n739), .A2(G311), .B1(new_n769), .B2(G303), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n771), .B2(new_n749), .C1(new_n759), .C2(new_n762), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n825), .A2(G283), .B1(new_n811), .B2(G294), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1037), .B(new_n1038), .C1(new_n1046), .C2(KEYINPUT49), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(KEYINPUT49), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1036), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1030), .B1(new_n1049), .B2(new_n808), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n978), .B2(new_n779), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n976), .B2(new_n970), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1021), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(G393));
  INV_X1    g0854(.A(new_n1020), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1000), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n698), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT108), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1000), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n997), .A2(new_n999), .A3(KEYINPUT108), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1060), .A2(new_n970), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT110), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n245), .A2(new_n782), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n780), .B1(new_n529), .B2(new_n211), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n798), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n749), .A2(new_n818), .B1(new_n939), .B2(new_n758), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n254), .B1(new_n745), .B2(new_n819), .C1(new_n394), .C2(new_n751), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n739), .A2(G50), .B1(new_n742), .B2(G87), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n756), .A2(new_n257), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G68), .B2(new_n811), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT109), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n749), .A2(new_n762), .B1(new_n956), .B2(new_n758), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT52), .Z(new_n1077));
  OAI221_X1 g0877(.A(new_n398), .B1(new_n745), .B2(new_n771), .C1(new_n773), .C2(new_n751), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n813), .A2(new_n601), .B1(new_n741), .B2(new_n312), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n756), .A2(new_n610), .B1(new_n754), .B2(new_n766), .ZN(new_n1080));
  OR4_X1    g0880(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1074), .A2(KEYINPUT109), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1075), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1066), .B1(new_n1083), .B2(new_n736), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n779), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1084), .B1(new_n987), .B2(new_n1085), .ZN(new_n1086));
  AND3_X1   g0886(.A1(new_n1062), .A2(new_n1063), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1063), .B1(new_n1062), .B2(new_n1086), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1058), .B1(new_n1087), .B2(new_n1088), .ZN(G390));
  NAND3_X1  g0889(.A1(new_n710), .A2(new_n673), .A3(new_n831), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n829), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n858), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n863), .A2(new_n865), .B1(new_n887), .B2(new_n882), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n891), .B1(new_n1093), .B2(KEYINPUT38), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n889), .A2(KEYINPUT102), .A3(new_n873), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n881), .B2(new_n885), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1097), .A2(new_n895), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1092), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n858), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n732), .A2(new_n832), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n895), .B1(new_n851), .B2(new_n858), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT111), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1103), .A2(new_n1104), .B1(new_n894), .B2(new_n898), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n662), .A2(new_n843), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n836), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n662), .A2(KEYINPUT100), .A3(new_n843), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n828), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n896), .B1(new_n1109), .B2(new_n1100), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1110), .A2(KEYINPUT111), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1099), .B(new_n1102), .C1(new_n1105), .C2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n894), .A2(new_n898), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n1110), .B2(KEYINPUT111), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1114), .A2(new_n1115), .B1(new_n1092), .B2(new_n1098), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n916), .A2(G330), .A3(new_n917), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT112), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT112), .A4(G330), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1112), .B(new_n970), .C1(new_n1116), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n806), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n798), .B1(new_n287), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1072), .B1(G283), .B2(new_n748), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n312), .B2(new_n813), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n254), .B1(new_n769), .B2(G97), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1127), .B1(new_n610), .B2(new_n758), .C1(new_n773), .C2(new_n745), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n351), .A2(new_n741), .B1(new_n754), .B2(new_n534), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1126), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT114), .Z(new_n1131));
  OAI22_X1  g0931(.A1(new_n813), .A2(new_n943), .B1(new_n741), .B2(new_n202), .ZN(new_n1132));
  INV_X1    g0932(.A(G128), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n749), .A2(new_n1133), .B1(new_n939), .B2(new_n756), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n758), .A2(new_n822), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n254), .B1(new_n751), .B2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1136), .B(new_n1138), .C1(G125), .C2(new_n746), .ZN(new_n1139));
  OR3_X1    g0939(.A1(new_n754), .A2(KEYINPUT53), .A3(new_n818), .ZN(new_n1140));
  OAI21_X1  g0940(.A(KEYINPUT53), .B1(new_n754), .B2(new_n818), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1135), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT115), .B1(new_n1131), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1143), .A2(new_n808), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1131), .A2(KEYINPUT115), .A3(new_n1142), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1124), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n1113), .B2(new_n778), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1122), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1112), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n448), .A2(G330), .A3(new_n916), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n642), .A2(new_n908), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT113), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n916), .A2(new_n1152), .A3(G330), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n833), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1152), .B1(new_n916), .B2(G330), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1100), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1101), .A2(new_n1091), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1100), .B1(new_n732), .B2(new_n832), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1119), .A2(new_n1159), .A3(new_n1120), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n851), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1151), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n698), .B1(new_n1149), .B2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1112), .B(new_n1162), .C1(new_n1116), .C2(new_n1121), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1148), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(G378));
  INV_X1    g0967(.A(KEYINPUT118), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n641), .A2(new_n298), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n295), .A2(new_n671), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1170), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n307), .A2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1171), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1174), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1168), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1174), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(new_n1175), .A3(KEYINPUT118), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(G330), .C1(new_n924), .C2(new_n918), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n916), .A2(new_n917), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT40), .B1(new_n1097), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n919), .A2(new_n911), .A3(new_n876), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n690), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1184), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n907), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1189), .B1(new_n921), .B2(new_n690), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1193), .A2(new_n900), .A3(new_n906), .A4(new_n1184), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1192), .A2(KEYINPUT119), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT119), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1151), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1165), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT57), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1192), .A2(KEYINPUT57), .A3(new_n1194), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n697), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n797), .B1(new_n202), .B2(new_n806), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n742), .A2(G58), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n254), .A2(G41), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n746), .A2(G283), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1031), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT116), .Z(new_n1210));
  OAI22_X1  g1010(.A1(new_n758), .A2(new_n312), .B1(new_n751), .B2(new_n320), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n529), .A2(new_n813), .B1(new_n749), .B2(new_n610), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(new_n1210), .A2(new_n946), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n1213), .A2(KEYINPUT58), .B1(new_n1207), .B2(new_n1214), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G150), .A2(new_n825), .B1(new_n748), .B2(G125), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT117), .Z(new_n1217));
  NAND2_X1  g1017(.A1(new_n769), .A2(G137), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n1133), .B2(new_n758), .C1(new_n754), .C2(new_n1137), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G132), .B2(new_n739), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1217), .A2(new_n1220), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1223));
  AOI211_X1 g1023(.A(G33), .B(G41), .C1(new_n746), .C2(G124), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n939), .B2(new_n741), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1222), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1215), .B(new_n1226), .C1(KEYINPUT58), .C2(new_n1213), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1205), .B1(new_n808), .B2(new_n1227), .C1(new_n1183), .C2(new_n778), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1197), .B2(new_n970), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1204), .A2(new_n1230), .ZN(G375));
  NAND3_X1  g1031(.A1(new_n1158), .A2(new_n1161), .A3(new_n1151), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1163), .A2(new_n1003), .A3(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n969), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1100), .A2(new_n777), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n798), .B1(G68), .B2(new_n1123), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n748), .A2(G132), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT121), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n254), .B1(new_n751), .B2(new_n818), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G128), .B2(new_n746), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1238), .B(new_n1240), .C1(new_n943), .C2(new_n759), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n811), .A2(G159), .B1(new_n742), .B2(G58), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1242), .B1(new_n202), .B2(new_n756), .C1(new_n813), .C2(new_n1137), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n398), .B1(new_n741), .B2(new_n257), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT120), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n758), .A2(new_n766), .B1(new_n745), .B2(new_n601), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G107), .B2(new_n769), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n825), .A2(new_n544), .B1(new_n811), .B2(G97), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G116), .A2(new_n739), .B1(new_n748), .B2(G294), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n1241), .A2(new_n1243), .B1(new_n1245), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1236), .B1(new_n1251), .B2(new_n736), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1234), .B1(new_n1235), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1233), .A2(new_n1253), .ZN(G381));
  OR2_X1    g1054(.A1(G375), .A2(KEYINPUT122), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G375), .A2(KEYINPUT122), .ZN(new_n1256));
  INV_X1    g1056(.A(G387), .ZN(new_n1257));
  INV_X1    g1057(.A(G384), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1021), .A2(new_n804), .A3(new_n1052), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NOR4_X1   g1060(.A1(new_n1260), .A2(G378), .A3(G390), .A4(G381), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1255), .A2(new_n1256), .A3(new_n1261), .ZN(G407));
  INV_X1    g1062(.A(G213), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1263), .A2(G343), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1255), .A2(new_n1166), .A3(new_n1256), .A4(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1066(.A(KEYINPUT62), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT60), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1232), .B1(new_n1162), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT123), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT123), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1271), .B(new_n1232), .C1(new_n1162), .C2(new_n1268), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1232), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n698), .B1(new_n1273), .B2(KEYINPUT60), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1270), .A2(new_n1272), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1253), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1258), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(G384), .A3(new_n1253), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  OAI211_X1 g1079(.A(G378), .B(new_n1230), .C1(new_n1200), .C2(new_n1203), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1196), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1192), .A2(new_n1194), .A3(KEYINPUT119), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1199), .A3(new_n1003), .A4(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1192), .A2(new_n1194), .A3(new_n970), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(new_n1228), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1166), .ZN(new_n1286));
  AOI211_X1 g1086(.A(new_n1264), .B(new_n1279), .C1(new_n1280), .C2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT124), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1267), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1280), .A2(new_n1286), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1264), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1264), .A2(G2897), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1279), .B(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT61), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1279), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1290), .A2(new_n1291), .A3(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1297), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1289), .A2(new_n1295), .A3(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT125), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G390), .A2(new_n1257), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1062), .A2(new_n1086), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(KEYINPUT110), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1062), .A2(new_n1063), .A3(new_n1086), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(G387), .A3(new_n1058), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1053), .A2(new_n804), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1307), .A2(new_n1259), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1301), .A2(new_n1306), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1301), .B2(new_n1306), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1300), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(G390), .A2(new_n1257), .ZN(new_n1312));
  AOI21_X1  g1112(.A(G387), .B1(new_n1305), .B2(new_n1058), .ZN(new_n1313));
  OAI22_X1  g1113(.A1(new_n1312), .A2(new_n1313), .B1(new_n1259), .B2(new_n1307), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1301), .A2(new_n1306), .A3(new_n1308), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1314), .A2(KEYINPUT125), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1311), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1299), .A2(new_n1317), .ZN(new_n1318));
  OR2_X1    g1118(.A1(new_n1287), .A2(KEYINPUT63), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1287), .A2(KEYINPUT63), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .A4(new_n1295), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1318), .A2(new_n1322), .ZN(G405));
  AOI21_X1  g1123(.A(G378), .B1(new_n1204), .B2(new_n1230), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT126), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1280), .A2(new_n1325), .ZN(new_n1326));
  OR2_X1    g1126(.A1(new_n1324), .A2(new_n1326), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1279), .A2(KEYINPUT127), .ZN(new_n1328));
  NOR3_X1   g1128(.A1(new_n1309), .A2(new_n1310), .A3(new_n1300), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT125), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1328), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1311), .B(new_n1316), .C1(KEYINPUT127), .C2(new_n1279), .ZN(new_n1332));
  AOI22_X1  g1132(.A1(new_n1324), .A2(KEYINPUT126), .B1(KEYINPUT127), .B2(new_n1279), .ZN(new_n1333));
  AND4_X1   g1133(.A1(new_n1327), .A2(new_n1331), .A3(new_n1332), .A4(new_n1333), .ZN(new_n1334));
  AOI22_X1  g1134(.A1(new_n1331), .A2(new_n1332), .B1(new_n1327), .B2(new_n1333), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(G402));
endmodule


