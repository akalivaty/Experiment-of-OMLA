//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  XNOR2_X1  g000(.A(G116), .B(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT5), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  OAI211_X1 g004(.A(new_n188), .B(G113), .C1(KEYINPUT5), .C2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G104), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT78), .A2(G107), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT78), .A2(G107), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n193), .B1(new_n196), .B2(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G101), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n192), .A2(G104), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT79), .A2(G101), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT79), .A2(G101), .ZN(new_n201));
  NOR3_X1   g015(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n195), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT3), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT78), .A2(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(KEYINPUT77), .B1(new_n193), .B2(KEYINPUT3), .ZN(new_n208));
  OAI211_X1 g022(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n204), .C2(G107), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n202), .B(new_n207), .C1(new_n208), .C2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n212));
  INV_X1    g026(.A(G113), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n215));
  NAND3_X1  g029(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n187), .B(new_n214), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n191), .A2(new_n198), .A3(new_n211), .A4(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G101), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT77), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n223), .A2(new_n209), .B1(new_n196), .B2(new_n205), .ZN(new_n224));
  INV_X1    g038(.A(new_n199), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n220), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n211), .A2(KEYINPUT4), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n225), .B(new_n207), .C1(new_n210), .C2(new_n208), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(G101), .ZN(new_n231));
  INV_X1    g045(.A(new_n187), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n217), .A2(new_n215), .ZN(new_n233));
  NOR2_X1   g047(.A1(KEYINPUT2), .A2(G113), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n218), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n219), .B1(new_n228), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G110), .B(G122), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n219), .B(new_n239), .C1(new_n228), .C2(new_n237), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(KEYINPUT6), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT6), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n238), .A2(new_n244), .A3(new_n240), .ZN(new_n245));
  INV_X1    g059(.A(G143), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(G146), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT64), .ZN(new_n248));
  INV_X1    g062(.A(G146), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(G143), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n246), .A2(KEYINPUT64), .A3(G146), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n247), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT0), .B(G128), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n249), .A2(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n246), .A2(G146), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  OAI22_X1  g071(.A1(new_n252), .A2(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G125), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n254), .A2(new_n255), .A3(new_n260), .A4(G128), .ZN(new_n261));
  INV_X1    g075(.A(G128), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n262), .B1(new_n254), .B2(KEYINPUT1), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n261), .B1(new_n252), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n259), .B1(G125), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G224), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(G953), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n265), .B(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n243), .A2(new_n245), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT7), .B1(new_n266), .B2(G953), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n239), .B(KEYINPUT8), .Z(new_n272));
  NAND2_X1  g086(.A1(new_n198), .A2(new_n211), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n191), .A2(new_n218), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n272), .B1(new_n275), .B2(new_n219), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n265), .A2(new_n270), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n271), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(G902), .B1(new_n278), .B2(new_n242), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n269), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(G210), .B1(G237), .B2(G902), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT84), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n269), .A2(new_n279), .A3(new_n281), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n269), .A2(new_n279), .A3(new_n281), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT84), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT95), .B(G952), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n289), .A2(G953), .ZN(new_n290));
  NAND2_X1  g104(.A1(G234), .A2(G237), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n291), .A2(G902), .A3(G953), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT21), .B(G898), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G214), .B1(G237), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n286), .A2(new_n288), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n246), .A2(G128), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n262), .A2(G143), .ZN(new_n302));
  INV_X1    g116(.A(G134), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  XOR2_X1   g119(.A(G116), .B(G122), .Z(new_n306));
  NAND2_X1  g120(.A1(new_n203), .A2(new_n206), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G116), .B(G122), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n196), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n305), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n262), .A2(G143), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n302), .B1(new_n312), .B2(KEYINPUT13), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT13), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n301), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G134), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n246), .A2(G128), .ZN(new_n317));
  OAI21_X1  g131(.A(G134), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n318), .A2(new_n304), .B1(new_n196), .B2(new_n309), .ZN(new_n319));
  INV_X1    g133(.A(G122), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(G116), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n192), .B1(new_n321), .B2(KEYINPUT14), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(new_n306), .B2(KEYINPUT14), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n311), .A2(new_n316), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT9), .B(G234), .ZN(new_n325));
  INV_X1    g139(.A(G217), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n325), .A2(new_n326), .A3(G953), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT94), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n308), .A2(new_n310), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n316), .A3(new_n304), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n319), .A2(new_n323), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT94), .ZN(new_n333));
  INV_X1    g147(.A(new_n327), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n330), .A2(new_n331), .A3(new_n327), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(KEYINPUT93), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT93), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(new_n324), .B2(new_n327), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n328), .B(new_n335), .C1(new_n337), .C2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G902), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G478), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(KEYINPUT15), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n344), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n340), .A2(new_n341), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT91), .ZN(new_n349));
  XOR2_X1   g163(.A(G113), .B(G122), .Z(new_n350));
  XOR2_X1   g164(.A(KEYINPUT90), .B(G104), .Z(new_n351));
  XOR2_X1   g165(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g166(.A(KEYINPUT89), .ZN(new_n353));
  INV_X1    g167(.A(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G125), .ZN(new_n355));
  INV_X1    g169(.A(G125), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G140), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n357), .A3(KEYINPUT72), .ZN(new_n358));
  OR3_X1    g172(.A1(new_n356), .A2(KEYINPUT72), .A3(G140), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT19), .ZN(new_n361));
  XNOR2_X1  g175(.A(G125), .B(G140), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(KEYINPUT19), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(G146), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n358), .A2(new_n359), .A3(KEYINPUT16), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT16), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n355), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n249), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n353), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G237), .A2(G953), .ZN(new_n371));
  AOI21_X1  g185(.A(G143), .B1(new_n371), .B2(G214), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(G143), .A3(G214), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(KEYINPUT66), .A2(G131), .ZN(new_n376));
  NOR2_X1   g190(.A1(KEYINPUT66), .A2(G131), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n373), .A2(new_n378), .A3(new_n374), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n369), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT19), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n384), .B1(new_n358), .B2(new_n359), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n249), .B1(new_n385), .B2(new_n363), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(KEYINPUT89), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n370), .A2(new_n382), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n358), .A2(new_n359), .A3(G146), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(new_n362), .B2(new_n249), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n358), .A2(new_n359), .A3(new_n390), .A4(G146), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT87), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT87), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(new_n396), .A3(new_n393), .ZN(new_n397));
  INV_X1    g211(.A(new_n374), .ZN(new_n398));
  NAND2_X1  g212(.A1(KEYINPUT18), .A2(G131), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT88), .B1(new_n399), .B2(KEYINPUT85), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n398), .A2(new_n372), .A3(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n373), .B(new_n374), .C1(KEYINPUT88), .C2(new_n399), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n401), .B1(new_n402), .B2(new_n400), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n395), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n352), .B1(new_n388), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT17), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n380), .A2(new_n406), .A3(new_n381), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n366), .A2(new_n249), .A3(new_n368), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n375), .A2(KEYINPUT17), .A3(new_n379), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n407), .A2(new_n383), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n404), .A2(new_n352), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n349), .B1(new_n405), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(G475), .A2(G902), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n405), .B2(new_n411), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT20), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n352), .B1(new_n404), .B2(new_n410), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n411), .A2(new_n417), .A3(KEYINPUT92), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n404), .A2(new_n410), .ZN(new_n419));
  INV_X1    g233(.A(new_n352), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(KEYINPUT92), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n341), .ZN(new_n422));
  OAI21_X1  g236(.A(G475), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  OAI221_X1 g237(.A(new_n413), .B1(new_n349), .B2(KEYINPUT20), .C1(new_n405), .C2(new_n411), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n416), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n300), .A2(new_n348), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G953), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G227), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT76), .ZN(new_n429));
  XNOR2_X1  g243(.A(G110), .B(G140), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n246), .A2(KEYINPUT64), .A3(G146), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT64), .B1(new_n246), .B2(G146), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n254), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n253), .ZN(new_n436));
  INV_X1    g250(.A(new_n256), .ZN(new_n437));
  INV_X1    g251(.A(new_n257), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n435), .A2(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n439), .B(new_n231), .C1(new_n226), .C2(new_n227), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT11), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n303), .B2(G137), .ZN(new_n442));
  INV_X1    g256(.A(G137), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(KEYINPUT11), .A3(G134), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n303), .A2(G137), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G131), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n378), .A2(new_n442), .A3(new_n444), .A4(new_n445), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT10), .ZN(new_n451));
  INV_X1    g265(.A(new_n261), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n247), .B2(new_n260), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n254), .A2(KEYINPUT80), .A3(KEYINPUT1), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(G128), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n452), .B1(new_n456), .B2(new_n256), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n451), .B1(new_n273), .B2(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n198), .A2(new_n211), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n264), .A2(KEYINPUT10), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n440), .A2(new_n450), .A3(new_n458), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT81), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n260), .B1(G143), .B2(new_n249), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n262), .B1(new_n464), .B2(KEYINPUT80), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n437), .B1(new_n465), .B2(new_n454), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n211), .B(new_n198), .C1(new_n466), .C2(new_n452), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n467), .A2(new_n451), .B1(new_n459), .B2(new_n460), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n450), .A4(new_n440), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n432), .B1(new_n463), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n450), .B1(new_n468), .B2(new_n440), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n463), .A2(new_n470), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT82), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n273), .A2(new_n457), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n264), .B1(new_n198), .B2(new_n211), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n449), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT12), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(KEYINPUT12), .B(new_n449), .C1(new_n477), .C2(new_n478), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n475), .A2(new_n476), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n432), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n463), .A2(new_n470), .B1(new_n482), .B2(new_n481), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(new_n476), .ZN(new_n487));
  OAI211_X1 g301(.A(G469), .B(new_n474), .C1(new_n485), .C2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G469), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n475), .A2(new_n483), .A3(new_n431), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n431), .B1(new_n475), .B2(new_n473), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n489), .B(new_n341), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n489), .A2(new_n341), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n488), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT83), .ZN(new_n496));
  OAI21_X1  g310(.A(G221), .B1(new_n325), .B2(G902), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n496), .B1(new_n495), .B2(new_n497), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n426), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT96), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n262), .A2(G119), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT23), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n262), .A2(KEYINPUT23), .A3(G119), .ZN(new_n505));
  INV_X1    g319(.A(G110), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n189), .A2(G128), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n504), .A2(new_n505), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n502), .A2(new_n507), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT24), .B(G110), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n508), .A2(new_n511), .B1(new_n249), .B2(new_n362), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n383), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n427), .A2(G221), .A3(G234), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT73), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT22), .B(G137), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n408), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(new_n369), .ZN(new_n519));
  INV_X1    g333(.A(new_n510), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n520), .A2(KEYINPUT70), .A3(new_n502), .A4(new_n507), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT70), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n509), .B2(new_n510), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n189), .A2(G128), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n507), .B(new_n505), .C1(new_n525), .C2(KEYINPUT23), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(KEYINPUT71), .A3(G110), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT71), .B1(new_n526), .B2(G110), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n524), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n513), .B(new_n517), .C1(new_n519), .C2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n526), .A2(G110), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT71), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n527), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n536), .B(new_n524), .C1(new_n518), .C2(new_n369), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n517), .B1(new_n537), .B2(new_n513), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n326), .B1(G234), .B2(new_n341), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(G902), .ZN(new_n541));
  XOR2_X1   g355(.A(new_n541), .B(KEYINPUT75), .Z(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n540), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n341), .B1(new_n532), .B2(new_n538), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT74), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT25), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT25), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n544), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n371), .A2(G210), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT27), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT26), .B(G101), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n439), .A2(new_n449), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n235), .A2(new_n218), .ZN(new_n559));
  INV_X1    g373(.A(new_n445), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n303), .A2(G137), .ZN(new_n561));
  OAI21_X1  g375(.A(G131), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n264), .A2(new_n448), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n558), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(KEYINPUT28), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n258), .A2(KEYINPUT65), .B1(new_n448), .B2(new_n447), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT65), .ZN(new_n567));
  OAI221_X1 g381(.A(new_n567), .B1(new_n256), .B2(new_n257), .C1(new_n252), .C2(new_n253), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n448), .A2(new_n562), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n566), .A2(new_n568), .B1(new_n264), .B2(new_n569), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n570), .A2(new_n559), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n557), .B1(new_n565), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n558), .A2(new_n563), .A3(KEYINPUT30), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n236), .B(new_n574), .C1(new_n570), .C2(KEYINPUT30), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT68), .B1(new_n564), .B2(new_n557), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n564), .A2(KEYINPUT68), .A3(new_n557), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n575), .B(KEYINPUT31), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT68), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n558), .A2(new_n559), .A3(new_n563), .ZN(new_n581));
  INV_X1    g395(.A(new_n557), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n564), .A2(KEYINPUT68), .A3(new_n557), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT31), .B1(new_n585), .B2(new_n575), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n573), .B1(new_n579), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT32), .ZN(new_n588));
  NOR2_X1   g402(.A1(G472), .A2(G902), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT31), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n577), .A2(new_n576), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n258), .A2(KEYINPUT65), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n568), .A3(new_n449), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT30), .B1(new_n594), .B2(new_n563), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n558), .A2(KEYINPUT30), .A3(new_n563), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n595), .A2(new_n559), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n591), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n572), .B1(new_n598), .B2(new_n578), .ZN(new_n599));
  INV_X1    g413(.A(new_n589), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT32), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n590), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n575), .A2(new_n564), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n582), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT29), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n565), .A2(new_n571), .A3(new_n557), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT69), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n559), .B1(new_n558), .B2(new_n563), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n608), .B(KEYINPUT28), .C1(new_n581), .C2(new_n609), .ZN(new_n610));
  OR2_X1    g424(.A1(new_n581), .A2(KEYINPUT28), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n558), .A2(new_n563), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n236), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n564), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n608), .B1(new_n615), .B2(KEYINPUT28), .ZN(new_n616));
  OR2_X1    g430(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n557), .A2(KEYINPUT29), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n607), .B(new_n341), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(G472), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n553), .B1(new_n602), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT96), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n426), .B(new_n622), .C1(new_n498), .C2(new_n499), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n501), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT97), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n200), .A2(new_n201), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G3));
  OR2_X1    g441(.A1(new_n498), .A2(new_n499), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n599), .A2(new_n600), .ZN(new_n629));
  INV_X1    g443(.A(G472), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n587), .B2(new_n341), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n553), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n298), .B1(new_n283), .B2(new_n285), .ZN(new_n634));
  INV_X1    g448(.A(new_n296), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n340), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n332), .A2(new_n334), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(KEYINPUT33), .A3(new_n336), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n343), .A2(G902), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n342), .A2(new_n343), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n425), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n636), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n633), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT34), .B(G104), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  OR2_X1    g463(.A1(new_n414), .A2(new_n415), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n414), .A2(new_n415), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n650), .A2(new_n348), .A3(new_n423), .A4(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n636), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n633), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT35), .B(G107), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  OAI21_X1  g470(.A(new_n513), .B1(new_n519), .B2(new_n530), .ZN(new_n657));
  INV_X1    g471(.A(new_n517), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(G902), .B1(new_n659), .B2(new_n531), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n549), .B1(new_n660), .B2(KEYINPUT74), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n551), .A3(new_n540), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n517), .A2(KEYINPUT36), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n657), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n542), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n667), .A2(new_n631), .A3(new_n629), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n501), .A2(new_n623), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT37), .B(G110), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT98), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n669), .B(new_n671), .ZN(G12));
  AOI22_X1  g486(.A1(new_n590), .A2(new_n601), .B1(new_n619), .B2(G472), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n281), .B1(new_n269), .B2(new_n279), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n297), .B1(new_n287), .B2(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n673), .A2(new_n675), .A3(new_n667), .ZN(new_n676));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n293), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n292), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n652), .A2(new_n680), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n676), .B(new_n681), .C1(new_n498), .C2(new_n499), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n679), .B(KEYINPUT39), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n628), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n685), .B1(new_n498), .B2(new_n499), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n287), .A2(new_n674), .A3(KEYINPUT84), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n285), .A2(new_n284), .ZN(new_n690));
  OAI21_X1  g504(.A(KEYINPUT38), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT38), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n286), .A2(new_n692), .A3(new_n288), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n615), .A2(new_n582), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n696), .B(KEYINPUT99), .Z(new_n697));
  NOR2_X1   g511(.A1(new_n592), .A2(new_n597), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n341), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(G472), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n602), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n425), .A2(new_n348), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n702), .A2(new_n298), .A3(new_n666), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n695), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n686), .A2(new_n688), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G143), .ZN(G45));
  AND3_X1   g520(.A1(new_n425), .A2(new_n644), .A3(new_n679), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n676), .B(new_n707), .C1(new_n498), .C2(new_n499), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  INV_X1    g523(.A(new_n621), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n489), .A2(KEYINPUT100), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n475), .A2(new_n473), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n712), .A2(new_n432), .B1(new_n471), .B2(new_n483), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n711), .B1(new_n713), .B2(G902), .ZN(new_n714));
  INV_X1    g528(.A(new_n711), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n341), .B(new_n715), .C1(new_n490), .C2(new_n491), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n497), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n646), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND2_X1  g535(.A1(new_n718), .A2(new_n653), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT101), .B(G116), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G18));
  AND3_X1   g538(.A1(new_n340), .A2(new_n341), .A3(new_n346), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n346), .B1(new_n340), .B2(new_n341), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AND4_X1   g541(.A1(new_n727), .A2(new_n416), .A3(new_n423), .A4(new_n424), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n283), .A2(new_n285), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n297), .A4(new_n635), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n717), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n673), .A2(new_n667), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  OAI21_X1  g548(.A(G472), .B1(new_n599), .B2(G902), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n582), .B1(new_n612), .B2(new_n616), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n736), .B1(new_n579), .B2(new_n586), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n589), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n552), .A2(new_n735), .A3(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n717), .A2(new_n739), .A3(new_n296), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT102), .B1(new_n702), .B2(new_n675), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT102), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n634), .A2(new_n742), .A3(new_n348), .A4(new_n425), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(KEYINPUT103), .B(G122), .Z(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G24));
  INV_X1    g561(.A(KEYINPUT104), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n735), .A2(new_n738), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n707), .A3(new_n666), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n634), .A2(new_n497), .A3(new_n714), .A4(new_n716), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n735), .A2(new_n666), .A3(new_n738), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n425), .A2(new_n644), .A3(new_n679), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n717), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n756), .A3(KEYINPUT104), .A4(new_n634), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G125), .ZN(G27));
  INV_X1    g573(.A(KEYINPUT106), .ZN(new_n760));
  INV_X1    g574(.A(new_n497), .ZN(new_n761));
  AOI211_X1 g575(.A(new_n761), .B(new_n298), .C1(new_n286), .C2(new_n288), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n488), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n712), .A2(new_n432), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n475), .A2(new_n483), .A3(new_n431), .ZN(new_n766));
  AOI21_X1  g580(.A(G902), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n493), .B1(new_n767), .B2(new_n489), .ZN(new_n768));
  AOI211_X1 g582(.A(new_n432), .B(new_n472), .C1(new_n470), .C2(new_n463), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n431), .B1(new_n486), .B2(new_n476), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n475), .A2(new_n483), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT82), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n769), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(KEYINPUT105), .A3(G469), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n764), .A2(new_n768), .A3(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n762), .A2(new_n775), .A3(new_n621), .A4(new_n707), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT42), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n760), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n762), .A2(new_n775), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n781), .A2(KEYINPUT42), .A3(new_n621), .A4(new_n707), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n776), .A2(new_n777), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(KEYINPUT106), .A3(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G131), .ZN(G33));
  NAND4_X1  g600(.A1(new_n762), .A2(new_n775), .A3(new_n621), .A4(new_n681), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G134), .ZN(G36));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n789), .B(new_n769), .C1(new_n770), .C2(new_n772), .ZN(new_n790));
  OAI21_X1  g604(.A(G469), .B1(new_n773), .B2(KEYINPUT45), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n790), .B1(new_n791), .B2(KEYINPUT107), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT107), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n793), .B(G469), .C1(new_n773), .C2(KEYINPUT45), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n493), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n492), .B1(new_n795), .B2(KEYINPUT46), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  AOI211_X1 g611(.A(new_n797), .B(new_n493), .C1(new_n792), .C2(new_n794), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n666), .B1(new_n631), .B2(new_n629), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n416), .A2(new_n423), .A3(new_n424), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT108), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n801), .B(new_n644), .C1(new_n802), .C2(KEYINPUT43), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n416), .A2(new_n423), .A3(new_n802), .A4(new_n424), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT43), .ZN(new_n805));
  INV_X1    g619(.A(new_n644), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n804), .B(new_n805), .C1(new_n425), .C2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n800), .B1(new_n803), .B2(new_n807), .ZN(new_n808));
  OR3_X1    g622(.A1(new_n808), .A2(KEYINPUT109), .A3(KEYINPUT44), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT109), .B1(new_n808), .B2(KEYINPUT44), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n297), .B1(new_n689), .B2(new_n690), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n808), .B2(KEYINPUT44), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n799), .A2(new_n813), .A3(new_n497), .A4(new_n685), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  OAI21_X1  g629(.A(new_n497), .B1(new_n796), .B2(new_n798), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT47), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(KEYINPUT47), .B(new_n497), .C1(new_n796), .C2(new_n798), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n673), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n821), .A2(new_n811), .A3(new_n552), .A4(new_n754), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G140), .ZN(G42));
  INV_X1    g638(.A(new_n716), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n472), .B1(new_n463), .B2(new_n470), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n766), .B1(new_n431), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n715), .B1(new_n827), .B2(new_n341), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  XOR2_X1   g643(.A(new_n829), .B(KEYINPUT110), .Z(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n761), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n818), .A2(new_n819), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n803), .A2(new_n807), .ZN(new_n833));
  INV_X1    g647(.A(new_n292), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n552), .A3(new_n834), .A4(new_n749), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n811), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n811), .A2(new_n717), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n834), .A3(new_n833), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n839), .A2(new_n753), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n701), .A2(new_n553), .A3(new_n292), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n838), .A3(new_n801), .A4(new_n806), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT50), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n829), .A2(new_n845), .A3(new_n497), .A4(new_n298), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT114), .B1(new_n717), .B2(new_n297), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n694), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n844), .B1(new_n848), .B2(new_n835), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n717), .A2(new_n297), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n850), .A2(new_n845), .B1(new_n691), .B2(new_n693), .ZN(new_n851));
  AOI211_X1 g665(.A(new_n292), .B(new_n739), .C1(new_n803), .C2(new_n807), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT50), .A4(new_n847), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n843), .A2(KEYINPUT51), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n837), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n841), .A2(new_n838), .ZN(new_n857));
  OAI221_X1 g671(.A(new_n290), .B1(new_n835), .B2(new_n751), .C1(new_n857), .C2(new_n645), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n839), .A2(new_n710), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n860), .A2(KEYINPUT48), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(KEYINPUT48), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n856), .A2(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n849), .A2(new_n853), .A3(KEYINPUT115), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT115), .B1(new_n849), .B2(new_n853), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n843), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n837), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(KEYINPUT116), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n867), .B1(new_n832), .B2(new_n836), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n872), .B1(new_n873), .B2(KEYINPUT51), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n864), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n666), .A2(new_n761), .A3(new_n680), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n744), .A2(new_n701), .A3(new_n775), .A4(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n758), .A2(new_n682), .A3(new_n708), .A4(new_n877), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT52), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n758), .A2(new_n682), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT52), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n348), .A2(new_n680), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(new_n423), .A3(new_n651), .A4(new_n650), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n673), .A2(new_n667), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n811), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n887), .B(new_n888), .C1(new_n498), .C2(new_n499), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n762), .A2(new_n775), .A3(new_n755), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n889), .A2(new_n787), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n780), .A2(new_n784), .A3(new_n891), .ZN(new_n892));
  AND4_X1   g706(.A1(new_n348), .A2(new_n416), .A3(new_n423), .A4(new_n424), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT111), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n893), .A2(new_n894), .B1(new_n425), .B2(new_n644), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT111), .B1(new_n425), .B2(new_n727), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n300), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n897), .B(new_n632), .C1(new_n498), .C2(new_n499), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n744), .A2(new_n740), .B1(new_n731), .B2(new_n732), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n621), .B(new_n756), .C1(new_n646), .C2(new_n653), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n624), .A2(new_n901), .A3(new_n669), .ZN(new_n902));
  NOR4_X1   g716(.A1(new_n879), .A2(new_n884), .A3(new_n892), .A4(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n892), .A2(new_n902), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT52), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n878), .B(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT53), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT54), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT112), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n892), .ZN(new_n911));
  INV_X1    g725(.A(new_n902), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n906), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n882), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n782), .A2(new_n783), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n881), .A2(new_n915), .A3(new_n891), .A4(KEYINPUT53), .ZN(new_n916));
  OR3_X1    g730(.A1(new_n879), .A2(new_n902), .A3(new_n916), .ZN(new_n917));
  XOR2_X1   g731(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n918));
  NAND3_X1  g732(.A1(new_n914), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(KEYINPUT112), .B(KEYINPUT54), .C1(new_n903), .C2(new_n907), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n875), .A2(new_n910), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  OR2_X1    g735(.A1(G952), .A2(G953), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n830), .B(KEYINPUT49), .Z(new_n924));
  NOR3_X1   g738(.A1(new_n553), .A2(new_n761), .A3(new_n298), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(new_n801), .A3(new_n644), .ZN(new_n926));
  OR4_X1    g740(.A1(new_n695), .A2(new_n924), .A3(new_n701), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n923), .A2(new_n927), .ZN(G75));
  NOR3_X1   g742(.A1(new_n879), .A2(new_n902), .A3(new_n916), .ZN(new_n929));
  OAI211_X1 g743(.A(G210), .B(G902), .C1(new_n907), .C2(new_n929), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n930), .A2(KEYINPUT117), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(KEYINPUT117), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n243), .A2(new_n245), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n268), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT55), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n935), .A2(KEYINPUT56), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n931), .A2(new_n932), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n427), .A2(G952), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT56), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n930), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n938), .B1(new_n940), .B2(new_n935), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n937), .A2(new_n941), .ZN(G51));
  XNOR2_X1  g756(.A(new_n493), .B(KEYINPUT57), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n918), .B1(new_n914), .B2(new_n917), .ZN(new_n944));
  INV_X1    g758(.A(new_n918), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n907), .A2(new_n929), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n943), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n827), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n341), .B1(new_n914), .B2(new_n917), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n792), .A2(new_n794), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT118), .Z(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n938), .B1(new_n948), .B2(new_n952), .ZN(G54));
  NAND2_X1  g767(.A1(KEYINPUT58), .A2(G475), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT119), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n949), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n405), .A2(new_n411), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n958), .A2(new_n959), .A3(new_n938), .ZN(G60));
  NAND2_X1  g774(.A1(new_n638), .A2(new_n640), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT120), .ZN(new_n962));
  NAND2_X1  g776(.A1(G478), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT59), .Z(new_n964));
  NOR2_X1   g778(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n944), .B2(new_n946), .ZN(new_n966));
  INV_X1    g780(.A(new_n938), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n964), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n914), .B1(new_n913), .B2(new_n884), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT112), .B1(new_n970), .B2(KEYINPUT54), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n920), .A2(new_n919), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n968), .B1(new_n973), .B2(new_n962), .ZN(G63));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT121), .Z(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT60), .Z(new_n977));
  OAI211_X1 g791(.A(new_n664), .B(new_n977), .C1(new_n907), .C2(new_n929), .ZN(new_n978));
  NOR2_X1   g792(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n938), .A2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n977), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n914), .B2(new_n917), .ZN(new_n982));
  INV_X1    g796(.A(new_n539), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n978), .B(new_n980), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT123), .Z(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n984), .B(new_n987), .ZN(G66));
  INV_X1    g802(.A(new_n294), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n427), .B1(new_n989), .B2(G224), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n990), .B1(new_n902), .B2(new_n427), .ZN(new_n991));
  INV_X1    g805(.A(G898), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n933), .B1(new_n992), .B2(G953), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n991), .B(new_n993), .ZN(G69));
  NOR2_X1   g808(.A1(new_n595), .A2(new_n596), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n361), .A2(new_n364), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n997), .B1(new_n677), .B2(new_n427), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n820), .A2(new_n822), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n744), .A2(new_n621), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n799), .A2(new_n497), .A3(new_n685), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n880), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n1002), .A2(new_n708), .A3(new_n787), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n814), .A2(new_n1001), .A3(new_n785), .A4(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n999), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n998), .B1(new_n1005), .B2(new_n427), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT62), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n686), .A2(new_n688), .A3(new_n704), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1002), .A2(new_n708), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n705), .A2(KEYINPUT62), .A3(new_n708), .A4(new_n1002), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n687), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n895), .A2(new_n896), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1013), .A2(new_n621), .A3(new_n888), .A4(new_n1014), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n814), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1012), .A2(new_n1016), .A3(new_n823), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n997), .B1(new_n1017), .B2(new_n427), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1006), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n427), .B1(G227), .B2(G900), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT124), .Z(new_n1021));
  XNOR2_X1  g835(.A(new_n1019), .B(new_n1021), .ZN(G72));
  NAND4_X1  g836(.A1(new_n1012), .A2(new_n1016), .A3(new_n823), .A4(new_n912), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT126), .ZN(new_n1024));
  XNOR2_X1  g838(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n630), .A2(new_n341), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1025), .B(new_n1026), .Z(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  AND3_X1   g842(.A1(new_n1023), .A2(new_n1024), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1024), .B1(new_n1023), .B2(new_n1028), .ZN(new_n1030));
  OAI211_X1 g844(.A(new_n557), .B(new_n603), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1005), .A2(new_n912), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT127), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1032), .A2(new_n1033), .A3(new_n1028), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n999), .A2(new_n1004), .A3(new_n902), .ZN(new_n1035));
  OAI21_X1  g849(.A(KEYINPUT127), .B1(new_n1035), .B2(new_n1027), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n603), .A2(new_n557), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n698), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1027), .B1(new_n1039), .B2(new_n604), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n938), .B1(new_n970), .B2(new_n1040), .ZN(new_n1041));
  AND3_X1   g855(.A1(new_n1031), .A2(new_n1038), .A3(new_n1041), .ZN(G57));
endmodule


