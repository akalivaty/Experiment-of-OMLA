

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XNOR2_X1 U326 ( .A(n348), .B(KEYINPUT33), .ZN(n349) );
  XNOR2_X1 U327 ( .A(n350), .B(n349), .ZN(n352) );
  XNOR2_X1 U328 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n416) );
  XNOR2_X1 U329 ( .A(n417), .B(n416), .ZN(n532) );
  XNOR2_X1 U330 ( .A(n357), .B(n392), .ZN(n358) );
  XNOR2_X1 U331 ( .A(n359), .B(n358), .ZN(n363) );
  NOR2_X1 U332 ( .A1(n535), .A2(n457), .ZN(n570) );
  XNOR2_X1 U333 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U334 ( .A(n465), .B(n464), .ZN(G1351GAT) );
  XOR2_X1 U335 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n300) );
  XOR2_X1 U336 ( .A(G169GAT), .B(KEYINPUT85), .Z(n295) );
  NAND2_X1 U337 ( .A1(G227GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n295), .B(n294), .ZN(n298) );
  XOR2_X1 U339 ( .A(G71GAT), .B(G120GAT), .Z(n297) );
  XNOR2_X1 U340 ( .A(G99GAT), .B(G176GAT), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n350) );
  XNOR2_X1 U342 ( .A(n298), .B(n350), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n300), .B(n299), .ZN(n302) );
  XNOR2_X1 U344 ( .A(G134GAT), .B(G127GAT), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n301), .B(KEYINPUT0), .ZN(n445) );
  XOR2_X1 U346 ( .A(n302), .B(n445), .Z(n310) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(G15GAT), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n303), .B(G113GAT), .ZN(n343) );
  XOR2_X1 U349 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n305) );
  XNOR2_X1 U350 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U352 ( .A(n306), .B(G183GAT), .Z(n308) );
  XNOR2_X1 U353 ( .A(KEYINPUT17), .B(G190GAT), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n433) );
  XNOR2_X1 U355 ( .A(n343), .B(n433), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n310), .B(n309), .ZN(n535) );
  XOR2_X1 U357 ( .A(KEYINPUT89), .B(KEYINPUT92), .Z(n312) );
  XNOR2_X1 U358 ( .A(G204GAT), .B(KEYINPUT90), .ZN(n311) );
  XNOR2_X1 U359 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U360 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n314) );
  NAND2_X1 U361 ( .A1(G228GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U363 ( .A(n316), .B(n315), .Z(n320) );
  XOR2_X1 U364 ( .A(KEYINPUT21), .B(G211GAT), .Z(n318) );
  XNOR2_X1 U365 ( .A(G197GAT), .B(G218GAT), .ZN(n317) );
  XNOR2_X1 U366 ( .A(n318), .B(n317), .ZN(n419) );
  XNOR2_X1 U367 ( .A(n419), .B(KEYINPUT23), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n323) );
  XOR2_X1 U369 ( .A(G78GAT), .B(KEYINPUT75), .Z(n322) );
  XNOR2_X1 U370 ( .A(G148GAT), .B(G106GAT), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n361) );
  XOR2_X1 U372 ( .A(n323), .B(n361), .Z(n329) );
  XNOR2_X1 U373 ( .A(G50GAT), .B(G22GAT), .ZN(n324) );
  XNOR2_X1 U374 ( .A(n324), .B(G141GAT), .ZN(n342) );
  XOR2_X1 U375 ( .A(G155GAT), .B(G162GAT), .Z(n326) );
  XNOR2_X1 U376 ( .A(KEYINPUT91), .B(KEYINPUT3), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U378 ( .A(KEYINPUT2), .B(n327), .Z(n438) );
  XNOR2_X1 U379 ( .A(n342), .B(n438), .ZN(n328) );
  XNOR2_X1 U380 ( .A(n329), .B(n328), .ZN(n477) );
  XOR2_X1 U381 ( .A(KEYINPUT47), .B(KEYINPUT111), .Z(n409) );
  XOR2_X1 U382 ( .A(KEYINPUT46), .B(KEYINPUT110), .Z(n330) );
  XNOR2_X1 U383 ( .A(KEYINPUT109), .B(n330), .ZN(n365) );
  XOR2_X1 U384 ( .A(KEYINPUT29), .B(KEYINPUT71), .Z(n332) );
  XNOR2_X1 U385 ( .A(KEYINPUT70), .B(KEYINPUT68), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n337) );
  XNOR2_X1 U387 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n333), .B(KEYINPUT7), .ZN(n367) );
  XOR2_X1 U389 ( .A(n367), .B(G1GAT), .Z(n335) );
  NAND2_X1 U390 ( .A1(G229GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n347) );
  XOR2_X1 U393 ( .A(KEYINPUT69), .B(G197GAT), .Z(n340) );
  XNOR2_X1 U394 ( .A(G169GAT), .B(G36GAT), .ZN(n338) );
  XOR2_X1 U395 ( .A(n338), .B(G8GAT), .Z(n418) );
  XOR2_X1 U396 ( .A(KEYINPUT30), .B(n418), .Z(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U398 ( .A(n341), .B(KEYINPUT72), .Z(n345) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n576) );
  INV_X1 U402 ( .A(n576), .ZN(n552) );
  AND2_X1 U403 ( .A1(G230GAT), .A2(G233GAT), .ZN(n348) );
  INV_X1 U404 ( .A(KEYINPUT32), .ZN(n351) );
  NAND2_X1 U405 ( .A1(n352), .A2(n351), .ZN(n355) );
  INV_X1 U406 ( .A(n352), .ZN(n353) );
  NAND2_X1 U407 ( .A1(n353), .A2(KEYINPUT32), .ZN(n354) );
  NAND2_X1 U408 ( .A1(n355), .A2(n354), .ZN(n359) );
  XOR2_X1 U409 ( .A(G85GAT), .B(KEYINPUT76), .Z(n366) );
  XOR2_X1 U410 ( .A(n366), .B(KEYINPUT31), .Z(n357) );
  XNOR2_X1 U411 ( .A(G57GAT), .B(KEYINPUT74), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n356), .B(KEYINPUT13), .ZN(n392) );
  XNOR2_X1 U413 ( .A(G92GAT), .B(G64GAT), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n360), .B(G204GAT), .ZN(n429) );
  XNOR2_X1 U415 ( .A(n361), .B(n429), .ZN(n362) );
  XNOR2_X1 U416 ( .A(n363), .B(n362), .ZN(n580) );
  XNOR2_X1 U417 ( .A(KEYINPUT41), .B(n580), .ZN(n555) );
  NAND2_X1 U418 ( .A1(n552), .A2(n555), .ZN(n364) );
  XNOR2_X1 U419 ( .A(n365), .B(n364), .ZN(n407) );
  XOR2_X1 U420 ( .A(n367), .B(n366), .Z(n369) );
  NAND2_X1 U421 ( .A1(G232GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n369), .B(n368), .ZN(n385) );
  XOR2_X1 U423 ( .A(KEYINPUT78), .B(KEYINPUT10), .Z(n371) );
  XNOR2_X1 U424 ( .A(KEYINPUT11), .B(KEYINPUT77), .ZN(n370) );
  XNOR2_X1 U425 ( .A(n371), .B(n370), .ZN(n383) );
  XOR2_X1 U426 ( .A(G92GAT), .B(G106GAT), .Z(n373) );
  XNOR2_X1 U427 ( .A(G99GAT), .B(G218GAT), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n381) );
  XOR2_X1 U429 ( .A(G162GAT), .B(G134GAT), .Z(n375) );
  XNOR2_X1 U430 ( .A(G43GAT), .B(G50GAT), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U432 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n377) );
  XNOR2_X1 U433 ( .A(G36GAT), .B(G190GAT), .ZN(n376) );
  XNOR2_X1 U434 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U435 ( .A(n379), .B(n378), .Z(n380) );
  XNOR2_X1 U436 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U437 ( .A(n383), .B(n382), .Z(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n466) );
  INV_X1 U439 ( .A(n466), .ZN(n562) );
  XOR2_X1 U440 ( .A(G78GAT), .B(G1GAT), .Z(n387) );
  XNOR2_X1 U441 ( .A(G15GAT), .B(G22GAT), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U443 ( .A(KEYINPUT81), .B(G155GAT), .Z(n389) );
  XNOR2_X1 U444 ( .A(G8GAT), .B(G183GAT), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U446 ( .A(n391), .B(n390), .Z(n397) );
  XOR2_X1 U447 ( .A(n392), .B(G64GAT), .Z(n394) );
  NAND2_X1 U448 ( .A1(G231GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U449 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U450 ( .A(G71GAT), .B(n395), .ZN(n396) );
  XNOR2_X1 U451 ( .A(n397), .B(n396), .ZN(n405) );
  XOR2_X1 U452 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n399) );
  XNOR2_X1 U453 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U455 ( .A(G211GAT), .B(KEYINPUT82), .Z(n401) );
  XNOR2_X1 U456 ( .A(G127GAT), .B(KEYINPUT15), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U458 ( .A(n403), .B(n402), .Z(n404) );
  XNOR2_X1 U459 ( .A(n405), .B(n404), .ZN(n571) );
  NOR2_X1 U460 ( .A1(n562), .A2(n571), .ZN(n406) );
  NAND2_X1 U461 ( .A1(n407), .A2(n406), .ZN(n408) );
  XNOR2_X1 U462 ( .A(n409), .B(n408), .ZN(n415) );
  XOR2_X1 U463 ( .A(KEYINPUT67), .B(KEYINPUT45), .Z(n411) );
  XNOR2_X1 U464 ( .A(KEYINPUT36), .B(n562), .ZN(n586) );
  NAND2_X1 U465 ( .A1(n586), .A2(n571), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n413) );
  XOR2_X1 U467 ( .A(n576), .B(KEYINPUT73), .Z(n458) );
  NAND2_X1 U468 ( .A1(n580), .A2(n458), .ZN(n412) );
  NOR2_X1 U469 ( .A1(n413), .A2(n412), .ZN(n414) );
  NOR2_X1 U470 ( .A1(n415), .A2(n414), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n419), .B(n418), .ZN(n427) );
  NAND2_X1 U472 ( .A1(G226GAT), .A2(G233GAT), .ZN(n425) );
  XOR2_X1 U473 ( .A(KEYINPUT97), .B(KEYINPUT99), .Z(n421) );
  XNOR2_X1 U474 ( .A(KEYINPUT79), .B(KEYINPUT98), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n423) );
  XOR2_X1 U476 ( .A(G176GAT), .B(KEYINPUT78), .Z(n422) );
  XNOR2_X1 U477 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U479 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U480 ( .A(n428), .B(KEYINPUT95), .Z(n431) );
  XNOR2_X1 U481 ( .A(n429), .B(KEYINPUT96), .ZN(n430) );
  XNOR2_X1 U482 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U483 ( .A(n433), .B(n432), .Z(n524) );
  NOR2_X1 U484 ( .A1(n532), .A2(n524), .ZN(n434) );
  XNOR2_X1 U485 ( .A(n434), .B(KEYINPUT54), .ZN(n453) );
  XOR2_X1 U486 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n436) );
  XNOR2_X1 U487 ( .A(KEYINPUT94), .B(KEYINPUT93), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n452) );
  XOR2_X1 U490 ( .A(G148GAT), .B(G57GAT), .Z(n440) );
  XNOR2_X1 U491 ( .A(G113GAT), .B(G120GAT), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U493 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n442) );
  XNOR2_X1 U494 ( .A(G141GAT), .B(G1GAT), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U496 ( .A(n444), .B(n443), .Z(n450) );
  XOR2_X1 U497 ( .A(G85GAT), .B(n445), .Z(n447) );
  NAND2_X1 U498 ( .A1(G225GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U500 ( .A(G29GAT), .B(n448), .ZN(n449) );
  XNOR2_X1 U501 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U502 ( .A(n452), .B(n451), .ZN(n522) );
  NAND2_X1 U503 ( .A1(n453), .A2(n522), .ZN(n454) );
  XNOR2_X1 U504 ( .A(n454), .B(KEYINPUT65), .ZN(n575) );
  NAND2_X1 U505 ( .A1(n477), .A2(n575), .ZN(n456) );
  INV_X1 U506 ( .A(KEYINPUT55), .ZN(n455) );
  XNOR2_X1 U507 ( .A(n456), .B(n455), .ZN(n457) );
  INV_X1 U508 ( .A(n458), .ZN(n536) );
  NAND2_X1 U509 ( .A1(n570), .A2(n536), .ZN(n461) );
  XOR2_X1 U510 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n459) );
  XNOR2_X1 U511 ( .A(n459), .B(G169GAT), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n461), .B(n460), .ZN(G1348GAT) );
  NAND2_X1 U513 ( .A1(n570), .A2(n562), .ZN(n465) );
  XOR2_X1 U514 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n463) );
  XNOR2_X1 U515 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n462) );
  NAND2_X1 U516 ( .A1(n571), .A2(n466), .ZN(n467) );
  XNOR2_X1 U517 ( .A(n467), .B(KEYINPUT83), .ZN(n468) );
  XNOR2_X1 U518 ( .A(n468), .B(KEYINPUT16), .ZN(n484) );
  XOR2_X1 U519 ( .A(n524), .B(KEYINPUT27), .Z(n475) );
  INV_X1 U520 ( .A(n475), .ZN(n469) );
  NOR2_X1 U521 ( .A1(n522), .A2(n469), .ZN(n530) );
  XOR2_X1 U522 ( .A(n477), .B(KEYINPUT28), .Z(n492) );
  INV_X1 U523 ( .A(n535), .ZN(n472) );
  XNOR2_X1 U524 ( .A(KEYINPUT88), .B(n472), .ZN(n470) );
  NOR2_X1 U525 ( .A1(n492), .A2(n470), .ZN(n471) );
  NAND2_X1 U526 ( .A1(n530), .A2(n471), .ZN(n483) );
  NOR2_X1 U527 ( .A1(n477), .A2(n472), .ZN(n474) );
  XNOR2_X1 U528 ( .A(KEYINPUT100), .B(KEYINPUT26), .ZN(n473) );
  XNOR2_X1 U529 ( .A(n474), .B(n473), .ZN(n574) );
  NAND2_X1 U530 ( .A1(n475), .A2(n574), .ZN(n480) );
  OR2_X1 U531 ( .A1(n535), .A2(n524), .ZN(n476) );
  NAND2_X1 U532 ( .A1(n477), .A2(n476), .ZN(n478) );
  XOR2_X1 U533 ( .A(KEYINPUT25), .B(n478), .Z(n479) );
  NAND2_X1 U534 ( .A1(n480), .A2(n479), .ZN(n481) );
  NAND2_X1 U535 ( .A1(n481), .A2(n522), .ZN(n482) );
  NAND2_X1 U536 ( .A1(n483), .A2(n482), .ZN(n495) );
  NAND2_X1 U537 ( .A1(n484), .A2(n495), .ZN(n511) );
  NAND2_X1 U538 ( .A1(n580), .A2(n536), .ZN(n500) );
  NOR2_X1 U539 ( .A1(n511), .A2(n500), .ZN(n485) );
  XNOR2_X1 U540 ( .A(n485), .B(KEYINPUT101), .ZN(n493) );
  NOR2_X1 U541 ( .A1(n522), .A2(n493), .ZN(n487) );
  XNOR2_X1 U542 ( .A(KEYINPUT102), .B(KEYINPUT34), .ZN(n486) );
  XNOR2_X1 U543 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U544 ( .A(G1GAT), .B(n488), .Z(G1324GAT) );
  NOR2_X1 U545 ( .A1(n524), .A2(n493), .ZN(n489) );
  XOR2_X1 U546 ( .A(G8GAT), .B(n489), .Z(G1325GAT) );
  NOR2_X1 U547 ( .A1(n535), .A2(n493), .ZN(n491) );
  XNOR2_X1 U548 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  INV_X1 U550 ( .A(n492), .ZN(n533) );
  NOR2_X1 U551 ( .A1(n533), .A2(n493), .ZN(n494) );
  XOR2_X1 U552 ( .A(G22GAT), .B(n494), .Z(G1327GAT) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n504) );
  INV_X1 U554 ( .A(n571), .ZN(n583) );
  NAND2_X1 U555 ( .A1(n583), .A2(n495), .ZN(n496) );
  XNOR2_X1 U556 ( .A(KEYINPUT103), .B(n496), .ZN(n497) );
  NAND2_X1 U557 ( .A1(n497), .A2(n586), .ZN(n499) );
  XOR2_X1 U558 ( .A(KEYINPUT37), .B(KEYINPUT104), .Z(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(n521) );
  NOR2_X1 U560 ( .A1(n521), .A2(n500), .ZN(n502) );
  XNOR2_X1 U561 ( .A(KEYINPUT38), .B(KEYINPUT105), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(n509) );
  NOR2_X1 U563 ( .A1(n522), .A2(n509), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  NOR2_X1 U565 ( .A1(n524), .A2(n509), .ZN(n505) );
  XOR2_X1 U566 ( .A(KEYINPUT106), .B(n505), .Z(n506) );
  XNOR2_X1 U567 ( .A(G36GAT), .B(n506), .ZN(G1329GAT) );
  NOR2_X1 U568 ( .A1(n535), .A2(n509), .ZN(n507) );
  XOR2_X1 U569 ( .A(KEYINPUT40), .B(n507), .Z(n508) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(n508), .ZN(G1330GAT) );
  NOR2_X1 U571 ( .A1(n509), .A2(n533), .ZN(n510) );
  XOR2_X1 U572 ( .A(G50GAT), .B(n510), .Z(G1331GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT107), .B(n555), .Z(n566) );
  NAND2_X1 U574 ( .A1(n576), .A2(n566), .ZN(n520) );
  OR2_X1 U575 ( .A1(n520), .A2(n511), .ZN(n516) );
  NOR2_X1 U576 ( .A1(n522), .A2(n516), .ZN(n512) );
  XOR2_X1 U577 ( .A(n512), .B(KEYINPUT42), .Z(n513) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(n513), .ZN(G1332GAT) );
  NOR2_X1 U579 ( .A1(n524), .A2(n516), .ZN(n514) );
  XOR2_X1 U580 ( .A(G64GAT), .B(n514), .Z(G1333GAT) );
  NOR2_X1 U581 ( .A1(n535), .A2(n516), .ZN(n515) );
  XOR2_X1 U582 ( .A(G71GAT), .B(n515), .Z(G1334GAT) );
  NOR2_X1 U583 ( .A1(n533), .A2(n516), .ZN(n518) );
  XNOR2_X1 U584 ( .A(KEYINPUT43), .B(KEYINPUT108), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(n519), .ZN(G1335GAT) );
  OR2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n527) );
  NOR2_X1 U588 ( .A1(n522), .A2(n527), .ZN(n523) );
  XOR2_X1 U589 ( .A(G85GAT), .B(n523), .Z(G1336GAT) );
  NOR2_X1 U590 ( .A1(n524), .A2(n527), .ZN(n525) );
  XOR2_X1 U591 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  NOR2_X1 U592 ( .A1(n535), .A2(n527), .ZN(n526) );
  XOR2_X1 U593 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  NOR2_X1 U594 ( .A1(n533), .A2(n527), .ZN(n528) );
  XOR2_X1 U595 ( .A(KEYINPUT44), .B(n528), .Z(n529) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n538) );
  INV_X1 U598 ( .A(n530), .ZN(n531) );
  NOR2_X1 U599 ( .A1(n532), .A2(n531), .ZN(n550) );
  NAND2_X1 U600 ( .A1(n550), .A2(n533), .ZN(n534) );
  NOR2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n546), .A2(n536), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n539), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n541) );
  NAND2_X1 U606 ( .A1(n546), .A2(n566), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n543) );
  XOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT114), .Z(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  NAND2_X1 U610 ( .A1(n571), .A2(n546), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n544), .B(KEYINPUT50), .ZN(n545) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U614 ( .A1(n546), .A2(n562), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G134GAT), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U617 ( .A1(n574), .A2(n550), .ZN(n551) );
  XNOR2_X1 U618 ( .A(KEYINPUT117), .B(n551), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n552), .A2(n563), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(KEYINPUT118), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n557) );
  NAND2_X1 U623 ( .A1(n563), .A2(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT53), .Z(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U627 ( .A1(n571), .A2(n563), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n560), .B(KEYINPUT120), .ZN(n561) );
  XNOR2_X1 U629 ( .A(G155GAT), .B(n561), .ZN(G1346GAT) );
  XOR2_X1 U630 ( .A(G162GAT), .B(KEYINPUT121), .Z(n565) );
  NAND2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1347GAT) );
  NAND2_X1 U633 ( .A1(n570), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(n569), .ZN(G1349GAT) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT124), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n585) );
  NOR2_X1 U641 ( .A1(n576), .A2(n585), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n585), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n585), .ZN(n584) );
  XOR2_X1 U649 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  INV_X1 U650 ( .A(n585), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

