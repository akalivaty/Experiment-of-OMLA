//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1215, new_n1216, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n210), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n213), .B1(new_n217), .B2(new_n218), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G50), .B(G68), .Z(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(KEYINPUT80), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT8), .B(G58), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT69), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G58), .ZN(new_n248));
  OR3_X1    g0048(.A1(new_n246), .A2(new_n248), .A3(KEYINPUT8), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT78), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n247), .A2(KEYINPUT78), .A3(new_n249), .A4(new_n253), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT68), .B1(new_n210), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n260), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n259), .A2(new_n214), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n262), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n256), .A2(new_n266), .B1(new_n267), .B2(new_n250), .ZN(new_n268));
  INV_X1    g0068(.A(G68), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT75), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n272), .A2(KEYINPUT75), .A3(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n215), .A3(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n271), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n279), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n276), .A2(new_n215), .A3(new_n277), .A4(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n269), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT16), .ZN(new_n284));
  AND2_X1   g0084(.A1(G58), .A2(G68), .ZN(new_n285));
  OAI21_X1  g0085(.A(G20), .B1(new_n285), .B2(new_n201), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT77), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G159), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n287), .B1(new_n286), .B2(new_n289), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n283), .A2(new_n284), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n259), .A2(new_n214), .A3(new_n261), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n286), .A2(new_n289), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT7), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT3), .B(G33), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(new_n297), .B2(G20), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n273), .A2(new_n274), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(KEYINPUT7), .A3(new_n215), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n295), .B1(new_n301), .B2(G68), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n294), .B1(new_n302), .B2(KEYINPUT16), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n268), .B1(new_n293), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G41), .A2(G45), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT67), .B1(new_n305), .B2(G1), .ZN(new_n306));
  AND2_X1   g0106(.A1(G1), .A2(G13), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G33), .A2(G41), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT67), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n310), .B(new_n252), .C1(G41), .C2(G45), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n306), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G232), .ZN(new_n313));
  INV_X1    g0113(.A(G274), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n307), .B2(new_n308), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n315), .B(new_n252), .C1(G41), .C2(G45), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n276), .A2(new_n277), .ZN(new_n318));
  INV_X1    g0118(.A(G1698), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(G223), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT79), .ZN(new_n321));
  AOI21_X1  g0121(.A(G1698), .B1(new_n276), .B2(new_n277), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT79), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(new_n323), .A3(G223), .ZN(new_n324));
  AND2_X1   g0124(.A1(G226), .A2(G1698), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n318), .A2(new_n325), .B1(G33), .B2(G87), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n321), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n317), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G179), .ZN(new_n332));
  AOI211_X1 g0132(.A(new_n332), .B(new_n317), .C1(new_n327), .C2(new_n328), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n304), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT18), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n329), .A2(G179), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n330), .B2(new_n329), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT18), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(new_n338), .A3(new_n304), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n244), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT78), .B1(new_n251), .B2(new_n253), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n341), .A2(new_n265), .B1(new_n262), .B2(new_n251), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n278), .A2(new_n279), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n343), .A2(new_n282), .A3(new_n270), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G68), .ZN(new_n345));
  INV_X1    g0145(.A(new_n292), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(KEYINPUT16), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n294), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n297), .A2(new_n296), .A3(G20), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT7), .B1(new_n299), .B2(new_n215), .ZN(new_n350));
  OAI21_X1  g0150(.A(G68), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n295), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n348), .B1(new_n353), .B2(new_n284), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n342), .B1(new_n347), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT82), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n327), .A2(new_n328), .ZN(new_n357));
  INV_X1    g0157(.A(new_n317), .ZN(new_n358));
  AOI21_X1  g0158(.A(G200), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AND2_X1   g0159(.A1(KEYINPUT81), .A2(G190), .ZN(new_n360));
  NOR2_X1   g0160(.A1(KEYINPUT81), .A2(G190), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AOI211_X1 g0163(.A(new_n363), .B(new_n317), .C1(new_n327), .C2(new_n328), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n355), .B(new_n356), .C1(new_n359), .C2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT17), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(KEYINPUT80), .A2(KEYINPUT18), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n334), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n357), .A2(new_n362), .A3(new_n358), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(G200), .B2(new_n329), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n371), .A2(new_n356), .A3(KEYINPUT17), .A4(new_n355), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n367), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n340), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n375));
  OR2_X1    g0175(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n288), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n215), .A2(G33), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n377), .B1(new_n250), .B2(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n379), .A2(new_n294), .B1(new_n202), .B2(new_n267), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n264), .A2(G50), .A3(new_n253), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT9), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n382), .B(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n312), .A2(G226), .ZN(new_n385));
  INV_X1    g0185(.A(G77), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n299), .A2(new_n386), .ZN(new_n387));
  MUX2_X1   g0187(.A(G222), .B(G223), .S(G1698), .Z(new_n388));
  OAI211_X1 g0188(.A(new_n387), .B(new_n328), .C1(new_n299), .C2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n385), .A2(new_n389), .A3(new_n316), .ZN(new_n390));
  INV_X1    g0190(.A(G190), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(G200), .B2(new_n390), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n375), .B(new_n376), .C1(new_n384), .C2(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n382), .B(KEYINPUT9), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n396), .A2(KEYINPUT71), .A3(KEYINPUT10), .A4(new_n393), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n390), .A2(new_n330), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n382), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT70), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n382), .A2(KEYINPUT70), .A3(new_n399), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n403), .C1(G179), .C2(new_n390), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n398), .A2(new_n405), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n288), .A2(G50), .B1(G20), .B2(new_n269), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n386), .B2(new_n378), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(KEYINPUT11), .A3(new_n294), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT11), .B1(new_n408), .B2(new_n294), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT73), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n411), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT73), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(new_n409), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n269), .B1(new_n252), .B2(G20), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT12), .B1(new_n262), .B2(G68), .ZN(new_n417));
  OR3_X1    g0217(.A1(new_n262), .A2(KEYINPUT12), .A3(G68), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n264), .A2(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n412), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n306), .A2(G238), .A3(new_n309), .A4(new_n311), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n258), .A2(new_n205), .ZN(new_n422));
  NOR2_X1   g0222(.A1(G226), .A2(G1698), .ZN(new_n423));
  INV_X1    g0223(.A(G232), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n423), .B1(new_n424), .B2(G1698), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n422), .B1(new_n425), .B2(new_n297), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n316), .B(new_n421), .C1(new_n426), .C2(new_n309), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT13), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n424), .A2(G1698), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G226), .B2(G1698), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n430), .A2(new_n299), .B1(new_n258), .B2(new_n205), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n328), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT13), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n316), .A4(new_n421), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n428), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT14), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(G169), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n332), .B2(new_n435), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n436), .B1(new_n435), .B2(G169), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n420), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n428), .A2(G190), .A3(new_n434), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT72), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n428), .A2(new_n434), .A3(KEYINPUT72), .A4(G190), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G200), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(new_n428), .B2(new_n434), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n420), .A2(new_n447), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n445), .A2(new_n448), .A3(KEYINPUT74), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT74), .B1(new_n445), .B2(new_n448), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n440), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G20), .A2(G77), .ZN(new_n453));
  XNOR2_X1  g0253(.A(KEYINPUT15), .B(G87), .ZN(new_n454));
  INV_X1    g0254(.A(new_n288), .ZN(new_n455));
  OAI221_X1 g0255(.A(new_n453), .B1(new_n454), .B2(new_n378), .C1(new_n455), .C2(new_n245), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(new_n294), .B1(new_n386), .B2(new_n267), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n264), .A2(G77), .A3(new_n253), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n316), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(new_n312), .B2(G244), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n297), .A2(G238), .A3(G1698), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n297), .A2(G232), .A3(new_n319), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n463), .C1(new_n206), .C2(new_n297), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n328), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n459), .B1(new_n466), .B2(G190), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n446), .B2(new_n466), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n461), .A2(new_n465), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n469), .A2(new_n330), .B1(new_n457), .B2(new_n458), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n466), .A2(new_n332), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n374), .A2(new_n406), .A3(new_n452), .A4(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT23), .B1(new_n206), .B2(G20), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G116), .ZN(new_n478));
  OAI22_X1  g0278(.A1(new_n476), .A2(new_n477), .B1(G20), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT22), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n297), .A2(new_n215), .A3(G87), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT24), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n318), .A2(KEYINPUT22), .A3(new_n215), .A4(G87), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n483), .B1(new_n482), .B2(new_n484), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n294), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n258), .A2(G1), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n263), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT83), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n261), .A2(new_n214), .ZN(new_n491));
  INV_X1    g0291(.A(new_n488), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n491), .A2(new_n259), .A3(new_n262), .A4(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT83), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n490), .A2(new_n495), .A3(G107), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n262), .A2(G107), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT25), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n487), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT87), .ZN(new_n500));
  INV_X1    g0300(.A(G257), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G1698), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(G250), .B2(G1698), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n277), .B2(new_n276), .ZN(new_n504));
  INV_X1    g0304(.A(G294), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n258), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(KEYINPUT86), .B(new_n328), .C1(new_n504), .C2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT5), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT84), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n508), .B1(new_n509), .B2(G41), .ZN(new_n510));
  INV_X1    g0310(.A(G45), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(G1), .ZN(new_n512));
  INV_X1    g0312(.A(G41), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n510), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(G264), .A3(new_n309), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n315), .A2(new_n510), .A3(new_n512), .A4(new_n514), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n507), .A2(new_n518), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n272), .A2(KEYINPUT75), .A3(G33), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n520), .B1(new_n297), .B2(new_n275), .ZN(new_n521));
  OAI22_X1  g0321(.A1(new_n521), .A2(new_n503), .B1(new_n258), .B2(new_n505), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT86), .B1(new_n522), .B2(new_n328), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n500), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n328), .B1(new_n504), .B2(new_n506), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT86), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n527), .A2(KEYINPUT87), .A3(new_n507), .A4(new_n518), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n330), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n525), .A2(new_n518), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(new_n332), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n499), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n499), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n524), .A2(new_n391), .A3(new_n528), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT88), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT88), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n524), .A2(new_n537), .A3(new_n528), .A4(new_n391), .ZN(new_n538));
  AOI21_X1  g0338(.A(G200), .B1(new_n525), .B2(new_n518), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n539), .B(KEYINPUT89), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n536), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n533), .B1(new_n534), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n515), .A2(G257), .A3(new_n309), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n297), .A2(G250), .A3(G1698), .ZN(new_n544));
  AND2_X1   g0344(.A1(KEYINPUT4), .A2(G244), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n273), .A2(new_n274), .A3(new_n545), .A4(new_n319), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G283), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n318), .A2(G244), .A3(new_n319), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT4), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n517), .B(new_n543), .C1(new_n551), .C2(new_n309), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n330), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT4), .B1(new_n322), .B2(G244), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n328), .B1(new_n554), .B2(new_n548), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n555), .A2(new_n332), .A3(new_n517), .A4(new_n543), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n490), .A2(new_n495), .A3(G97), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT6), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n558), .A2(new_n205), .A3(G107), .ZN(new_n559));
  XNOR2_X1  g0359(.A(G97), .B(G107), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n559), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n561), .A2(new_n215), .B1(new_n386), .B2(new_n455), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n206), .B1(new_n298), .B2(new_n300), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n294), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n267), .A2(new_n205), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n557), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n553), .A2(new_n556), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n552), .A2(G200), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n557), .A2(new_n564), .A3(new_n565), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n555), .A2(G190), .A3(new_n517), .A4(new_n543), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  OR2_X1    g0372(.A1(G238), .A2(G1698), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(G244), .B2(new_n319), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n277), .B2(new_n276), .ZN(new_n575));
  INV_X1    g0375(.A(new_n478), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n328), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(G250), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n328), .A2(new_n578), .A3(new_n512), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n512), .B2(new_n315), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G200), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n391), .B2(new_n581), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n490), .A2(new_n495), .A3(G87), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n521), .A2(G20), .A3(new_n269), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n378), .A2(KEYINPUT19), .A3(new_n205), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n422), .A2(G20), .B1(new_n207), .B2(G87), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(KEYINPUT19), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n294), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n454), .A2(new_n267), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n584), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n454), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n490), .A2(new_n495), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n589), .A3(new_n590), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n581), .A2(new_n330), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n577), .A2(new_n580), .A3(new_n332), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI22_X1  g0398(.A1(new_n583), .A2(new_n591), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT21), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n267), .A2(G116), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n493), .B2(G116), .ZN(new_n602));
  AOI21_X1  g0402(.A(G20), .B1(G33), .B2(G283), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n258), .A2(G97), .ZN(new_n604));
  INV_X1    g0404(.A(G116), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n603), .A2(new_n604), .B1(G20), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT20), .B1(new_n294), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT85), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n294), .A2(KEYINPUT20), .A3(new_n606), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n294), .A2(KEYINPUT85), .A3(new_n606), .A4(KEYINPUT20), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n602), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n501), .A2(new_n319), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(G264), .B2(new_n319), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n277), .B2(new_n276), .ZN(new_n615));
  INV_X1    g0415(.A(G303), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n297), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n328), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n515), .A2(G270), .A3(new_n309), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n619), .A2(new_n517), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G169), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n600), .B1(new_n612), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(G200), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n618), .A2(new_n620), .A3(new_n363), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n612), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n609), .A2(new_n608), .ZN(new_n627));
  INV_X1    g0427(.A(new_n607), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n628), .A3(new_n611), .ZN(new_n629));
  INV_X1    g0429(.A(new_n601), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n489), .B2(new_n605), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n618), .A2(new_n620), .A3(G179), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n330), .B1(new_n618), .B2(new_n620), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n632), .A2(KEYINPUT21), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n623), .A2(new_n626), .A3(new_n635), .A4(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n572), .A2(new_n599), .A3(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n475), .A2(new_n542), .A3(new_n639), .ZN(G372));
  NOR2_X1   g0440(.A1(new_n334), .A2(KEYINPUT18), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n338), .B1(new_n337), .B2(new_n304), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n472), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n449), .B2(new_n450), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n440), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n367), .A2(new_n372), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n644), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(KEYINPUT90), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(new_n398), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(KEYINPUT90), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n405), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n541), .A2(new_n534), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n623), .A2(new_n635), .A3(new_n637), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n532), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n572), .A2(new_n599), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n595), .A2(new_n598), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n596), .A2(new_n597), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n446), .B1(new_n577), .B2(new_n580), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n577), .A2(new_n580), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n661), .B1(G190), .B2(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n584), .A2(new_n589), .A3(new_n590), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n660), .A2(new_n594), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n569), .B1(new_n330), .B2(new_n552), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n665), .A2(KEYINPUT26), .A3(new_n666), .A4(new_n556), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n599), .B2(new_n567), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n659), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n658), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n475), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n653), .A2(new_n672), .ZN(G369));
  NAND3_X1  g0473(.A1(new_n252), .A2(new_n215), .A3(G13), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT91), .ZN(new_n676));
  INV_X1    g0476(.A(G213), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n674), .B2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n612), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT92), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n683), .B1(new_n638), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n684), .B2(new_n638), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n655), .A2(new_n683), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT93), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n542), .B1(new_n534), .B2(new_n682), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n532), .B2(new_n682), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n533), .A2(new_n682), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n655), .A2(new_n681), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n542), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n211), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n218), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT96), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n572), .B(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(new_n654), .A3(new_n665), .A4(new_n656), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n681), .B1(new_n708), .B2(new_n670), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n639), .A2(new_n654), .A3(new_n532), .A4(new_n682), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n555), .A2(new_n543), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n577), .A2(new_n525), .A3(new_n518), .A4(new_n580), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n713), .A2(new_n714), .A3(new_n633), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT94), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT30), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n714), .A2(new_n633), .ZN(new_n719));
  OAI211_X1 g0519(.A(KEYINPUT94), .B(new_n718), .C1(new_n719), .C2(new_n713), .ZN(new_n720));
  AOI21_X1  g0520(.A(G179), .B1(new_n577), .B2(new_n580), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n721), .A2(KEYINPUT95), .A3(new_n621), .ZN(new_n722));
  AOI21_X1  g0522(.A(KEYINPUT95), .B1(new_n721), .B2(new_n621), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n530), .B(new_n552), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n717), .A2(new_n720), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n681), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n712), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n730), .A2(G330), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n681), .B1(new_n658), .B2(new_n670), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(KEYINPUT29), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n711), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n705), .B1(new_n735), .B2(G1), .ZN(G364));
  AND2_X1   g0536(.A1(new_n215), .A2(G13), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n252), .B1(new_n737), .B2(G45), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n700), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n689), .A2(G330), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT97), .Z(new_n742));
  AOI211_X1 g0542(.A(new_n740), .B(new_n742), .C1(G330), .C2(new_n689), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n740), .B(KEYINPUT98), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n699), .A2(new_n299), .ZN(new_n746));
  AOI22_X1  g0546(.A1(G355), .A2(new_n746), .B1(new_n605), .B2(new_n699), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n242), .A2(new_n511), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n318), .A2(new_n699), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(G45), .B2(new_n218), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n747), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  OR3_X1    g0551(.A1(KEYINPUT99), .A2(G13), .A3(G33), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT99), .B1(G13), .B2(G33), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n214), .B1(G20), .B2(new_n330), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n745), .B1(new_n751), .B2(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n215), .A2(new_n332), .A3(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n391), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n299), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n363), .A2(new_n760), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n215), .A2(G179), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(G190), .A3(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n765), .A2(G322), .B1(G303), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G283), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n766), .A2(new_n391), .A3(G200), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n215), .A2(new_n332), .A3(new_n446), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT33), .B(G317), .Z(new_n776));
  OAI221_X1 g0576(.A(new_n769), .B1(new_n770), .B2(new_n771), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G179), .A2(G200), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT100), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n779), .A2(new_n215), .A3(G190), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n763), .B(new_n777), .C1(G329), .C2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(G20), .B1(new_n779), .B2(new_n391), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n773), .A2(new_n362), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n782), .A2(G294), .B1(new_n783), .B2(G326), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT102), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(KEYINPUT102), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n781), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n780), .A2(G159), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT32), .ZN(new_n789));
  INV_X1    g0589(.A(new_n761), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n299), .B1(new_n790), .B2(G77), .ZN(new_n791));
  INV_X1    g0591(.A(G87), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n791), .B1(new_n248), .B2(new_n764), .C1(new_n792), .C2(new_n767), .ZN(new_n793));
  INV_X1    g0593(.A(new_n782), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n205), .ZN(new_n795));
  INV_X1    g0595(.A(new_n771), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n774), .A2(G68), .B1(G107), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n783), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n202), .B2(new_n798), .ZN(new_n799));
  NOR4_X1   g0599(.A1(new_n789), .A2(new_n793), .A3(new_n795), .A4(new_n799), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n800), .A2(KEYINPUT101), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n787), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(KEYINPUT101), .B2(new_n800), .ZN(new_n803));
  INV_X1    g0603(.A(new_n757), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n759), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(new_n688), .B2(new_n756), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT103), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n743), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  NAND2_X1  g0609(.A1(new_n459), .A2(new_n681), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n468), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n472), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n472), .A2(new_n681), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n733), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n815), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n732), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n730), .A2(G330), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n740), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n820), .B2(new_n819), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n754), .A2(new_n757), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n745), .B1(new_n386), .B2(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT104), .Z(new_n825));
  AOI21_X1  g0625(.A(new_n297), .B1(new_n765), .B2(G294), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n771), .A2(new_n792), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G107), .B2(new_n768), .ZN(new_n828));
  INV_X1    g0628(.A(new_n780), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n826), .B(new_n828), .C1(new_n762), .C2(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n774), .A2(G283), .B1(new_n790), .B2(G116), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n616), .B2(new_n798), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n830), .A2(new_n795), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n521), .B1(G68), .B2(new_n796), .ZN(new_n834));
  INV_X1    g0634(.A(G132), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n202), .B2(new_n767), .C1(new_n829), .C2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G58), .B2(new_n782), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT105), .Z(new_n838));
  AOI22_X1  g0638(.A1(new_n783), .A2(G137), .B1(new_n790), .B2(G159), .ZN(new_n839));
  INV_X1    g0639(.A(G143), .ZN(new_n840));
  INV_X1    g0640(.A(G150), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n839), .B1(new_n840), .B2(new_n764), .C1(new_n841), .C2(new_n775), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT34), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n833), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n825), .B1(new_n844), .B2(new_n804), .C1(new_n817), .C2(new_n755), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n822), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G384));
  INV_X1    g0647(.A(new_n561), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n605), .B(new_n217), .C1(new_n848), .C2(KEYINPUT35), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(KEYINPUT35), .B2(new_n848), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT36), .Z(new_n851));
  NOR3_X1   g0651(.A1(new_n218), .A2(new_n285), .A3(new_n386), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT106), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n852), .A2(new_n853), .B1(new_n202), .B2(G68), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n252), .B(G13), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT40), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT107), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n292), .B1(new_n344), .B2(G68), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n348), .B1(new_n860), .B2(KEYINPUT16), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n284), .B1(new_n283), .B2(new_n292), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n342), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n859), .B1(new_n863), .B2(new_n679), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n347), .A2(new_n862), .A3(new_n294), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n268), .ZN(new_n866));
  INV_X1    g0666(.A(new_n679), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n866), .A2(KEYINPUT107), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n355), .B1(new_n359), .B2(new_n364), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n331), .A2(new_n333), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n870), .B1(new_n871), .B2(new_n863), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT37), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n304), .A2(new_n867), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n334), .A2(new_n870), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n869), .B1(new_n340), .B2(new_n373), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n877), .A2(new_n878), .A3(KEYINPUT38), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT38), .B1(new_n877), .B2(new_n878), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n420), .A2(new_n681), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n451), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n440), .B(new_n882), .C1(new_n449), .C2(new_n450), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n815), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n730), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n858), .B1(new_n881), .B2(new_n887), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n730), .A2(new_n886), .A3(KEYINPUT40), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n334), .A2(new_n870), .A3(new_n875), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n876), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n367), .A2(new_n335), .A3(new_n339), .A4(new_n372), .ZN(new_n893));
  INV_X1    g0693(.A(new_n875), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n892), .A2(KEYINPUT109), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT109), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n891), .A2(new_n896), .A3(new_n876), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n889), .B1(new_n898), .B2(new_n879), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n888), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n475), .A2(new_n730), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(G330), .A3(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT111), .Z(new_n905));
  NOR3_X1   g0705(.A1(new_n898), .A2(new_n879), .A3(KEYINPUT39), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  INV_X1    g0708(.A(new_n869), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n367), .A2(new_n369), .A3(new_n372), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT80), .B1(new_n641), .B2(new_n642), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n876), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n337), .A2(new_n866), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n864), .A2(new_n868), .A3(new_n914), .A4(new_n870), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n913), .B1(KEYINPUT37), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n908), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n877), .A2(new_n878), .A3(KEYINPUT38), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n907), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT110), .B1(new_n906), .B2(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n440), .A2(new_n681), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT108), .Z(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n892), .A2(KEYINPUT109), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n893), .A2(new_n894), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n924), .A2(new_n897), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n908), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n907), .A3(new_n918), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT39), .B1(new_n879), .B2(new_n880), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT110), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n920), .A2(new_n923), .A3(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n881), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n884), .A2(new_n885), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n818), .B2(new_n814), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n933), .A2(new_n935), .B1(new_n644), .B2(new_n679), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n475), .B1(new_n711), .B2(new_n734), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n653), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n937), .B(new_n939), .Z(new_n940));
  OAI22_X1  g0740(.A1(new_n905), .A2(new_n940), .B1(new_n252), .B2(new_n737), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n905), .A2(new_n940), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n857), .B1(new_n941), .B2(new_n942), .ZN(G367));
  NAND2_X1  g0743(.A1(new_n235), .A2(new_n749), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n757), .B(new_n756), .C1(new_n699), .C2(new_n592), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n745), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n756), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n591), .A2(new_n681), .ZN(new_n948));
  MUX2_X1   g0748(.A(new_n659), .B(new_n665), .S(new_n948), .Z(new_n949));
  AOI22_X1  g0749(.A1(new_n765), .A2(G303), .B1(new_n783), .B2(G311), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n951), .A2(KEYINPUT114), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(KEYINPUT114), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n521), .B1(new_n205), .B2(new_n771), .C1(new_n775), .C2(new_n505), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n767), .A2(new_n605), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(KEYINPUT46), .ZN(new_n957));
  XOR2_X1   g0757(.A(KEYINPUT115), .B(G317), .Z(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n780), .A2(new_n959), .B1(new_n956), .B2(KEYINPUT46), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n782), .A2(G107), .B1(G283), .B2(new_n790), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT113), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n955), .A2(new_n957), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n782), .A2(G68), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n841), .B2(new_n764), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT116), .Z(new_n966));
  INV_X1    g0766(.A(G137), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n297), .B1(new_n202), .B2(new_n761), .C1(new_n829), .C2(new_n967), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n774), .A2(G159), .B1(G58), .B2(new_n768), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n969), .B1(new_n386), .B2(new_n771), .C1(new_n840), .C2(new_n798), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n963), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT47), .Z(new_n973));
  OAI221_X1 g0773(.A(new_n946), .B1(new_n947), .B2(new_n949), .C1(new_n973), .C2(new_n804), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n566), .A2(new_n681), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n707), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n666), .A2(new_n556), .A3(new_n681), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(new_n695), .A3(new_n697), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT45), .Z(new_n980));
  AOI21_X1  g0780(.A(new_n978), .B1(new_n695), .B2(new_n697), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT44), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n694), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n980), .A2(new_n982), .A3(new_n694), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n697), .B1(new_n693), .B2(new_n696), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n690), .B(new_n987), .Z(new_n988));
  NAND4_X1  g0788(.A1(new_n985), .A2(new_n735), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT112), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AND3_X1   g0791(.A1(new_n980), .A2(new_n982), .A3(new_n694), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n694), .B1(new_n980), .B2(new_n982), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n988), .A2(new_n735), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT112), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n735), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n700), .B(KEYINPUT41), .Z(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n739), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n978), .A2(new_n542), .A3(new_n696), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(KEYINPUT42), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n707), .A2(new_n533), .A3(new_n975), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n681), .B1(new_n1003), .B2(new_n567), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n1001), .B2(KEYINPUT42), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n1002), .A2(new_n1005), .B1(KEYINPUT43), .B2(new_n949), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n984), .A2(new_n978), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1008), .B(new_n1009), .Z(new_n1010));
  OAI21_X1  g0810(.A(new_n974), .B1(new_n1000), .B2(new_n1010), .ZN(G387));
  NOR2_X1   g0811(.A1(new_n995), .A2(new_n701), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n735), .B2(new_n988), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n988), .A2(new_n739), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n702), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n746), .A2(new_n1015), .B1(new_n206), .B2(new_n699), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n232), .A2(new_n511), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n245), .A2(G50), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT50), .Z(new_n1019));
  OAI211_X1 g0819(.A(new_n702), .B(new_n511), .C1(new_n269), .C2(new_n386), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n749), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1016), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n745), .B1(new_n1022), .B2(new_n758), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n521), .B1(G97), .B2(new_n796), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n775), .B2(new_n250), .C1(new_n829), .C2(new_n841), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n783), .A2(G159), .B1(new_n790), .B2(G68), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n202), .B2(new_n764), .C1(new_n386), .C2(new_n767), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1025), .B(new_n1027), .C1(new_n592), .C2(new_n782), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G322), .A2(new_n783), .B1(new_n774), .B2(G311), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n616), .B2(new_n761), .C1(new_n764), .C2(new_n958), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT48), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n782), .A2(G283), .B1(G294), .B2(new_n768), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT49), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n521), .B1(new_n605), .B2(new_n771), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G326), .B2(new_n780), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT117), .Z(new_n1040));
  NOR2_X1   g0840(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1028), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1023), .B1(new_n804), .B2(new_n1043), .C1(new_n693), .C2(new_n947), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1013), .A2(new_n1014), .A3(new_n1044), .ZN(G393));
  OAI221_X1 g0845(.A(new_n700), .B1(new_n994), .B2(new_n995), .C1(new_n991), .C2(new_n996), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n749), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n758), .B1(new_n205), .B2(new_n211), .C1(new_n239), .C2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n744), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n775), .A2(new_n616), .B1(new_n761), .B2(new_n505), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n297), .B(new_n1050), .C1(G107), .C2(new_n796), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n765), .A2(G311), .B1(new_n783), .B2(G317), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT52), .Z(new_n1053));
  OAI211_X1 g0853(.A(new_n1051), .B(new_n1053), .C1(new_n605), .C2(new_n794), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n780), .A2(G322), .B1(G283), .B2(new_n768), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT118), .Z(new_n1056));
  AOI211_X1 g0856(.A(new_n521), .B(new_n827), .C1(new_n780), .C2(G143), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n774), .A2(G50), .B1(G68), .B2(new_n768), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n245), .C2(new_n761), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n765), .A2(G159), .B1(new_n783), .B2(G150), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1060), .A2(KEYINPUT51), .B1(G77), .B2(new_n782), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(KEYINPUT51), .B2(new_n1060), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n1054), .A2(new_n1056), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1049), .B1(new_n1063), .B2(new_n757), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n978), .B2(new_n947), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n994), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(new_n1066), .B2(new_n738), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1046), .A2(new_n1068), .ZN(G390));
  OR3_X1    g0869(.A1(new_n820), .A2(new_n815), .A3(new_n934), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT119), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n935), .B2(new_n923), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n813), .B1(new_n732), .B2(new_n817), .ZN(new_n1074));
  OAI211_X1 g0874(.A(KEYINPUT119), .B(new_n922), .C1(new_n1074), .C2(new_n934), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n920), .B2(new_n931), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n813), .B1(new_n709), .B2(new_n812), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1078), .A2(new_n934), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n927), .A2(new_n918), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n1080), .A3(new_n922), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1071), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n928), .A2(new_n930), .A3(new_n929), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n930), .B1(new_n928), .B2(new_n929), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1070), .B(new_n1081), .C1(new_n1086), .C2(new_n1076), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n731), .A2(new_n475), .A3(KEYINPUT120), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT120), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n820), .B2(new_n474), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n653), .A2(new_n1092), .A3(new_n938), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1074), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n884), .A2(new_n885), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n731), .B2(new_n817), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1094), .B1(new_n1071), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n731), .A2(KEYINPUT121), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT121), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n817), .B1(new_n820), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n934), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n1070), .A3(new_n1078), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1093), .B1(new_n1097), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1088), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1083), .A2(new_n1087), .A3(new_n1103), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n700), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1083), .A2(new_n1087), .A3(new_n739), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT54), .B(G143), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n775), .A2(new_n967), .B1(new_n761), .B2(new_n1109), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n764), .A2(new_n835), .B1(new_n202), .B2(new_n771), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n780), .A2(G125), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n299), .B(new_n1113), .C1(G128), .C2(new_n783), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n782), .A2(G159), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n767), .A2(new_n841), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT53), .ZN(new_n1117));
  AND4_X1   g0917(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G77), .A2(new_n782), .B1(new_n765), .B2(G116), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT122), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n790), .A2(G97), .B1(new_n796), .B2(G68), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1121), .B1(new_n798), .B2(new_n770), .C1(new_n206), .C2(new_n775), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n299), .B1(new_n792), .B2(new_n767), .C1(new_n829), .C2(new_n505), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1120), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n757), .B1(new_n1118), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n745), .B1(new_n250), .B2(new_n823), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1125), .B(new_n1126), .C1(new_n1086), .C2(new_n755), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1108), .A2(KEYINPUT123), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT123), .B1(new_n1108), .B2(new_n1127), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1107), .B1(new_n1128), .B2(new_n1129), .ZN(G378));
  NAND2_X1  g0930(.A1(new_n382), .A2(new_n867), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n406), .B(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1132), .B(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n888), .A2(new_n1135), .A3(G330), .A4(new_n899), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n887), .B1(new_n917), .B2(new_n918), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n899), .B(G330), .C1(KEYINPUT40), .C2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1132), .B(new_n1133), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AND4_X1   g0940(.A1(new_n932), .A2(new_n936), .A3(new_n1136), .A4(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n932), .A2(new_n936), .B1(new_n1140), .B2(new_n1136), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT125), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1140), .A2(new_n1136), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n937), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n932), .A2(new_n936), .A3(new_n1140), .A4(new_n1136), .ZN(new_n1147));
  AOI21_X1  g0947(.A(KEYINPUT125), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1093), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1106), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT57), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT57), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n700), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n823), .A2(new_n202), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n774), .A2(G97), .B1(G77), .B2(new_n768), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(new_n513), .A3(new_n521), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n765), .A2(G107), .B1(new_n783), .B2(G116), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n790), .A2(new_n592), .B1(new_n796), .B2(G58), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n964), .A3(new_n1162), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1160), .B(new_n1163), .C1(G283), .C2(new_n780), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT124), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1165), .A2(KEYINPUT58), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(KEYINPUT58), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G125), .A2(new_n783), .B1(new_n774), .B2(G132), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n782), .A2(G150), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1109), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n790), .A2(G137), .B1(new_n768), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n765), .A2(G128), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n780), .A2(G124), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G33), .B(G41), .C1(new_n796), .C2(G159), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1167), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n513), .B1(new_n521), .B2(new_n258), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1166), .B(new_n1179), .C1(new_n202), .C2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n740), .B(new_n1158), .C1(new_n1181), .C2(new_n804), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1139), .B2(new_n754), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1149), .B2(new_n739), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1157), .A2(new_n1184), .ZN(G375));
  NAND2_X1  g0985(.A1(new_n1102), .A2(new_n1097), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n934), .A2(new_n754), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n782), .A2(G50), .B1(G150), .B2(new_n790), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT126), .Z(new_n1189));
  AOI22_X1  g0989(.A1(new_n765), .A2(G137), .B1(G159), .B2(new_n768), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G132), .A2(new_n783), .B1(new_n774), .B2(new_n1170), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n318), .B1(new_n248), .B2(new_n771), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n780), .B2(G128), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n1193), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n764), .A2(new_n770), .B1(new_n205), .B2(new_n767), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n297), .B(new_n1195), .C1(G77), .C2(new_n796), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n775), .A2(new_n605), .B1(new_n761), .B2(new_n206), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G294), .B2(new_n783), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n782), .A2(new_n592), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n780), .A2(G303), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1196), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n804), .B1(new_n1194), .B2(new_n1201), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n745), .B(new_n1202), .C1(new_n269), .C2(new_n823), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1186), .A2(new_n739), .B1(new_n1187), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1104), .A2(new_n999), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1186), .A2(new_n1150), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(G381));
  INV_X1    g1007(.A(G375), .ZN(new_n1208));
  INV_X1    g1008(.A(G387), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1108), .A2(new_n1127), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1107), .A2(new_n1210), .ZN(new_n1211));
  OR2_X1    g1011(.A1(G393), .A2(G396), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(new_n1212), .A2(G390), .A3(G384), .A4(G381), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1208), .A2(new_n1209), .A3(new_n1211), .A4(new_n1213), .ZN(G407));
  NOR2_X1   g1014(.A1(new_n677), .A2(G343), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1208), .A2(new_n1211), .A3(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(G407), .A2(G213), .A3(new_n1216), .ZN(G409));
  NAND3_X1  g1017(.A1(G387), .A2(new_n1046), .A3(new_n1068), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(G393), .B(new_n808), .ZN(new_n1219));
  OAI211_X1 g1019(.A(G390), .B(new_n974), .C1(new_n1000), .C2(new_n1010), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1219), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(G378), .B(new_n1184), .C1(new_n1152), .C2(new_n1156), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1143), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1146), .A2(KEYINPUT125), .A3(new_n1147), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1151), .A2(new_n1226), .A3(new_n999), .A4(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1183), .B1(new_n1225), .B2(new_n739), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1211), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1215), .B1(new_n1224), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1206), .B1(new_n1104), .B2(KEYINPUT60), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1093), .A2(new_n1102), .A3(new_n1097), .A4(KEYINPUT60), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n700), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1204), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n846), .ZN(new_n1238));
  OAI211_X1 g1038(.A(G384), .B(new_n1204), .C1(new_n1234), .C2(new_n1236), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1215), .A2(G2897), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1240), .B(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT61), .B1(new_n1233), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1240), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1232), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT63), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1215), .B(new_n1240), .C1(new_n1224), .C2(new_n1231), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(KEYINPUT63), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1223), .A2(new_n1243), .A3(new_n1247), .A4(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT61), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1242), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n1232), .ZN(new_n1253));
  AND2_X1   g1053(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1254), .B1(new_n1248), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1245), .A2(new_n1255), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1253), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1250), .B1(new_n1259), .B2(new_n1223), .ZN(G405));
  NAND2_X1  g1060(.A1(G375), .A2(new_n1211), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n1224), .A3(new_n1240), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1240), .B1(new_n1261), .B2(new_n1224), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n1263), .A2(new_n1264), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1264), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(new_n1223), .A3(new_n1262), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(G402));
endmodule


