//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n552,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n586, new_n587, new_n588,
    new_n591, new_n593, new_n594, new_n595, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT68), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n463), .A2(new_n466), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(new_n468), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n462), .A2(G2105), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NOR3_X1   g052(.A1(new_n471), .A2(new_n475), .A3(new_n477), .ZN(G160));
  INV_X1    g053(.A(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n467), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  OAI22_X1  g056(.A1(new_n469), .A2(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR3_X1   g057(.A1(new_n462), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n465), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n485), .A2(KEYINPUT69), .A3(G2105), .A4(new_n463), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n463), .A2(new_n466), .A3(G2105), .A4(new_n468), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n482), .B1(new_n490), .B2(G124), .ZN(G162));
  NAND2_X1  g066(.A1(KEYINPUT4), .A2(G138), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n469), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n472), .A2(new_n468), .A3(G138), .A4(new_n467), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT71), .A2(G114), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT71), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n494), .A2(new_n495), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n463), .A2(new_n466), .A3(new_n468), .A4(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n503), .A2(new_n504), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n493), .B(new_n501), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  OR2_X1    g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(new_n517), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n511), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n514), .A2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND3_X1  g100(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n526));
  XOR2_X1   g101(.A(new_n526), .B(KEYINPUT72), .Z(new_n527));
  AOI21_X1  g102(.A(new_n527), .B1(G51), .B2(new_n518), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n509), .A2(new_n510), .B1(new_n516), .B2(new_n517), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n529), .A2(G89), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(KEYINPUT74), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  OR3_X1    g109(.A1(new_n530), .A2(new_n533), .A3(KEYINPUT74), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n528), .A2(new_n534), .A3(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  AOI22_X1  g112(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n513), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n518), .A2(G52), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n521), .B2(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n539), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  AOI22_X1  g119(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n513), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n518), .A2(G43), .ZN(new_n547));
  XNOR2_X1  g122(.A(KEYINPUT75), .B(G81), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n521), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(G188));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n518), .A2(new_n557), .A3(G53), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n529), .A2(G91), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n559), .B(new_n560), .C1(new_n513), .C2(new_n561), .ZN(G299));
  NAND2_X1  g137(.A1(new_n529), .A2(G87), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n518), .A2(G49), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(G288));
  AND2_X1   g141(.A1(new_n511), .A2(G61), .ZN(new_n567));
  NAND2_X1  g142(.A1(G73), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n529), .A2(G86), .B1(new_n518), .B2(G48), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(G305));
  AOI22_X1  g147(.A1(new_n529), .A2(G85), .B1(new_n518), .B2(G47), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n513), .B2(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(G301), .A2(G868), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n529), .A2(G92), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT10), .Z(new_n578));
  NAND2_X1  g153(.A1(new_n511), .A2(G66), .ZN(new_n579));
  INV_X1    g154(.A(G79), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n580), .B2(new_n515), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(G54), .B2(new_n518), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n576), .B1(new_n583), .B2(G868), .ZN(G284));
  XNOR2_X1  g159(.A(G284), .B(KEYINPUT77), .ZN(G321));
  INV_X1    g160(.A(G868), .ZN(new_n586));
  NOR2_X1   g161(.A1(G286), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g162(.A(G299), .B(KEYINPUT78), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n587), .B1(new_n586), .B2(new_n588), .ZN(G297));
  AOI21_X1  g164(.A(new_n587), .B1(new_n586), .B2(new_n588), .ZN(G280));
  INV_X1    g165(.A(G559), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n583), .B1(new_n591), .B2(G860), .ZN(G148));
  INV_X1    g167(.A(new_n550), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n583), .A2(new_n591), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT79), .ZN(new_n595));
  MUX2_X1   g170(.A(new_n593), .B(new_n595), .S(G868), .Z(G323));
  XNOR2_X1  g171(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g172(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n598));
  INV_X1    g173(.A(G111), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G2105), .ZN(new_n600));
  AND4_X1   g175(.A1(new_n467), .A2(new_n463), .A3(new_n466), .A4(new_n468), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G135), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n490), .B2(G123), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(G2096), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(G2096), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT80), .B(G2100), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT12), .Z(new_n611));
  XNOR2_X1  g186(.A(new_n609), .B(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n606), .A2(new_n607), .A3(new_n612), .ZN(G156));
  XOR2_X1   g188(.A(G2451), .B(G2454), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT16), .ZN(new_n615));
  XNOR2_X1  g190(.A(G1341), .B(G1348), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT81), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n615), .B(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT14), .ZN(new_n619));
  XNOR2_X1  g194(.A(G2427), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT15), .B(G2435), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n622), .B2(new_n621), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n618), .B(new_n624), .Z(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(G14), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(new_n628), .B2(new_n626), .ZN(G401));
  XNOR2_X1  g205(.A(G2072), .B(G2078), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT17), .Z(new_n634));
  XNOR2_X1  g209(.A(G2067), .B(G2678), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2084), .B(G2090), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n633), .B2(new_n635), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT83), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n636), .A2(new_n638), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n633), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT18), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n635), .A2(new_n638), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n644), .B1(new_n634), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(G2100), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT84), .B(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n647), .B(G2100), .ZN(new_n652));
  INV_X1    g227(.A(new_n650), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n651), .A2(new_n654), .ZN(G227));
  XOR2_X1   g230(.A(G1971), .B(G1976), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1956), .B(G2474), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1961), .B(G1966), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n657), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n657), .A2(new_n660), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT20), .Z(new_n664));
  AOI211_X1 g239(.A(new_n662), .B(new_n664), .C1(new_n657), .C2(new_n661), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1991), .B(G1996), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G229));
  XOR2_X1   g246(.A(KEYINPUT31), .B(G11), .Z(new_n672));
  INV_X1    g247(.A(G16), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n550), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n673), .B2(G19), .ZN(new_n675));
  INV_X1    g250(.A(G1341), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G29), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT30), .B(G28), .ZN(new_n679));
  AOI211_X1 g254(.A(new_n672), .B(new_n677), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n673), .A2(G5), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(G171), .B2(new_n673), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n682), .A2(G1961), .ZN(new_n683));
  AOI22_X1  g258(.A1(new_n676), .A2(new_n675), .B1(new_n682), .B2(G1961), .ZN(new_n684));
  INV_X1    g259(.A(G34), .ZN(new_n685));
  AOI21_X1  g260(.A(G29), .B1(new_n685), .B2(KEYINPUT24), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(KEYINPUT24), .B2(new_n685), .ZN(new_n687));
  INV_X1    g262(.A(G160), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n678), .ZN(new_n689));
  INV_X1    g264(.A(G2084), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g266(.A1(new_n680), .A2(new_n683), .A3(new_n684), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n673), .A2(G20), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT23), .Z(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G299), .B2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT93), .B(G1956), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G2078), .ZN(new_n698));
  NOR2_X1   g273(.A1(G164), .A2(new_n678), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G27), .B2(new_n678), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n697), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n692), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n583), .A2(new_n673), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G4), .B2(new_n673), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n705), .A2(G1348), .B1(G29), .B2(new_n604), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n702), .B(new_n706), .C1(G1348), .C2(new_n705), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n673), .A2(G21), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G168), .B2(new_n673), .ZN(new_n709));
  INV_X1    g284(.A(G1966), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n678), .A2(G26), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  INV_X1    g288(.A(G128), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n486), .B2(new_n489), .ZN(new_n715));
  INV_X1    g290(.A(G140), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n467), .A2(G116), .ZN(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n718));
  OAI22_X1  g293(.A1(new_n469), .A2(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n713), .B1(new_n720), .B2(new_n678), .ZN(new_n721));
  INV_X1    g296(.A(G2067), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n700), .A2(new_n698), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n711), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n476), .A2(G105), .ZN(new_n726));
  INV_X1    g301(.A(G141), .ZN(new_n727));
  AND3_X1   g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT26), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(KEYINPUT89), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT89), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(KEYINPUT26), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n728), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n728), .A2(new_n730), .A3(new_n732), .ZN(new_n734));
  OAI221_X1 g309(.A(new_n726), .B1(new_n469), .B2(new_n727), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G129), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n486), .B2(new_n489), .ZN(new_n737));
  NOR3_X1   g312(.A1(new_n735), .A2(new_n737), .A3(KEYINPUT90), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT90), .ZN(new_n739));
  INV_X1    g314(.A(new_n489), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n487), .A2(new_n488), .ZN(new_n741));
  OAI21_X1  g316(.A(G129), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n726), .B1(new_n734), .B2(new_n733), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n469), .A2(new_n727), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n739), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n738), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G29), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G29), .B2(G32), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT27), .B(G1996), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G2090), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n678), .A2(G35), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G162), .B2(new_n678), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT29), .Z(new_n755));
  AOI21_X1  g330(.A(new_n751), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n752), .B2(new_n755), .ZN(new_n757));
  NOR3_X1   g332(.A1(new_n707), .A2(new_n725), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n678), .A2(G33), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n601), .A2(G139), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT25), .Z(new_n762));
  AND2_X1   g337(.A1(new_n472), .A2(new_n468), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n763), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n760), .B(new_n762), .C1(new_n467), .C2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT87), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n759), .B1(new_n766), .B2(new_n678), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT88), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2072), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n690), .B2(new_n689), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n749), .A2(new_n750), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT91), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n758), .B1(new_n773), .B2(KEYINPUT92), .ZN(new_n774));
  NOR2_X1   g349(.A1(G16), .A2(G23), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT86), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G288), .B2(new_n673), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT33), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1976), .ZN(new_n779));
  MUX2_X1   g354(.A(G6), .B(G305), .S(G16), .Z(new_n780));
  XOR2_X1   g355(.A(KEYINPUT32), .B(G1981), .Z(new_n781));
  XOR2_X1   g356(.A(new_n780), .B(new_n781), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n673), .A2(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G166), .B2(new_n673), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1971), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n779), .A2(new_n782), .A3(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT34), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n678), .A2(G25), .ZN(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n791));
  INV_X1    g366(.A(G107), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(G2105), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT85), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G131), .B2(new_n601), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n490), .A2(G119), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n790), .B1(new_n798), .B2(new_n678), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT35), .B(G1991), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  MUX2_X1   g376(.A(G24), .B(G290), .S(G16), .Z(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(G1986), .Z(new_n803));
  NAND4_X1  g378(.A1(new_n788), .A2(new_n789), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT36), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n773), .A2(KEYINPUT92), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n774), .A2(new_n807), .ZN(G311));
  XNOR2_X1  g383(.A(G311), .B(KEYINPUT94), .ZN(G150));
  NAND2_X1  g384(.A1(new_n583), .A2(G559), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT38), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(new_n513), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n518), .A2(G55), .ZN(new_n814));
  INV_X1    g389(.A(G93), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n521), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n550), .B(new_n817), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n811), .B(new_n818), .Z(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n820));
  INV_X1    g395(.A(G860), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n817), .A2(new_n821), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT95), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT37), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT96), .ZN(G145));
  XNOR2_X1  g403(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT99), .B(G37), .Z(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n742), .A2(new_n745), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT90), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n735), .A2(new_n737), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(new_n739), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT97), .ZN(new_n838));
  INV_X1    g413(.A(new_n719), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n487), .B(KEYINPUT69), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n838), .B(new_n839), .C1(new_n840), .C2(new_n714), .ZN(new_n841));
  OAI21_X1  g416(.A(KEYINPUT97), .B1(new_n715), .B2(new_n719), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n841), .A2(new_n842), .A3(G164), .ZN(new_n843));
  AOI21_X1  g418(.A(G164), .B1(new_n841), .B2(new_n842), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n837), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n490), .A2(G128), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n838), .B1(new_n846), .B2(new_n839), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n715), .A2(KEYINPUT97), .A3(new_n719), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n507), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n841), .A2(new_n842), .A3(G164), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n849), .A2(new_n747), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n845), .A2(new_n851), .A3(new_n766), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n835), .B1(new_n843), .B2(new_n844), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n849), .A2(new_n833), .A3(new_n850), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n853), .A2(new_n854), .A3(new_n765), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n852), .A2(new_n855), .A3(new_n797), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n797), .B1(new_n852), .B2(new_n855), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n611), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n852), .A2(new_n855), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n798), .ZN(new_n860));
  INV_X1    g435(.A(new_n611), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n852), .A2(new_n855), .A3(new_n797), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(G106), .A2(G2105), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n864), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n865));
  INV_X1    g440(.A(G142), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n469), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n490), .B2(G130), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n858), .A2(new_n863), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n868), .B1(new_n858), .B2(new_n863), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n604), .B(G160), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(G162), .Z(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n832), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n876));
  INV_X1    g451(.A(new_n868), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n856), .A2(new_n857), .A3(new_n611), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n861), .B1(new_n860), .B2(new_n862), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n858), .A2(new_n863), .A3(new_n868), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT98), .B1(new_n882), .B2(new_n873), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n884));
  AOI211_X1 g459(.A(new_n884), .B(new_n874), .C1(new_n880), .C2(new_n881), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n875), .B(new_n876), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n873), .B1(new_n869), .B2(new_n870), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n884), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n882), .A2(KEYINPUT98), .A3(new_n873), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n876), .B1(new_n891), .B2(new_n875), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n830), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n875), .B1(new_n883), .B2(new_n885), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT100), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(new_n886), .A3(new_n829), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(G395));
  XNOR2_X1  g472(.A(new_n595), .B(new_n818), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n578), .A2(new_n582), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(G299), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT41), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n902), .B1(new_n900), .B2(new_n898), .ZN(new_n903));
  XOR2_X1   g478(.A(G303), .B(KEYINPUT102), .Z(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(G290), .ZN(new_n905));
  INV_X1    g480(.A(G288), .ZN(new_n906));
  XNOR2_X1  g481(.A(G305), .B(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n905), .B(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT42), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n903), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(G868), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(G868), .B2(new_n817), .ZN(G295));
  OAI21_X1  g487(.A(new_n911), .B1(G868), .B2(new_n817), .ZN(G331));
  XNOR2_X1  g488(.A(new_n818), .B(G301), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(G168), .ZN(new_n915));
  INV_X1    g490(.A(new_n900), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n901), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n917), .B1(new_n918), .B2(new_n915), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n832), .B1(new_n919), .B2(new_n908), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n908), .B2(new_n919), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(KEYINPUT43), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n923));
  INV_X1    g498(.A(new_n919), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n908), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(G37), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n919), .A2(new_n925), .A3(new_n908), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n931), .B1(new_n921), .B2(KEYINPUT43), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n927), .A2(new_n923), .A3(new_n928), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n934), .B1(new_n933), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(G397));
  INV_X1    g513(.A(KEYINPUT126), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n720), .B(new_n722), .ZN(new_n940));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n503), .B(KEYINPUT70), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n494), .A2(new_n495), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n498), .A2(new_n500), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n943), .B(new_n944), .C1(new_n469), .C2(new_n492), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n941), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(G160), .A2(G40), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n940), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G1996), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n833), .ZN(new_n954));
  OAI221_X1 g529(.A(new_n951), .B1(new_n953), .B2(new_n837), .C1(new_n952), .C2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n950), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n798), .A2(new_n800), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n798), .A2(new_n800), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(G290), .A2(G1986), .ZN(new_n961));
  AND2_X1   g536(.A1(G290), .A2(G1986), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n950), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT63), .ZN(new_n965));
  XOR2_X1   g540(.A(KEYINPUT105), .B(G1971), .Z(new_n966));
  OAI211_X1 g541(.A(KEYINPUT45), .B(new_n941), .C1(new_n942), .C2(new_n945), .ZN(new_n967));
  INV_X1    g542(.A(G40), .ZN(new_n968));
  NOR4_X1   g543(.A1(new_n471), .A2(new_n475), .A3(new_n968), .A4(new_n477), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT45), .B1(new_n507), .B2(new_n941), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n966), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n946), .A2(KEYINPUT50), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n507), .A2(new_n974), .A3(new_n941), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n973), .A2(new_n969), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n972), .B1(G2090), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(G8), .ZN(new_n978));
  NAND2_X1  g553(.A1(G303), .A2(G8), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT55), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT49), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT107), .B(G1981), .Z(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n570), .A2(new_n571), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1981), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n570), .B2(new_n571), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n982), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n988), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n990), .A2(KEYINPUT49), .A3(new_n985), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n943), .A2(new_n944), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n469), .A2(new_n492), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n503), .B(new_n504), .ZN(new_n995));
  AOI21_X1  g570(.A(G1384), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n969), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n989), .A2(new_n991), .A3(G8), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n906), .A2(G1976), .ZN(new_n999));
  OAI211_X1 g574(.A(G8), .B(new_n999), .C1(new_n946), .C2(new_n949), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT52), .ZN(new_n1001));
  INV_X1    g576(.A(G1976), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT52), .B1(G288), .B2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n997), .A2(G8), .A3(new_n999), .A4(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n998), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n978), .A2(new_n980), .B1(new_n981), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT106), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n972), .A2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT106), .B(new_n966), .C1(new_n970), .C2(new_n971), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1008), .B(new_n1009), .C1(G2090), .C2(new_n976), .ZN(new_n1010));
  INV_X1    g585(.A(new_n980), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(G8), .A3(new_n1011), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1005), .A2(new_n981), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1006), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n710), .B1(new_n970), .B2(new_n971), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT110), .B(new_n710), .C1(new_n970), .C2(new_n971), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n973), .A2(new_n975), .A3(new_n690), .A4(new_n969), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(G8), .B(G168), .C1(new_n1018), .C2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n965), .B1(new_n1014), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1010), .A2(G8), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1022), .B1(new_n1024), .B2(new_n980), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1005), .A2(new_n965), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1012), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n1012), .A2(new_n1005), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT108), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n998), .A2(new_n1002), .A3(new_n906), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1030), .B1(new_n1032), .B2(new_n986), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(KEYINPUT108), .A3(new_n985), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1033), .A2(G8), .A3(new_n997), .A4(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1028), .A2(new_n1029), .A3(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT56), .B(G2072), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n948), .A2(new_n967), .A3(new_n969), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT111), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n949), .B1(new_n996), .B2(KEYINPUT45), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT111), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(new_n948), .A4(new_n1037), .ZN(new_n1042));
  INV_X1    g617(.A(G1956), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n976), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n1046));
  XNOR2_X1  g621(.A(G299), .B(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1047), .A2(new_n1039), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT61), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1045), .A2(KEYINPUT114), .A3(new_n1048), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1053), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n593), .A2(KEYINPUT113), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n970), .A2(new_n971), .A3(G1996), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT58), .B(G1341), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n996), .B2(new_n969), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1057), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT59), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1063), .B(new_n1057), .C1(new_n1058), .C2(new_n1060), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1056), .A2(new_n1051), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT60), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1066), .B1(new_n583), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1348), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n976), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n969), .A2(new_n507), .A3(new_n941), .A4(new_n722), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT112), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n996), .A2(new_n1073), .A3(new_n722), .A4(new_n969), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1068), .A2(new_n1070), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n899), .A2(KEYINPUT115), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1068), .A2(new_n1070), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1070), .A2(new_n1075), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n1066), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT116), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1079), .A2(new_n1082), .A3(new_n1085), .A4(new_n1080), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1055), .A2(new_n1065), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1049), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n899), .B1(new_n1070), .B2(new_n1075), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1051), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT117), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1017), .A2(G168), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(new_n1093), .A3(G8), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1094), .A2(new_n1095), .A3(KEYINPUT51), .ZN(new_n1096));
  OAI211_X1 g671(.A(G8), .B(G286), .C1(new_n1018), .C2(new_n1021), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1092), .A2(KEYINPUT119), .A3(G8), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT51), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1096), .B(new_n1097), .C1(new_n1098), .C2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n948), .A2(new_n698), .A3(new_n967), .A4(new_n969), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G1961), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n976), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1040), .A2(KEYINPUT53), .A3(new_n698), .A4(new_n948), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1103), .B1(new_n1110), .B2(G171), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1105), .A2(new_n1104), .B1(new_n976), .B2(new_n1107), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1104), .A2(KEYINPUT120), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT53), .B1(new_n1104), .B2(KEYINPUT120), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1112), .B(G301), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1111), .A2(KEYINPUT121), .A3(new_n1115), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(G171), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1112), .A2(G301), .A3(new_n1109), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT54), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1124), .A2(new_n1014), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1102), .A2(new_n1120), .A3(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1091), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1087), .A2(KEYINPUT117), .A3(new_n1090), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1036), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1102), .A2(KEYINPUT62), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT122), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1102), .A2(KEYINPUT62), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1102), .A2(new_n1133), .A3(KEYINPUT62), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1014), .A2(new_n1122), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n964), .B1(new_n1129), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n951), .A2(new_n954), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n1138), .B(KEYINPUT125), .Z(new_n1139));
  INV_X1    g714(.A(KEYINPUT46), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n953), .A2(new_n1140), .ZN(new_n1141));
  XOR2_X1   g716(.A(new_n1141), .B(KEYINPUT124), .Z(new_n1142));
  NAND2_X1  g717(.A1(new_n953), .A2(new_n1140), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n1143), .B(KEYINPUT123), .Z(new_n1144));
  NAND3_X1  g719(.A1(new_n1139), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT47), .Z(new_n1146));
  NAND2_X1  g721(.A1(new_n950), .A2(new_n961), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n1147), .B(KEYINPUT48), .Z(new_n1148));
  NOR3_X1   g723(.A1(new_n1148), .A2(new_n955), .A3(new_n959), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n955), .A2(new_n958), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n720), .A2(new_n722), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n956), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1146), .A2(new_n1149), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n939), .B1(new_n1137), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT117), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1102), .A2(new_n1120), .A3(new_n1125), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1158), .A2(new_n1159), .A3(new_n1128), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1036), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1136), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n964), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1164), .A2(KEYINPUT126), .A3(new_n1153), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1155), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g741(.A1(G401), .A2(new_n460), .ZN(new_n1168));
  NAND3_X1  g742(.A1(new_n651), .A2(new_n654), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n1170));
  XNOR2_X1  g744(.A(new_n1169), .B(new_n1170), .ZN(new_n1171));
  INV_X1    g745(.A(G229), .ZN(new_n1172));
  OAI211_X1 g746(.A(new_n1171), .B(new_n1172), .C1(new_n929), .C2(new_n922), .ZN(new_n1173));
  AOI21_X1  g747(.A(new_n1173), .B1(new_n895), .B2(new_n886), .ZN(G308));
  NAND2_X1  g748(.A1(new_n895), .A2(new_n886), .ZN(new_n1175));
  NAND4_X1  g749(.A1(new_n1175), .A2(new_n1172), .A3(new_n930), .A4(new_n1171), .ZN(G225));
endmodule


