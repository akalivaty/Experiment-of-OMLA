//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT84), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G122), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n190), .B(KEYINPUT83), .Z(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  OR2_X1    g006(.A1(KEYINPUT68), .A2(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT68), .A2(G119), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n193), .A2(KEYINPUT69), .A3(G116), .A4(new_n194), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT68), .A2(G119), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT68), .A2(G119), .ZN(new_n197));
  INV_X1    g011(.A(G116), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT69), .B1(new_n198), .B2(G119), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n195), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT2), .B(G113), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G107), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n206), .A2(G107), .ZN(new_n209));
  OAI21_X1  g023(.A(G101), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(new_n206), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G104), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n211), .A2(new_n214), .A3(new_n215), .A4(new_n207), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT5), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n193), .A2(G116), .A3(new_n194), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n200), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n219), .B1(new_n221), .B2(new_n195), .ZN(new_n222));
  OAI21_X1  g036(.A(G113), .B1(new_n220), .B2(KEYINPUT5), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n205), .B(new_n218), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n203), .A3(new_n195), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n203), .B1(new_n221), .B2(new_n195), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n211), .A2(new_n214), .A3(new_n207), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G101), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT4), .A3(new_n216), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT4), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n233), .A3(G101), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n225), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT82), .B1(new_n229), .B2(new_n235), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n192), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n232), .A2(new_n234), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n205), .A2(new_n226), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n237), .A3(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n239), .A2(new_n243), .A3(new_n224), .A4(new_n190), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT6), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n189), .B1(new_n240), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n239), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n224), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n191), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n249), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n244), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT6), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n240), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n253));
  INV_X1    g067(.A(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT64), .A2(G146), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(G143), .A3(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n254), .A2(G143), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT65), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT65), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n257), .A2(new_n263), .A3(new_n259), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(G146), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n255), .A2(new_n256), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(new_n266), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT0), .B(G128), .ZN(new_n270));
  OR2_X1    g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G125), .ZN(new_n273));
  INV_X1    g087(.A(G128), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(KEYINPUT1), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n257), .A2(new_n259), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT67), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT67), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n257), .A2(new_n278), .A3(new_n259), .A4(new_n275), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G125), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n254), .A2(G143), .ZN(new_n282));
  AND2_X1   g096(.A1(KEYINPUT64), .A2(G146), .ZN(new_n283));
  NOR2_X1   g097(.A1(KEYINPUT64), .A2(G146), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n282), .B1(new_n285), .B2(G143), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n285), .B2(G143), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n286), .B1(new_n288), .B2(new_n274), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n280), .A2(new_n281), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n273), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT85), .B(G224), .Z(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(G953), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n291), .B(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n246), .A2(new_n250), .A3(new_n252), .A4(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT87), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n223), .B1(new_n202), .B2(KEYINPUT5), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n217), .B1(new_n297), .B2(new_n228), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n224), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n190), .B(KEYINPUT8), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT7), .B1(new_n292), .B2(G953), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n273), .A2(new_n290), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(new_n273), .B2(new_n290), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT86), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n301), .B(new_n304), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n291), .A2(new_n306), .A3(new_n302), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n296), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  AND3_X1   g124(.A1(new_n280), .A2(new_n281), .A3(new_n289), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n281), .B1(new_n265), .B2(new_n271), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n313), .A2(new_n303), .B1(new_n299), .B2(new_n300), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n302), .B1(new_n311), .B2(new_n312), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT86), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n314), .A2(KEYINPUT87), .A3(new_n308), .A4(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n310), .A2(new_n244), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G902), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n295), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(G210), .B1(G237), .B2(G902), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n295), .A2(new_n318), .A3(new_n319), .A4(new_n321), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n188), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT9), .B(G234), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT77), .ZN(new_n327));
  OAI21_X1  g141(.A(G221), .B1(new_n327), .B2(G902), .ZN(new_n328));
  INV_X1    g142(.A(G469), .ZN(new_n329));
  XNOR2_X1  g143(.A(G110), .B(G140), .ZN(new_n330));
  INV_X1    g144(.A(G953), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n331), .A2(G227), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n330), .B(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G137), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(KEYINPUT11), .A3(G134), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(G134), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G134), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(G137), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n335), .B(new_n337), .C1(new_n339), .C2(KEYINPUT11), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(G131), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n258), .B1(new_n285), .B2(G143), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n278), .B1(new_n343), .B2(new_n275), .ZN(new_n344));
  INV_X1    g158(.A(new_n279), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n274), .B1(new_n282), .B2(KEYINPUT1), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n347), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n257), .A2(new_n259), .ZN(new_n350));
  INV_X1    g164(.A(new_n348), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT78), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n218), .B1(new_n346), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n280), .A2(new_n289), .A3(new_n217), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n342), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT12), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n356), .B(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n289), .B1(new_n344), .B2(new_n345), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT70), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n280), .A2(KEYINPUT70), .A3(new_n289), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n361), .A2(KEYINPUT10), .A3(new_n362), .A4(new_n218), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n354), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n269), .A2(new_n270), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n366), .B1(new_n264), .B2(new_n262), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n241), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n363), .A2(new_n365), .A3(new_n342), .A4(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n333), .B1(new_n358), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n333), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n369), .A2(KEYINPUT79), .A3(new_n372), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n354), .A2(new_n364), .B1(new_n367), .B2(new_n241), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n363), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT80), .B1(new_n375), .B2(new_n341), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n377));
  AOI211_X1 g191(.A(new_n377), .B(new_n342), .C1(new_n374), .C2(new_n363), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n373), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT79), .B1(new_n369), .B2(new_n372), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n371), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT78), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT78), .B1(new_n350), .B2(new_n351), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n217), .B1(new_n386), .B2(new_n280), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n368), .B1(new_n387), .B2(KEYINPUT10), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n280), .A2(KEYINPUT70), .A3(new_n289), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT70), .B1(new_n280), .B2(new_n289), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n218), .A2(KEYINPUT10), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n341), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n377), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n375), .A2(KEYINPUT80), .A3(new_n341), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n380), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(new_n373), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(KEYINPUT81), .A3(new_n371), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n329), .B1(new_n383), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n372), .B1(new_n396), .B2(new_n369), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n369), .A2(new_n372), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n358), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n329), .B(new_n319), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n329), .A2(new_n319), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n325), .B(new_n328), .C1(new_n400), .C2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G237), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(new_n331), .A3(G210), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT27), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT26), .B(G101), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n339), .A2(new_n336), .ZN(new_n415));
  INV_X1    g229(.A(G131), .ZN(new_n416));
  MUX2_X1   g230(.A(new_n415), .B(new_n340), .S(new_n416), .Z(new_n417));
  NAND2_X1  g231(.A1(new_n359), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT66), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n341), .B1(new_n367), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n272), .A2(KEYINPUT66), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n361), .A2(new_n417), .A3(new_n362), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n367), .A2(new_n341), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(KEYINPUT30), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n242), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n229), .A3(new_n426), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n414), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n422), .A2(new_n242), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n429), .ZN(new_n432));
  XOR2_X1   g246(.A(KEYINPUT72), .B(KEYINPUT28), .Z(new_n433));
  INV_X1    g247(.A(KEYINPUT28), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n432), .A2(new_n433), .B1(new_n434), .B2(new_n429), .ZN(new_n435));
  AOI211_X1 g249(.A(KEYINPUT29), .B(new_n430), .C1(new_n414), .C2(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n425), .A2(new_n229), .A3(new_n426), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n229), .B1(new_n425), .B2(new_n426), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT28), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n429), .A2(new_n434), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n439), .A2(KEYINPUT29), .A3(new_n414), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n319), .ZN(new_n442));
  OAI21_X1  g256(.A(G472), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT73), .B1(new_n435), .B2(new_n414), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT73), .ZN(new_n445));
  INV_X1    g259(.A(new_n414), .ZN(new_n446));
  INV_X1    g260(.A(new_n433), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n431), .B2(new_n429), .ZN(new_n448));
  INV_X1    g262(.A(new_n440), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n445), .B(new_n446), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT71), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n429), .A2(new_n451), .A3(new_n414), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n451), .B1(new_n429), .B2(new_n414), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(KEYINPUT31), .B1(new_n454), .B2(new_n428), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT71), .B1(new_n437), .B2(new_n446), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n429), .A2(new_n451), .A3(new_n414), .ZN(new_n457));
  AND4_X1   g271(.A1(KEYINPUT31), .A2(new_n456), .A3(new_n428), .A4(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n444), .B(new_n450), .C1(new_n455), .C2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT32), .ZN(new_n460));
  NOR2_X1   g274(.A1(G472), .A2(G902), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n459), .B2(new_n461), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n443), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(G128), .B1(new_n193), .B2(new_n194), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(KEYINPUT23), .ZN(new_n466));
  NOR2_X1   g280(.A1(G119), .A2(G128), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT68), .B(G119), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n467), .B1(new_n468), .B2(G128), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n466), .B1(KEYINPUT23), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G110), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(G125), .B(G140), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT16), .ZN(new_n474));
  OR3_X1    g288(.A1(new_n281), .A2(KEYINPUT16), .A3(G140), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n254), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n474), .A2(G146), .A3(new_n475), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT24), .B(G110), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n469), .A2(new_n480), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n472), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n285), .A2(new_n473), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g298(.A(KEYINPUT74), .B(G110), .Z(new_n485));
  NAND2_X1  g299(.A1(new_n470), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n469), .A2(new_n480), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT75), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n482), .A2(new_n488), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT75), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT22), .B(G137), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n331), .A2(G221), .A3(G234), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n496), .B(KEYINPUT76), .Z(new_n497));
  NAND3_X1  g311(.A1(new_n490), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n491), .A2(new_n496), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n319), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT25), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n498), .A2(KEYINPUT25), .A3(new_n319), .A4(new_n499), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G217), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(G234), .B2(new_n319), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n498), .A2(new_n499), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n506), .A2(G902), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n507), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G122), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G116), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n198), .A2(G122), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n515), .A3(new_n213), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT93), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT91), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n519), .B1(new_n266), .B2(G128), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n274), .A2(KEYINPUT91), .A3(G143), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n266), .A2(G128), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n338), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n523), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G134), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n518), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT94), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n198), .A2(G122), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n528), .B(new_n515), .C1(new_n529), .C2(KEYINPUT14), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n513), .A2(G116), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT14), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n531), .B1(new_n532), .B2(new_n514), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT94), .B1(new_n515), .B2(KEYINPUT14), .ZN(new_n534));
  OAI211_X1 g348(.A(G107), .B(new_n530), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT95), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n515), .B1(new_n529), .B2(KEYINPUT14), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n540), .A2(KEYINPUT95), .A3(G107), .A4(new_n530), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n527), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G107), .B1(new_n529), .B2(new_n531), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n516), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT90), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n544), .A2(KEYINPUT90), .A3(new_n516), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT13), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n523), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n266), .A2(KEYINPUT13), .A3(G128), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n522), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI22_X1  g367(.A1(KEYINPUT92), .A2(new_n524), .B1(new_n553), .B2(G134), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n549), .B(new_n554), .C1(KEYINPUT92), .C2(new_n524), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n331), .A2(G217), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n327), .A2(new_n556), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n543), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n557), .B1(new_n543), .B2(new_n555), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n319), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT96), .ZN(new_n561));
  INV_X1    g375(.A(G478), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(KEYINPUT15), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT96), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n564), .B(new_n319), .C1(new_n558), .C2(new_n559), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n561), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n559), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n543), .A2(new_n555), .A3(new_n557), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n563), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n569), .A2(KEYINPUT97), .A3(new_n319), .A4(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT97), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(new_n560), .B2(new_n563), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n566), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G952), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(G953), .ZN(new_n576));
  NAND2_X1  g390(.A1(G234), .A2(G237), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(G902), .A3(G953), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT21), .B(G898), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n410), .A2(new_n331), .A3(G214), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n266), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n410), .A2(new_n331), .A3(G143), .A4(G214), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(KEYINPUT18), .A2(G131), .ZN(new_n588));
  OR3_X1    g402(.A1(new_n587), .A2(KEYINPUT89), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n588), .B1(new_n587), .B2(KEYINPUT89), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n483), .B1(new_n254), .B2(new_n473), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(G113), .B(G122), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(new_n206), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n587), .A2(G131), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT17), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n585), .A2(new_n416), .A3(new_n586), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n587), .A2(KEYINPUT17), .A3(G131), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n599), .A2(new_n478), .A3(new_n477), .A4(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n593), .A2(new_n595), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n595), .B1(new_n593), .B2(new_n601), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n319), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(G475), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n473), .B(KEYINPUT19), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n285), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n596), .A2(new_n598), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n609), .A3(new_n478), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n593), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n602), .B1(new_n611), .B2(new_n595), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT20), .ZN(new_n613));
  NOR2_X1   g427(.A1(G475), .A2(G902), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n612), .B2(new_n614), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n606), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n574), .A2(new_n583), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n409), .A2(new_n464), .A3(new_n512), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G101), .ZN(G3));
  AND2_X1   g435(.A1(new_n317), .A2(new_n244), .ZN(new_n622));
  AOI21_X1  g436(.A(G902), .B1(new_n622), .B2(new_n310), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n321), .B1(new_n623), .B2(new_n295), .ZN(new_n624));
  AND4_X1   g438(.A1(new_n319), .A2(new_n295), .A3(new_n318), .A4(new_n321), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n187), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n561), .A2(new_n562), .A3(new_n565), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT98), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n569), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n628), .A2(new_n629), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n567), .B(new_n568), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n319), .A2(G478), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n627), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n618), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n626), .A2(new_n583), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n328), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n398), .A2(KEYINPUT81), .A3(new_n371), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT81), .B1(new_n398), .B2(new_n371), .ZN(new_n641));
  OAI21_X1  g455(.A(G469), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n369), .B1(new_n376), .B2(new_n378), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n333), .ZN(new_n644));
  INV_X1    g458(.A(new_n403), .ZN(new_n645));
  AOI21_X1  g459(.A(G902), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n405), .B1(new_n646), .B2(new_n329), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n639), .B1(new_n642), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(G472), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n459), .B2(new_n319), .ZN(new_n650));
  INV_X1    g464(.A(new_n461), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n272), .A2(KEYINPUT66), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n367), .A2(new_n419), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n653), .A3(new_n341), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n229), .B1(new_n654), .B2(new_n418), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n433), .B1(new_n437), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n440), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n445), .B1(new_n657), .B2(new_n446), .ZN(new_n658));
  INV_X1    g472(.A(new_n450), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n456), .A2(new_n428), .A3(new_n457), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT31), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n454), .A2(KEYINPUT31), .A3(new_n428), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n651), .B1(new_n660), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n650), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n638), .A2(new_n512), .A3(new_n648), .A4(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT34), .B(G104), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G6));
  NAND2_X1  g484(.A1(new_n323), .A2(new_n324), .ZN(new_n671));
  INV_X1    g485(.A(new_n583), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n617), .A2(KEYINPUT99), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n612), .A2(new_n616), .A3(new_n614), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n612), .A2(KEYINPUT99), .A3(new_n616), .A4(new_n614), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n606), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n574), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND4_X1   g493(.A1(new_n187), .A2(new_n671), .A3(new_n672), .A4(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n680), .A2(new_n648), .A3(new_n667), .A4(new_n512), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT100), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT35), .B(G107), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G9));
  NAND2_X1  g498(.A1(new_n490), .A2(new_n493), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n685), .B1(KEYINPUT36), .B2(new_n497), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n497), .A2(KEYINPUT36), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n490), .A2(new_n493), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n510), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n504), .B2(new_n506), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n650), .A2(new_n666), .A3(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n691), .A2(new_n325), .A3(new_n648), .A4(new_n619), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT101), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT37), .B(G110), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G12));
  INV_X1    g509(.A(new_n689), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n507), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(G900), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n579), .B1(new_n581), .B2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n677), .A2(new_n678), .A3(new_n699), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n409), .A2(new_n464), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  XOR2_X1   g517(.A(new_n699), .B(KEYINPUT39), .Z(new_n704));
  AOI21_X1  g518(.A(KEYINPUT104), .B1(new_n648), .B2(new_n704), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n328), .B(new_n704), .C1(new_n400), .C2(new_n407), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(KEYINPUT40), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n648), .A2(KEYINPUT104), .A3(new_n704), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n706), .A2(new_n707), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT40), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n437), .A2(new_n438), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n454), .A2(new_n428), .B1(new_n446), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(G472), .B1(new_n715), .B2(G902), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n716), .B1(new_n462), .B2(new_n463), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT103), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n459), .A2(new_n461), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT32), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT103), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n723), .A3(new_n716), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n718), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n671), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n726), .B1(new_n323), .B2(new_n324), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n561), .A2(new_n563), .A3(new_n565), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n573), .A2(new_n571), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n618), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR4_X1   g547(.A1(new_n730), .A2(new_n188), .A3(new_n697), .A4(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n709), .A2(new_n713), .A3(new_n725), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G143), .ZN(G45));
  NOR3_X1   g550(.A1(new_n690), .A2(new_n637), .A3(new_n699), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n409), .A2(new_n464), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G146), .ZN(G48));
  AOI21_X1  g553(.A(new_n403), .B1(new_n643), .B2(new_n333), .ZN(new_n740));
  OAI21_X1  g554(.A(G469), .B1(new_n740), .B2(G902), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n328), .A3(new_n404), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n464), .A2(new_n638), .A3(new_n512), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NAND4_X1  g560(.A1(new_n464), .A2(new_n512), .A3(new_n680), .A4(new_n743), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  NOR2_X1   g562(.A1(new_n626), .A2(new_n742), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n697), .A2(new_n619), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n464), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G119), .ZN(G21));
  NAND2_X1  g566(.A1(new_n733), .A2(KEYINPUT106), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT106), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n574), .A2(new_n754), .A3(new_n618), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT107), .B1(new_n626), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT107), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n325), .A2(new_n758), .A3(new_n753), .A4(new_n755), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n742), .A2(new_n583), .ZN(new_n761));
  INV_X1    g575(.A(new_n650), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n455), .A2(new_n458), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n414), .B1(new_n439), .B2(new_n440), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n763), .B(new_n461), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n765), .B1(new_n663), .B2(new_n664), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT105), .B1(new_n767), .B2(new_n651), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n761), .A2(new_n512), .A3(new_n762), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n760), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g585(.A(KEYINPUT108), .B(G122), .Z(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G24));
  AOI21_X1  g587(.A(new_n650), .B1(new_n768), .B2(new_n766), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n737), .A3(new_n749), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G125), .ZN(G27));
  NAND3_X1  g590(.A1(new_n323), .A2(new_n187), .A3(new_n324), .ZN(new_n777));
  INV_X1    g591(.A(new_n371), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(new_n379), .B2(new_n380), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT109), .A4(new_n373), .ZN(new_n781));
  AOI211_X1 g595(.A(new_n329), .B(new_n778), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT110), .B1(new_n782), .B2(new_n407), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n369), .A2(new_n372), .ZN(new_n784));
  AOI22_X1  g598(.A1(KEYINPUT79), .A2(new_n784), .B1(new_n394), .B2(new_n395), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT109), .B1(new_n785), .B2(new_n397), .ZN(new_n786));
  INV_X1    g600(.A(new_n781), .ZN(new_n787));
  OAI211_X1 g601(.A(G469), .B(new_n371), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT110), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n789), .A3(new_n404), .A4(new_n406), .ZN(new_n790));
  AOI211_X1 g604(.A(new_n639), .B(new_n777), .C1(new_n783), .C2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT111), .B1(new_n462), .B2(new_n463), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n720), .A2(new_n793), .A3(new_n721), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n794), .A3(new_n443), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n637), .A2(new_n699), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n791), .A2(new_n795), .A3(new_n512), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n783), .A2(new_n790), .ZN(new_n798));
  INV_X1    g612(.A(new_n777), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n328), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n464), .A2(new_n512), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n637), .A2(KEYINPUT42), .A3(new_n699), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n797), .A2(KEYINPUT42), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(KEYINPUT112), .B(G131), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(G33));
  AOI21_X1  g620(.A(new_n511), .B1(new_n722), .B2(new_n443), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n791), .A2(new_n807), .A3(new_n700), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G134), .ZN(G36));
  INV_X1    g623(.A(KEYINPUT45), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n383), .A2(new_n810), .A3(new_n399), .ZN(new_n811));
  AOI211_X1 g625(.A(new_n810), .B(new_n778), .C1(new_n780), .C2(new_n781), .ZN(new_n812));
  OAI211_X1 g626(.A(G469), .B(new_n811), .C1(new_n812), .C2(KEYINPUT113), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n812), .A2(KEYINPUT113), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n406), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT46), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n815), .A2(new_n816), .B1(new_n329), .B2(new_n646), .ZN(new_n817));
  OAI211_X1 g631(.A(KEYINPUT46), .B(new_n406), .C1(new_n813), .C2(new_n814), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n639), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n618), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT114), .B1(new_n636), .B2(new_n820), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n821), .A2(KEYINPUT43), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n636), .A2(new_n820), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT43), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n822), .A2(new_n697), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n667), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(new_n827), .A3(KEYINPUT44), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT44), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n777), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n819), .A2(new_n704), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G137), .ZN(G39));
  INV_X1    g646(.A(new_n464), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n511), .A3(new_n796), .A4(new_n799), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT47), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n836), .B(new_n639), .C1(new_n817), .C2(new_n818), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n815), .A2(new_n816), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n404), .A3(new_n818), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT47), .B1(new_n839), .B2(new_n328), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n835), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g655(.A(KEYINPUT115), .B(G140), .Z(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(G42));
  NAND2_X1  g657(.A1(new_n741), .A2(new_n404), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n328), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n837), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n822), .A2(new_n825), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(new_n774), .A3(new_n512), .A4(new_n579), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n777), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n848), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n730), .A2(new_n188), .A3(new_n743), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT119), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT50), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n718), .A2(new_n724), .ZN(new_n858));
  NOR4_X1   g672(.A1(new_n511), .A2(new_n742), .A3(new_n777), .A4(new_n578), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OR3_X1    g674(.A1(new_n860), .A2(new_n618), .A3(new_n636), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n855), .A2(new_n856), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n579), .A2(new_n850), .A3(new_n743), .A4(new_n799), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n769), .A2(new_n762), .A3(new_n697), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n857), .A2(new_n861), .A3(new_n862), .A4(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n853), .A2(KEYINPUT51), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n749), .ZN(new_n868));
  OAI221_X1 g682(.A(new_n576), .B1(new_n851), .B2(new_n868), .C1(new_n860), .C2(new_n637), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n869), .A2(KEYINPUT121), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(KEYINPUT121), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n863), .A2(new_n512), .A3(new_n795), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT48), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n852), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n866), .B1(new_n846), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n867), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n620), .A2(new_n668), .A3(new_n744), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n747), .B1(new_n760), .B2(new_n770), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n678), .A2(new_n618), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n187), .A2(new_n671), .A3(new_n672), .A4(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(new_n648), .A3(new_n667), .A4(new_n512), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n692), .A2(new_n751), .A3(new_n884), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n880), .A2(new_n881), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n639), .B1(new_n783), .B2(new_n790), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n864), .A2(new_n887), .A3(new_n796), .A4(new_n799), .ZN(new_n888));
  NOR4_X1   g702(.A1(new_n690), .A2(new_n574), .A3(new_n677), .A4(new_n699), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n464), .A2(new_n889), .A3(new_n648), .A4(new_n799), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n808), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n886), .A2(new_n804), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n757), .A2(new_n759), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n697), .A2(new_n699), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n887), .A2(new_n893), .A3(new_n717), .A4(new_n894), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n409), .B(new_n464), .C1(new_n701), .C2(new_n737), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n775), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT52), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT53), .ZN(new_n899));
  OR3_X1    g713(.A1(new_n892), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n896), .A2(new_n775), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(KEYINPUT52), .A3(new_n895), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n903));
  XNOR2_X1  g717(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n897), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n897), .A2(new_n904), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT118), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n892), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n900), .B1(KEYINPUT53), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT54), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n908), .A2(new_n905), .A3(new_n902), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n886), .A2(new_n804), .A3(new_n891), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT53), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n899), .B1(new_n892), .B2(new_n898), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n911), .A2(new_n917), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n879), .A2(new_n918), .B1(G952), .B2(G953), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n823), .A2(new_n188), .A3(new_n639), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT49), .ZN(new_n921));
  INV_X1    g735(.A(new_n844), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n512), .B(new_n920), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT116), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n921), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n924), .A2(new_n858), .A3(new_n730), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n919), .A2(new_n926), .ZN(G75));
  AOI21_X1  g741(.A(new_n319), .B1(new_n914), .B2(new_n915), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT56), .B1(new_n928), .B2(G210), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n246), .A2(new_n250), .A3(new_n252), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n294), .ZN(new_n931));
  XNOR2_X1  g745(.A(KEYINPUT122), .B(KEYINPUT55), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n929), .A2(new_n933), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n331), .A2(G952), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(G51));
  NAND2_X1  g751(.A1(new_n914), .A2(new_n915), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n916), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n405), .B(KEYINPUT57), .Z(new_n940));
  OAI22_X1  g754(.A1(new_n939), .A2(new_n940), .B1(new_n401), .B2(new_n403), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n813), .A2(new_n814), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n928), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n936), .B1(new_n941), .B2(new_n943), .ZN(G54));
  NAND2_X1  g758(.A1(KEYINPUT58), .A2(G475), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT123), .Z(new_n946));
  AND3_X1   g760(.A1(new_n928), .A2(new_n612), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n612), .B1(new_n928), .B2(new_n946), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n947), .A2(new_n948), .A3(new_n936), .ZN(G60));
  INV_X1    g763(.A(new_n634), .ZN(new_n950));
  NAND2_X1  g764(.A1(G478), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT59), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n950), .B1(new_n918), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n936), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n950), .A2(new_n952), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n954), .B1(new_n939), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n953), .A2(new_n956), .ZN(G63));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT60), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n938), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n936), .B1(new_n961), .B2(new_n508), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n959), .B1(new_n914), .B2(new_n915), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n686), .A2(new_n688), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n964), .B1(new_n963), .B2(new_n965), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n962), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n962), .B(KEYINPUT61), .C1(new_n966), .C2(new_n967), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(G66));
  NOR2_X1   g786(.A1(new_n292), .A2(new_n582), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n973), .A2(new_n331), .ZN(new_n974));
  INV_X1    g788(.A(new_n886), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(new_n331), .ZN(new_n976));
  INV_X1    g790(.A(G898), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n930), .B1(new_n977), .B2(G953), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n976), .B(new_n978), .ZN(G69));
  NAND2_X1  g793(.A1(new_n841), .A2(new_n831), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n705), .A2(new_n708), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n637), .B1(new_n678), .B2(new_n618), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n981), .A2(new_n807), .A3(new_n799), .A4(new_n982), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n735), .A2(KEYINPUT62), .A3(new_n901), .ZN(new_n984));
  AOI21_X1  g798(.A(KEYINPUT62), .B1(new_n735), .B2(new_n901), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n331), .B1(new_n980), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n424), .A2(new_n427), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(new_n607), .Z(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n990), .B1(G900), .B2(G953), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n795), .A2(new_n512), .A3(new_n893), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n839), .A2(new_n994), .A3(new_n328), .A4(new_n704), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT125), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n819), .A2(KEYINPUT125), .A3(new_n704), .A4(new_n994), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n797), .A2(KEYINPUT42), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n802), .A2(new_n803), .ZN(new_n1001));
  AND4_X1   g815(.A1(new_n1000), .A2(new_n1001), .A3(new_n901), .A4(new_n808), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n999), .A2(new_n831), .A3(new_n841), .A4(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n993), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n991), .A2(new_n992), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n992), .B1(new_n991), .B2(new_n1004), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n331), .B1(G227), .B2(G900), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  NOR3_X1   g822(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n993), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n841), .A2(new_n831), .A3(new_n1002), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n997), .A2(new_n998), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1010), .B1(new_n1013), .B2(new_n331), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n735), .A2(new_n901), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT62), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n735), .A2(KEYINPUT62), .A3(new_n901), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1019), .A2(new_n831), .A3(new_n841), .A4(new_n983), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n989), .B1(new_n1020), .B2(new_n331), .ZN(new_n1021));
  OAI21_X1  g835(.A(KEYINPUT126), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n991), .A2(new_n1004), .A3(new_n992), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1007), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n1009), .A2(new_n1024), .ZN(G72));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n428), .A2(new_n429), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1029), .A2(new_n446), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1028), .B1(new_n1030), .B2(new_n661), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n910), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT127), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1027), .B1(new_n1003), .B2(new_n975), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1035), .A2(new_n428), .A3(new_n429), .A4(new_n446), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1027), .B1(new_n1020), .B2(new_n975), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1037), .A2(new_n414), .A3(new_n1029), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1036), .A2(new_n1038), .A3(new_n954), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1034), .A2(new_n1039), .ZN(G57));
endmodule


