//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G146), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT64), .B1(new_n189), .B2(G143), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(new_n187), .A3(G146), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n188), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n189), .A2(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n187), .A2(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n194), .A2(new_n198), .ZN(new_n199));
  AOI22_X1  g013(.A1(new_n193), .A2(new_n194), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n190), .A2(new_n192), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n203), .B1(new_n195), .B2(KEYINPUT1), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n204), .A3(new_n195), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n206));
  OAI21_X1  g020(.A(G128), .B1(new_n188), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n197), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n201), .B1(new_n210), .B2(G125), .ZN(new_n211));
  INV_X1    g025(.A(G224), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G953), .ZN(new_n213));
  XOR2_X1   g027(.A(new_n211), .B(new_n213), .Z(new_n214));
  INV_X1    g028(.A(KEYINPUT6), .ZN(new_n215));
  XNOR2_X1  g029(.A(G110), .B(G122), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G107), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT80), .B1(new_n218), .B2(G104), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT80), .ZN(new_n220));
  INV_X1    g034(.A(G104), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G107), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT3), .B1(new_n221), .B2(G107), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n218), .A3(G104), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G101), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n223), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n219), .A2(new_n224), .A3(new_n222), .A4(new_n226), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G101), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(KEYINPUT4), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G116), .B(G119), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT2), .B(G113), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(KEYINPUT66), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n235), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT66), .B1(new_n237), .B2(new_n233), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n235), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n230), .A2(new_n241), .A3(G101), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n232), .A2(new_n236), .A3(new_n240), .A4(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n218), .A2(G104), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n221), .A2(G107), .ZN(new_n245));
  OAI21_X1  g059(.A(G101), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n230), .B2(G101), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT81), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n233), .A2(KEYINPUT5), .ZN(new_n250));
  INV_X1    g064(.A(G116), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n251), .A2(KEYINPUT5), .A3(G119), .ZN(new_n252));
  INV_X1    g066(.A(G113), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n250), .A2(new_n254), .B1(new_n237), .B2(new_n233), .ZN(new_n255));
  OAI211_X1 g069(.A(KEYINPUT81), .B(new_n246), .C1(new_n230), .C2(G101), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n249), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n243), .A2(KEYINPUT85), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT85), .B1(new_n243), .B2(new_n257), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n217), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n243), .A2(new_n257), .A3(new_n216), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n215), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n243), .A2(new_n257), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT85), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n243), .A2(new_n257), .A3(KEYINPUT85), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT6), .B1(new_n267), .B2(new_n217), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n214), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT7), .B1(new_n212), .B2(G953), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n211), .B(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n271), .A2(new_n261), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n216), .B(KEYINPUT8), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n255), .B(KEYINPUT86), .Z(new_n274));
  NAND2_X1  g088(.A1(new_n249), .A2(new_n256), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n255), .B1(new_n229), .B2(new_n246), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n273), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(G902), .B1(new_n272), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n269), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(G210), .B1(G237), .B2(G902), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT87), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n281), .B1(new_n269), .B2(new_n279), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT87), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n269), .A2(new_n281), .A3(new_n279), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n284), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT88), .ZN(new_n290));
  OAI21_X1  g104(.A(G214), .B1(G237), .B2(G902), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n288), .B1(new_n285), .B2(new_n286), .ZN(new_n293));
  AOI211_X1 g107(.A(KEYINPUT87), .B(new_n281), .C1(new_n269), .C2(new_n279), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT88), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G125), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n298), .A2(KEYINPUT16), .A3(G140), .ZN(new_n299));
  NAND2_X1  g113(.A1(KEYINPUT74), .A2(G125), .ZN(new_n300));
  INV_X1    g114(.A(G140), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n300), .B(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n299), .B1(new_n302), .B2(KEYINPUT16), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(new_n189), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n305));
  OAI211_X1 g119(.A(G119), .B(new_n203), .C1(new_n305), .C2(KEYINPUT23), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n305), .B(KEYINPUT23), .C1(new_n203), .C2(G119), .ZN(new_n307));
  XOR2_X1   g121(.A(new_n306), .B(new_n307), .Z(new_n308));
  INV_X1    g122(.A(G110), .ZN(new_n309));
  XOR2_X1   g123(.A(G119), .B(G128), .Z(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT24), .B(G110), .ZN(new_n311));
  OAI22_X1  g125(.A1(new_n308), .A2(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OR2_X1    g126(.A1(new_n304), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT22), .B(G137), .ZN(new_n314));
  INV_X1    g128(.A(G953), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(G221), .A3(G234), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n314), .B(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n310), .A2(new_n311), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(KEYINPUT75), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(new_n309), .B2(new_n308), .ZN(new_n321));
  XNOR2_X1  g135(.A(G125), .B(G140), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n322), .A2(KEYINPUT76), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(KEYINPUT76), .ZN(new_n324));
  AOI21_X1  g138(.A(G146), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n303), .A2(G146), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n313), .B(new_n318), .C1(new_n321), .C2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n321), .A2(new_n328), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n318), .B1(new_n331), .B2(new_n313), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT25), .B1(new_n333), .B2(G902), .ZN(new_n334));
  INV_X1    g148(.A(G217), .ZN(new_n335));
  INV_X1    g149(.A(G902), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n335), .B1(G234), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT25), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n338), .B(new_n336), .C1(new_n330), .C2(new_n332), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n334), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n333), .B(KEYINPUT77), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n337), .A2(G902), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT67), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n209), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G134), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G137), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n347), .A2(G137), .ZN(new_n350));
  OAI21_X1  g164(.A(G131), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT11), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n352), .B1(new_n347), .B2(G137), .ZN(new_n353));
  INV_X1    g167(.A(G137), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(KEYINPUT11), .A3(G134), .ZN(new_n355));
  INV_X1    g169(.A(G131), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n353), .A2(new_n355), .A3(new_n356), .A4(new_n348), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n205), .A2(new_n208), .A3(KEYINPUT67), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n346), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n353), .A2(new_n348), .A3(new_n355), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G131), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n357), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n200), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(KEYINPUT30), .A3(new_n365), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n359), .A2(new_n209), .B1(new_n364), .B2(new_n200), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT65), .B1(new_n367), .B2(KEYINPUT30), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n240), .A2(new_n236), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT65), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT30), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n364), .A2(new_n200), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n358), .B1(new_n208), .B2(new_n205), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n371), .B(new_n372), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n366), .A2(new_n368), .A3(new_n370), .A4(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n361), .A2(new_n365), .A3(new_n369), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT26), .B(G101), .ZN(new_n378));
  INV_X1    g192(.A(G237), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n315), .A3(G210), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n378), .B(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n381), .B(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n376), .A2(new_n377), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT31), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n376), .A2(KEYINPUT31), .A3(new_n377), .A4(new_n383), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n383), .B(KEYINPUT69), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n236), .B(new_n240), .C1(new_n373), .C2(new_n374), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n377), .A2(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(KEYINPUT71), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT28), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n377), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n392), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(new_n377), .B2(new_n390), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(KEYINPUT71), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n389), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n388), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT72), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G472), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n388), .A2(new_n400), .A3(KEYINPUT72), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n403), .A2(new_n404), .A3(new_n336), .A4(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT32), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n405), .A2(new_n336), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n409), .A2(KEYINPUT32), .A3(new_n404), .A4(new_n403), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT29), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n376), .A2(new_n377), .ZN(new_n412));
  INV_X1    g226(.A(new_n383), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n399), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n393), .A3(new_n395), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n411), .B(new_n414), .C1(new_n416), .C2(new_n389), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n361), .A2(new_n365), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(new_n370), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n395), .B1(new_n419), .B2(new_n394), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n383), .A2(KEYINPUT29), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n417), .B(new_n336), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G472), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n408), .A2(new_n410), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT9), .B(G234), .ZN(new_n425));
  OAI21_X1  g239(.A(G221), .B1(new_n425), .B2(G902), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(KEYINPUT78), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n379), .A2(new_n315), .A3(G214), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(new_n187), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G131), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n428), .B(G143), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n356), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT17), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n434), .A2(KEYINPUT91), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(KEYINPUT91), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n429), .A2(KEYINPUT17), .A3(G131), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n435), .A2(new_n304), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G113), .B(G122), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(new_n221), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT18), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n431), .B1(new_n441), .B2(new_n356), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n302), .A2(new_n189), .ZN(new_n443));
  OAI221_X1 g257(.A(new_n442), .B1(new_n430), .B2(new_n441), .C1(new_n325), .C2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n438), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n444), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n323), .A2(new_n324), .ZN(new_n447));
  XOR2_X1   g261(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT19), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n302), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n449), .A2(KEYINPUT90), .A3(new_n189), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n430), .A2(new_n432), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n452), .A2(new_n327), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n449), .A2(new_n189), .A3(new_n451), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n446), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n445), .B1(new_n458), .B2(new_n440), .ZN(new_n459));
  NOR2_X1   g273(.A1(G475), .A2(G902), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT20), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n463), .A3(new_n460), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n315), .A2(G952), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n466), .B1(G234), .B2(G237), .ZN(new_n467));
  NAND2_X1  g281(.A1(G234), .A2(G237), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n468), .A2(G902), .A3(G953), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(G898), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n251), .A2(G122), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n218), .B1(new_n473), .B2(KEYINPUT14), .ZN(new_n474));
  XNOR2_X1  g288(.A(G116), .B(G122), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n187), .A2(G128), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT92), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n203), .A2(G143), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n347), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n347), .B1(new_n478), .B2(new_n479), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n476), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n425), .A2(new_n335), .A3(G953), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(KEYINPUT93), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT93), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n478), .A2(new_n486), .A3(new_n347), .A4(new_n479), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n475), .B(new_n218), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT13), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n478), .A2(new_n490), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n478), .A2(new_n490), .B1(new_n203), .B2(G143), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n347), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n483), .B(new_n484), .C1(new_n489), .C2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT94), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n495), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n483), .B1(new_n489), .B2(new_n493), .ZN(new_n498));
  INV_X1    g312(.A(new_n484), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n496), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G478), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n502), .A2(KEYINPUT15), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n501), .A2(new_n336), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n503), .B1(new_n501), .B2(new_n336), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n445), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n440), .B1(new_n438), .B2(new_n444), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n336), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(G475), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n465), .A2(new_n472), .A3(new_n506), .A4(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G469), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(new_n336), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT84), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT81), .B1(new_n229), .B2(new_n246), .ZN(new_n515));
  INV_X1    g329(.A(new_n256), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n517), .A2(KEYINPUT10), .A3(new_n346), .A4(new_n360), .ZN(new_n518));
  INV_X1    g332(.A(new_n364), .ZN(new_n519));
  INV_X1    g333(.A(new_n205), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n193), .A2(new_n204), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n229), .B(new_n246), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT10), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n232), .A2(new_n200), .A3(new_n242), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n518), .A2(new_n519), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  XOR2_X1   g340(.A(G110), .B(G140), .Z(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT79), .ZN(new_n528));
  INV_X1    g342(.A(G227), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(G953), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n528), .B(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n514), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n346), .A2(KEYINPUT10), .A3(new_n360), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n524), .B(new_n525), .C1(new_n533), .C2(new_n275), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n514), .B(new_n531), .C1(new_n534), .C2(new_n364), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT82), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n538), .B(new_n210), .C1(new_n515), .C2(new_n516), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n522), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n209), .B1(new_n249), .B2(new_n256), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(new_n538), .ZN(new_n542));
  OAI211_X1 g356(.A(KEYINPUT12), .B(new_n364), .C1(new_n540), .C2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT83), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n521), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n247), .B1(new_n546), .B2(new_n205), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n547), .B1(new_n541), .B2(new_n538), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT82), .B1(new_n517), .B2(new_n209), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n550), .A2(KEYINPUT83), .A3(KEYINPUT12), .A4(new_n364), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n364), .B1(new_n540), .B2(new_n542), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT12), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n545), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n537), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n534), .A2(new_n364), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n526), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n531), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(G902), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n513), .B1(new_n561), .B2(new_n512), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n555), .A2(new_n526), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n559), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n526), .A2(new_n557), .A3(new_n531), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(G469), .A3(new_n565), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n427), .B(new_n511), .C1(new_n562), .C2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n297), .A2(new_n344), .A3(new_n424), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(G101), .ZN(G3));
  OAI211_X1 g383(.A(new_n409), .B(new_n403), .C1(KEYINPUT95), .C2(new_n404), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n404), .A2(KEYINPUT95), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n405), .A2(new_n336), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT72), .B1(new_n388), .B2(new_n400), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n570), .A2(new_n344), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n562), .A2(new_n566), .ZN(new_n576));
  INV_X1    g390(.A(new_n427), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n283), .A2(KEYINPUT96), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT96), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n288), .B1(new_n285), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n291), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n459), .A2(new_n463), .A3(new_n460), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n463), .B1(new_n459), .B2(new_n460), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n510), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT98), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n494), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n484), .A2(KEYINPUT97), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(new_n588), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n483), .B(new_n591), .C1(new_n489), .C2(new_n493), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n498), .A2(new_n590), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n589), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT33), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n496), .A2(new_n596), .A3(new_n497), .A4(new_n500), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n502), .A2(G902), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n501), .A2(new_n336), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n502), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n587), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(new_n471), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n579), .A2(new_n584), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT34), .B(G104), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G6));
  INV_X1    g422(.A(new_n587), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n504), .A2(new_n505), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n471), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n579), .A2(new_n584), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT35), .B(G107), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G9));
  NOR2_X1   g429(.A1(new_n318), .A2(KEYINPUT36), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n331), .A2(KEYINPUT99), .A3(new_n313), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT99), .B1(new_n331), .B2(new_n313), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n619), .ZN(new_n621));
  INV_X1    g435(.A(new_n616), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n617), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n620), .A2(new_n623), .A3(new_n343), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n331), .A2(new_n313), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n317), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n329), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n338), .B1(new_n627), .B2(new_n336), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n339), .A2(new_n337), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n624), .B(KEYINPUT100), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT100), .B1(new_n340), .B2(new_n624), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n633), .A2(new_n574), .A3(new_n570), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n297), .A2(new_n634), .A3(new_n567), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT37), .B(G110), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT101), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n635), .B(new_n637), .ZN(G12));
  AOI21_X1  g452(.A(new_n427), .B1(new_n562), .B2(new_n566), .ZN(new_n639));
  INV_X1    g453(.A(new_n467), .ZN(new_n640));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n469), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n611), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n584), .A2(new_n639), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n424), .A2(new_n633), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(new_n203), .ZN(G30));
  XOR2_X1   g463(.A(new_n643), .B(KEYINPUT39), .Z(new_n650));
  OR2_X1    g464(.A1(new_n578), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n651), .A2(KEYINPUT40), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n289), .A2(KEYINPUT38), .ZN(new_n653));
  OR3_X1    g467(.A1(new_n293), .A2(KEYINPUT38), .A3(new_n294), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n340), .A2(new_n624), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n506), .B1(new_n465), .B2(new_n510), .ZN(new_n658));
  AND4_X1   g472(.A1(new_n291), .A2(new_n655), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n651), .A2(KEYINPUT40), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n408), .A2(new_n410), .ZN(new_n661));
  INV_X1    g475(.A(new_n389), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n384), .B1(new_n419), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n336), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(G472), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  AND4_X1   g480(.A1(new_n652), .A2(new_n659), .A3(new_n660), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n187), .ZN(G45));
  NOR2_X1   g482(.A1(new_n604), .A2(new_n644), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n584), .A2(new_n639), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n647), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT102), .B(G146), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G48));
  NAND2_X1  g487(.A1(new_n561), .A2(new_n512), .ZN(new_n674));
  AOI22_X1  g488(.A1(new_n537), .A2(new_n555), .B1(new_n558), .B2(new_n559), .ZN(new_n675));
  OAI21_X1  g489(.A(G469), .B1(new_n675), .B2(G902), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n674), .A2(new_n577), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n583), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n678), .A2(new_n344), .A3(new_n424), .A4(new_n605), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT41), .B(G113), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G15));
  NAND4_X1  g495(.A1(new_n678), .A2(new_n344), .A3(new_n424), .A4(new_n612), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G116), .ZN(G18));
  INV_X1    g497(.A(new_n511), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n678), .A2(new_n424), .A3(new_n684), .A4(new_n633), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT103), .B(G119), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G21));
  OAI211_X1 g501(.A(new_n291), .B(new_n658), .C1(new_n580), .C2(new_n582), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n688), .A2(new_n471), .A3(new_n677), .ZN(new_n689));
  OAI21_X1  g503(.A(G472), .B1(new_n572), .B2(new_n573), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT104), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n692), .B(G472), .C1(new_n572), .C2(new_n573), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n420), .A2(new_n389), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n388), .ZN(new_n695));
  NOR2_X1   g509(.A1(G472), .A2(G902), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n691), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n689), .A2(new_n698), .A3(new_n344), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G122), .ZN(G24));
  NAND4_X1  g514(.A1(new_n691), .A2(new_n656), .A3(new_n693), .A4(new_n697), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI22_X1  g517(.A1(new_n690), .A2(KEYINPUT104), .B1(new_n695), .B2(new_n696), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n704), .A2(KEYINPUT105), .A3(new_n656), .A4(new_n693), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n669), .B(KEYINPUT106), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n678), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G125), .ZN(G27));
  AND2_X1   g523(.A1(new_n424), .A2(new_n344), .ZN(new_n710));
  INV_X1    g524(.A(new_n291), .ZN(new_n711));
  NOR4_X1   g525(.A1(new_n293), .A2(new_n294), .A3(new_n711), .A4(new_n427), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n565), .A2(KEYINPUT107), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n565), .A2(KEYINPUT107), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n563), .A2(new_n559), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G469), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n562), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n710), .A2(new_n707), .A3(KEYINPUT42), .A4(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT42), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n424), .A2(new_n712), .A3(new_n344), .A4(new_n717), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n669), .B(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n720), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT108), .B(G131), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G33));
  INV_X1    g541(.A(new_n645), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n721), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n347), .ZN(G36));
  NAND4_X1  g544(.A1(new_n284), .A2(new_n291), .A3(new_n287), .A4(new_n288), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n600), .A2(new_n602), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n587), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI211_X1 g550(.A(KEYINPUT110), .B(KEYINPUT43), .C1(new_n733), .C2(new_n587), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI211_X1 g552(.A(new_n657), .B(new_n738), .C1(new_n574), .C2(new_n570), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n731), .B1(new_n739), .B2(KEYINPUT44), .ZN(new_n740));
  INV_X1    g554(.A(new_n674), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n713), .A2(new_n714), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n564), .A2(KEYINPUT45), .A3(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n531), .B1(new_n555), .B2(new_n526), .ZN(new_n745));
  INV_X1    g559(.A(new_n565), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n743), .A2(new_n747), .A3(G469), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT109), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n512), .B1(new_n715), .B2(KEYINPUT45), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n751), .A3(new_n747), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n513), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n741), .B1(new_n753), .B2(KEYINPUT46), .ZN(new_n754));
  INV_X1    g568(.A(new_n513), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n751), .B1(new_n750), .B2(new_n747), .ZN(new_n756));
  AND4_X1   g570(.A1(new_n751), .A2(new_n743), .A3(G469), .A4(new_n747), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI211_X1 g574(.A(new_n427), .B(new_n650), .C1(new_n754), .C2(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n740), .B(new_n761), .C1(KEYINPUT44), .C2(new_n739), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT47), .ZN(new_n765));
  OAI211_X1 g579(.A(KEYINPUT46), .B(new_n755), .C1(new_n756), .C2(new_n757), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n674), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n749), .A2(new_n752), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT46), .B1(new_n768), .B2(new_n755), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n577), .B(new_n765), .C1(new_n767), .C2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n764), .A2(KEYINPUT47), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n754), .A2(new_n760), .ZN(new_n773));
  INV_X1    g587(.A(new_n771), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n577), .A3(new_n765), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n587), .A2(new_n603), .A3(new_n643), .ZN(new_n777));
  NOR4_X1   g591(.A1(new_n424), .A2(new_n344), .A3(new_n777), .A4(new_n731), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  NOR2_X1   g594(.A1(G952), .A2(G953), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(KEYINPUT118), .Z(new_n782));
  NAND2_X1  g596(.A1(new_n674), .A2(new_n676), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n712), .A2(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n785), .A2(new_n738), .A3(new_n640), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n706), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n661), .A2(new_n344), .A3(new_n467), .A4(new_n665), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n609), .A2(new_n733), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n788), .A2(new_n785), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n677), .A2(new_n291), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n792), .B1(new_n655), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n793), .A2(new_n653), .A3(new_n654), .A4(KEYINPUT117), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n736), .A2(new_n467), .A3(new_n737), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n798), .A2(new_n344), .A3(new_n698), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n797), .A2(KEYINPUT50), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT50), .B1(new_n797), .B2(new_n799), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n791), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n731), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n427), .B1(new_n754), .B2(new_n760), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n774), .B1(new_n808), .B2(new_n765), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n770), .A2(new_n771), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT115), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n772), .A2(new_n812), .A3(new_n775), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n783), .A2(new_n577), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n807), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n802), .B1(new_n817), .B2(KEYINPUT116), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n772), .A2(new_n812), .A3(new_n775), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n812), .B1(new_n772), .B2(new_n775), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT116), .B1(new_n821), .B2(new_n806), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT51), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n791), .B(KEYINPUT51), .C1(new_n800), .C2(new_n801), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n772), .A2(new_n775), .A3(new_n816), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n806), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n786), .A2(new_n710), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT48), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n788), .A2(new_n604), .A3(new_n785), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n466), .B(new_n832), .C1(new_n678), .C2(new_n799), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n829), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n577), .A2(new_n717), .A3(new_n657), .A4(new_n643), .ZN(new_n835));
  INV_X1    g649(.A(new_n688), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n666), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n647), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n578), .A2(new_n583), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n838), .B(new_n839), .C1(new_n645), .C2(new_n669), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n708), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n647), .B1(new_n646), .B2(new_n670), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n723), .B1(new_n703), .B2(new_n705), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n844), .B1(new_n845), .B2(new_n678), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(KEYINPUT52), .A3(new_n837), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n729), .B1(new_n719), .B2(new_n724), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n568), .A2(new_n635), .A3(new_n679), .A4(new_n682), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n587), .A2(new_n610), .A3(new_n644), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT100), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n656), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(new_n853), .A3(new_n630), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n731), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n855), .A2(new_n424), .A3(new_n639), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n845), .B2(new_n718), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n471), .B1(new_n611), .B2(new_n604), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n579), .A2(new_n297), .A3(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n859), .A2(new_n685), .A3(new_n699), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n849), .A2(new_n850), .A3(new_n857), .A4(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n848), .A2(new_n861), .A3(KEYINPUT53), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT53), .B1(new_n848), .B2(new_n861), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT52), .B1(new_n846), .B2(new_n837), .ZN(new_n867));
  AND4_X1   g681(.A1(KEYINPUT52), .A2(new_n708), .A3(new_n837), .A4(new_n840), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n849), .A2(new_n850), .A3(new_n857), .A4(new_n860), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n848), .A2(new_n861), .A3(KEYINPUT53), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT54), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n834), .B1(new_n865), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n782), .B1(new_n824), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n876));
  INV_X1    g690(.A(new_n734), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n344), .A2(new_n291), .A3(new_n577), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT112), .Z(new_n879));
  AOI211_X1 g693(.A(new_n877), .B(new_n879), .C1(KEYINPUT49), .C2(new_n783), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT113), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n653), .B(new_n654), .C1(KEYINPUT49), .C2(new_n783), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n881), .A2(new_n666), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n875), .A2(new_n876), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n782), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT51), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n821), .A2(KEYINPUT116), .A3(new_n806), .ZN(new_n888));
  INV_X1    g702(.A(new_n802), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n887), .B1(new_n890), .B2(new_n822), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n829), .A2(new_n831), .A3(new_n833), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n864), .B1(new_n862), .B2(new_n863), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n871), .A2(KEYINPUT54), .A3(new_n872), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n886), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT119), .B1(new_n896), .B2(new_n883), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n885), .A2(new_n897), .ZN(G75));
  OAI211_X1 g712(.A(G210), .B(G902), .C1(new_n862), .C2(new_n863), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT56), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n262), .A2(new_n268), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(new_n214), .Z(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT55), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n899), .A2(new_n900), .A3(new_n904), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n315), .A2(G952), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT120), .Z(new_n909));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT121), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n906), .A2(new_n912), .A3(new_n907), .A4(new_n909), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(G51));
  XNOR2_X1  g728(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(new_n513), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n893), .A2(new_n894), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n918));
  INV_X1    g732(.A(new_n675), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n336), .B1(new_n871), .B2(new_n872), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(new_n752), .A3(new_n749), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n917), .A2(new_n919), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(KEYINPUT123), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n908), .B1(new_n923), .B2(new_n925), .ZN(G54));
  NAND3_X1  g740(.A1(new_n921), .A2(KEYINPUT58), .A3(G475), .ZN(new_n927));
  INV_X1    g741(.A(new_n459), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n930), .A3(new_n908), .ZN(G60));
  NAND2_X1  g745(.A1(G478), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT59), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n893), .A2(new_n894), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n598), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n936), .A2(new_n909), .A3(new_n937), .ZN(G63));
  NAND2_X1  g752(.A1(new_n871), .A2(new_n872), .ZN(new_n939));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT60), .Z(new_n941));
  NAND4_X1  g755(.A1(new_n939), .A2(new_n620), .A3(new_n623), .A4(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n939), .A2(new_n941), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n909), .B(new_n942), .C1(new_n943), .C2(new_n342), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(G66));
  NOR3_X1   g760(.A1(new_n470), .A2(new_n212), .A3(new_n315), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n850), .A2(new_n860), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n947), .B1(new_n949), .B2(new_n315), .ZN(new_n950));
  INV_X1    g764(.A(G898), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n902), .B1(new_n951), .B2(G953), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n950), .B(new_n952), .Z(G69));
  NAND3_X1  g767(.A1(new_n366), .A2(new_n368), .A3(new_n375), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n449), .A2(new_n451), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n954), .B(new_n955), .Z(new_n956));
  NAND3_X1  g770(.A1(new_n761), .A2(new_n710), .A3(new_n836), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n849), .A2(new_n846), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n762), .A2(new_n779), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n956), .B1(new_n959), .B2(new_n315), .ZN(new_n960));
  INV_X1    g774(.A(new_n708), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n667), .A2(new_n961), .A3(new_n844), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT62), .ZN(new_n963));
  INV_X1    g777(.A(new_n651), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n611), .A2(new_n604), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT124), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n964), .A2(new_n710), .A3(new_n803), .A4(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n762), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n963), .A2(new_n779), .A3(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT125), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n963), .A2(new_n779), .A3(new_n968), .A4(KEYINPUT125), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n956), .A2(new_n315), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n960), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n315), .B1(G227), .B2(G900), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT126), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n641), .B1(new_n956), .B2(new_n529), .ZN(new_n978));
  OAI22_X1  g792(.A1(new_n975), .A2(new_n977), .B1(new_n315), .B2(new_n978), .ZN(G72));
  NAND2_X1  g793(.A1(new_n412), .A2(new_n383), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n971), .A2(new_n949), .A3(new_n972), .ZN(new_n981));
  NAND2_X1  g795(.A1(G472), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT63), .Z(new_n983));
  AOI21_X1  g797(.A(new_n980), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n983), .B1(new_n959), .B2(new_n948), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n985), .A2(new_n377), .A3(new_n413), .A4(new_n376), .ZN(new_n986));
  INV_X1    g800(.A(new_n983), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(new_n414), .B2(new_n384), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT127), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n939), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n986), .B(new_n990), .C1(G952), .C2(new_n315), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n984), .A2(new_n991), .ZN(G57));
endmodule


