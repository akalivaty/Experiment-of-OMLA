

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U550 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U551 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U552 ( .A1(G543), .A2(G651), .ZN(n651) );
  AND2_X1 U553 ( .A1(n695), .A2(n694), .ZN(n514) );
  XOR2_X1 U554 ( .A(n725), .B(KEYINPUT100), .Z(n515) );
  AND2_X1 U555 ( .A1(n808), .A2(n807), .ZN(n516) );
  AND2_X1 U556 ( .A1(n719), .A2(G1996), .ZN(n693) );
  INV_X1 U557 ( .A(n940), .ZN(n698) );
  NAND2_X1 U558 ( .A1(n515), .A2(n734), .ZN(n745) );
  XNOR2_X1 U559 ( .A(KEYINPUT32), .B(n743), .ZN(n762) );
  NAND2_X1 U560 ( .A1(n784), .A2(n690), .ZN(n735) );
  NOR2_X1 U561 ( .A1(G164), .A2(G1384), .ZN(n784) );
  NAND2_X1 U562 ( .A1(n816), .A2(n516), .ZN(n809) );
  NOR2_X1 U563 ( .A1(n574), .A2(n573), .ZN(n575) );
  OR2_X1 U564 ( .A1(n810), .A2(n809), .ZN(n824) );
  XOR2_X1 U565 ( .A(KEYINPUT1), .B(n547), .Z(n655) );
  NOR2_X1 U566 ( .A1(G651), .A2(n635), .ZN(n646) );
  NAND2_X1 U567 ( .A1(n577), .A2(n576), .ZN(n940) );
  INV_X1 U568 ( .A(G2105), .ZN(n520) );
  AND2_X1 U569 ( .A1(n520), .A2(G2104), .ZN(n885) );
  NAND2_X1 U570 ( .A1(G102), .A2(n885), .ZN(n519) );
  NOR2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  XOR2_X2 U572 ( .A(KEYINPUT17), .B(n517), .Z(n886) );
  NAND2_X1 U573 ( .A1(G138), .A2(n886), .ZN(n518) );
  NAND2_X1 U574 ( .A1(n519), .A2(n518), .ZN(n524) );
  NOR2_X1 U575 ( .A1(G2104), .A2(n520), .ZN(n890) );
  NAND2_X1 U576 ( .A1(G126), .A2(n890), .ZN(n522) );
  AND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n893) );
  NAND2_X1 U578 ( .A1(G114), .A2(n893), .ZN(n521) );
  NAND2_X1 U579 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U580 ( .A1(n524), .A2(n523), .ZN(G164) );
  NAND2_X1 U581 ( .A1(G101), .A2(n885), .ZN(n525) );
  XOR2_X1 U582 ( .A(KEYINPUT64), .B(n525), .Z(n526) );
  XNOR2_X1 U583 ( .A(n526), .B(KEYINPUT23), .ZN(n528) );
  NAND2_X1 U584 ( .A1(G113), .A2(n893), .ZN(n527) );
  AND2_X1 U585 ( .A1(n528), .A2(n527), .ZN(n689) );
  NAND2_X1 U586 ( .A1(G137), .A2(n886), .ZN(n530) );
  NAND2_X1 U587 ( .A1(G125), .A2(n890), .ZN(n529) );
  AND2_X1 U588 ( .A1(n530), .A2(n529), .ZN(n687) );
  AND2_X1 U589 ( .A1(n689), .A2(n687), .ZN(G160) );
  XOR2_X1 U590 ( .A(G2438), .B(G2454), .Z(n532) );
  XNOR2_X1 U591 ( .A(G2435), .B(G2430), .ZN(n531) );
  XNOR2_X1 U592 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U593 ( .A(n533), .B(KEYINPUT104), .Z(n535) );
  XNOR2_X1 U594 ( .A(G1348), .B(G1341), .ZN(n534) );
  XNOR2_X1 U595 ( .A(n535), .B(n534), .ZN(n539) );
  XOR2_X1 U596 ( .A(G2446), .B(G2451), .Z(n537) );
  XNOR2_X1 U597 ( .A(G2443), .B(G2427), .ZN(n536) );
  XNOR2_X1 U598 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U599 ( .A(n539), .B(n538), .Z(n540) );
  AND2_X1 U600 ( .A1(G14), .A2(n540), .ZN(G401) );
  AND2_X1 U601 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U602 ( .A(G132), .ZN(G219) );
  INV_X1 U603 ( .A(G82), .ZN(G220) );
  INV_X1 U604 ( .A(G69), .ZN(G235) );
  INV_X1 U605 ( .A(G57), .ZN(G237) );
  NAND2_X1 U606 ( .A1(n651), .A2(G90), .ZN(n541) );
  XOR2_X1 U607 ( .A(KEYINPUT67), .B(n541), .Z(n543) );
  XOR2_X1 U608 ( .A(G543), .B(KEYINPUT0), .Z(n635) );
  INV_X1 U609 ( .A(G651), .ZN(n546) );
  NOR2_X1 U610 ( .A1(n635), .A2(n546), .ZN(n648) );
  NAND2_X1 U611 ( .A1(n648), .A2(G77), .ZN(n542) );
  NAND2_X1 U612 ( .A1(n543), .A2(n542), .ZN(n545) );
  XNOR2_X1 U613 ( .A(KEYINPUT68), .B(KEYINPUT9), .ZN(n544) );
  XNOR2_X1 U614 ( .A(n545), .B(n544), .ZN(n551) );
  NAND2_X1 U615 ( .A1(n646), .A2(G52), .ZN(n549) );
  NOR2_X1 U616 ( .A1(G543), .A2(n546), .ZN(n547) );
  NAND2_X1 U617 ( .A1(G64), .A2(n655), .ZN(n548) );
  AND2_X1 U618 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U619 ( .A1(n551), .A2(n550), .ZN(G301) );
  XNOR2_X1 U620 ( .A(KEYINPUT76), .B(KEYINPUT6), .ZN(n556) );
  NAND2_X1 U621 ( .A1(n655), .A2(G63), .ZN(n554) );
  NAND2_X1 U622 ( .A1(n646), .A2(G51), .ZN(n552) );
  XOR2_X1 U623 ( .A(KEYINPUT75), .B(n552), .Z(n553) );
  NAND2_X1 U624 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U625 ( .A(n556), .B(n555), .Z(n563) );
  XNOR2_X1 U626 ( .A(KEYINPUT74), .B(KEYINPUT5), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n651), .A2(G89), .ZN(n557) );
  XNOR2_X1 U628 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U629 ( .A1(G76), .A2(n648), .ZN(n558) );
  NAND2_X1 U630 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U631 ( .A(n561), .B(n560), .ZN(n562) );
  NAND2_X1 U632 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n564), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U634 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U636 ( .A(n565), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U637 ( .A(G223), .ZN(n826) );
  NAND2_X1 U638 ( .A1(n826), .A2(G567), .ZN(n566) );
  XOR2_X1 U639 ( .A(KEYINPUT11), .B(n566), .Z(G234) );
  XNOR2_X1 U640 ( .A(KEYINPUT71), .B(KEYINPUT13), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n651), .A2(G81), .ZN(n567) );
  XNOR2_X1 U642 ( .A(n567), .B(KEYINPUT12), .ZN(n569) );
  NAND2_X1 U643 ( .A1(G68), .A2(n648), .ZN(n568) );
  NAND2_X1 U644 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U645 ( .A(n571), .B(n570), .ZN(n574) );
  NAND2_X1 U646 ( .A1(n655), .A2(G56), .ZN(n572) );
  XOR2_X1 U647 ( .A(KEYINPUT14), .B(n572), .Z(n573) );
  XNOR2_X1 U648 ( .A(n575), .B(KEYINPUT72), .ZN(n577) );
  NAND2_X1 U649 ( .A1(G43), .A2(n646), .ZN(n576) );
  INV_X1 U650 ( .A(G860), .ZN(n599) );
  OR2_X1 U651 ( .A1(n940), .A2(n599), .ZN(G153) );
  NAND2_X1 U652 ( .A1(G92), .A2(n651), .ZN(n579) );
  NAND2_X1 U653 ( .A1(G79), .A2(n648), .ZN(n578) );
  NAND2_X1 U654 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U655 ( .A1(G54), .A2(n646), .ZN(n581) );
  NAND2_X1 U656 ( .A1(G66), .A2(n655), .ZN(n580) );
  NAND2_X1 U657 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U659 ( .A(KEYINPUT15), .B(n584), .Z(n948) );
  NOR2_X1 U660 ( .A1(n948), .A2(G868), .ZN(n585) );
  XNOR2_X1 U661 ( .A(n585), .B(KEYINPUT73), .ZN(n587) );
  NAND2_X1 U662 ( .A1(G868), .A2(G301), .ZN(n586) );
  NAND2_X1 U663 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G53), .A2(n646), .ZN(n589) );
  NAND2_X1 U665 ( .A1(G65), .A2(n655), .ZN(n588) );
  NAND2_X1 U666 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U667 ( .A(KEYINPUT70), .B(n590), .ZN(n593) );
  NAND2_X1 U668 ( .A1(G78), .A2(n648), .ZN(n591) );
  XNOR2_X1 U669 ( .A(KEYINPUT69), .B(n591), .ZN(n592) );
  NOR2_X1 U670 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n651), .A2(G91), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n595), .A2(n594), .ZN(G299) );
  INV_X1 U673 ( .A(G868), .ZN(n596) );
  NOR2_X1 U674 ( .A1(G286), .A2(n596), .ZN(n598) );
  NOR2_X1 U675 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U676 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U677 ( .A1(n599), .A2(G559), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n600), .A2(n948), .ZN(n601) );
  XNOR2_X1 U679 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n940), .ZN(n604) );
  NAND2_X1 U681 ( .A1(n948), .A2(G868), .ZN(n602) );
  NOR2_X1 U682 ( .A1(G559), .A2(n602), .ZN(n603) );
  NOR2_X1 U683 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U684 ( .A1(G123), .A2(n890), .ZN(n605) );
  XOR2_X1 U685 ( .A(KEYINPUT18), .B(n605), .Z(n606) );
  XNOR2_X1 U686 ( .A(n606), .B(KEYINPUT77), .ZN(n608) );
  NAND2_X1 U687 ( .A1(G111), .A2(n893), .ZN(n607) );
  NAND2_X1 U688 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U689 ( .A1(G99), .A2(n885), .ZN(n610) );
  NAND2_X1 U690 ( .A1(G135), .A2(n886), .ZN(n609) );
  NAND2_X1 U691 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U692 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U693 ( .A(KEYINPUT78), .B(n613), .ZN(n995) );
  XOR2_X1 U694 ( .A(G2096), .B(n995), .Z(n614) );
  NOR2_X1 U695 ( .A1(G2100), .A2(n614), .ZN(n615) );
  XNOR2_X1 U696 ( .A(KEYINPUT79), .B(n615), .ZN(G156) );
  NAND2_X1 U697 ( .A1(n948), .A2(G559), .ZN(n666) );
  XNOR2_X1 U698 ( .A(n940), .B(n666), .ZN(n616) );
  NOR2_X1 U699 ( .A1(n616), .A2(G860), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G93), .A2(n651), .ZN(n618) );
  NAND2_X1 U701 ( .A1(G80), .A2(n648), .ZN(n617) );
  NAND2_X1 U702 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U703 ( .A(KEYINPUT80), .B(n619), .ZN(n623) );
  NAND2_X1 U704 ( .A1(G55), .A2(n646), .ZN(n621) );
  NAND2_X1 U705 ( .A1(G67), .A2(n655), .ZN(n620) );
  NAND2_X1 U706 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U707 ( .A1(n623), .A2(n622), .ZN(n669) );
  XNOR2_X1 U708 ( .A(n624), .B(n669), .ZN(G145) );
  NAND2_X1 U709 ( .A1(G88), .A2(n651), .ZN(n626) );
  NAND2_X1 U710 ( .A1(G62), .A2(n655), .ZN(n625) );
  NAND2_X1 U711 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n648), .A2(G75), .ZN(n627) );
  XOR2_X1 U713 ( .A(KEYINPUT82), .B(n627), .Z(n628) );
  NOR2_X1 U714 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n646), .A2(G50), .ZN(n630) );
  NAND2_X1 U716 ( .A1(n631), .A2(n630), .ZN(G303) );
  INV_X1 U717 ( .A(G303), .ZN(G166) );
  NAND2_X1 U718 ( .A1(G49), .A2(n646), .ZN(n633) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n632) );
  NAND2_X1 U720 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U721 ( .A1(n655), .A2(n634), .ZN(n637) );
  NAND2_X1 U722 ( .A1(n635), .A2(G87), .ZN(n636) );
  NAND2_X1 U723 ( .A1(n637), .A2(n636), .ZN(G288) );
  NAND2_X1 U724 ( .A1(G73), .A2(n648), .ZN(n638) );
  XNOR2_X1 U725 ( .A(n638), .B(KEYINPUT2), .ZN(n645) );
  NAND2_X1 U726 ( .A1(G48), .A2(n646), .ZN(n640) );
  NAND2_X1 U727 ( .A1(G86), .A2(n651), .ZN(n639) );
  NAND2_X1 U728 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U729 ( .A1(G61), .A2(n655), .ZN(n641) );
  XNOR2_X1 U730 ( .A(KEYINPUT81), .B(n641), .ZN(n642) );
  NOR2_X1 U731 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U732 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U733 ( .A1(n646), .A2(G47), .ZN(n647) );
  XNOR2_X1 U734 ( .A(n647), .B(KEYINPUT66), .ZN(n650) );
  NAND2_X1 U735 ( .A1(G72), .A2(n648), .ZN(n649) );
  NAND2_X1 U736 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U737 ( .A1(G85), .A2(n651), .ZN(n652) );
  XNOR2_X1 U738 ( .A(KEYINPUT65), .B(n652), .ZN(n653) );
  NOR2_X1 U739 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U740 ( .A1(n655), .A2(G60), .ZN(n656) );
  NAND2_X1 U741 ( .A1(n657), .A2(n656), .ZN(G290) );
  XNOR2_X1 U742 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n659) );
  XNOR2_X1 U743 ( .A(G288), .B(KEYINPUT19), .ZN(n658) );
  XNOR2_X1 U744 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U745 ( .A(n660), .B(G305), .ZN(n663) );
  INV_X1 U746 ( .A(G299), .ZN(n711) );
  XNOR2_X1 U747 ( .A(n711), .B(n669), .ZN(n661) );
  XNOR2_X1 U748 ( .A(n661), .B(n940), .ZN(n662) );
  XNOR2_X1 U749 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U750 ( .A(G166), .B(n664), .ZN(n665) );
  XNOR2_X1 U751 ( .A(n665), .B(G290), .ZN(n833) );
  XNOR2_X1 U752 ( .A(KEYINPUT85), .B(n666), .ZN(n667) );
  XNOR2_X1 U753 ( .A(n833), .B(n667), .ZN(n668) );
  NAND2_X1 U754 ( .A1(n668), .A2(G868), .ZN(n671) );
  OR2_X1 U755 ( .A1(G868), .A2(n669), .ZN(n670) );
  NAND2_X1 U756 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U757 ( .A1(G2084), .A2(G2078), .ZN(n672) );
  XOR2_X1 U758 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U761 ( .A1(n675), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(KEYINPUT86), .B(G44), .ZN(n676) );
  XNOR2_X1 U763 ( .A(n676), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U764 ( .A1(G661), .A2(G483), .ZN(n685) );
  NOR2_X1 U765 ( .A1(G237), .A2(G235), .ZN(n677) );
  NAND2_X1 U766 ( .A1(G120), .A2(n677), .ZN(n678) );
  XNOR2_X1 U767 ( .A(KEYINPUT87), .B(n678), .ZN(n679) );
  NAND2_X1 U768 ( .A1(n679), .A2(G108), .ZN(n830) );
  NAND2_X1 U769 ( .A1(n830), .A2(G567), .ZN(n684) );
  NOR2_X1 U770 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U771 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U772 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U773 ( .A1(G96), .A2(n682), .ZN(n831) );
  NAND2_X1 U774 ( .A1(n831), .A2(G2106), .ZN(n683) );
  NAND2_X1 U775 ( .A1(n684), .A2(n683), .ZN(n909) );
  NOR2_X1 U776 ( .A1(n685), .A2(n909), .ZN(n686) );
  XNOR2_X1 U777 ( .A(n686), .B(KEYINPUT88), .ZN(n829) );
  NAND2_X1 U778 ( .A1(G36), .A2(n829), .ZN(G176) );
  AND2_X1 U779 ( .A1(n687), .A2(G40), .ZN(n688) );
  NAND2_X1 U780 ( .A1(n689), .A2(n688), .ZN(n783) );
  INV_X1 U781 ( .A(n783), .ZN(n690) );
  NAND2_X1 U782 ( .A1(G8), .A2(n735), .ZN(n767) );
  NOR2_X1 U783 ( .A1(G1981), .A2(G305), .ZN(n691) );
  XOR2_X1 U784 ( .A(n691), .B(KEYINPUT24), .Z(n692) );
  NOR2_X1 U785 ( .A1(n767), .A2(n692), .ZN(n772) );
  INV_X1 U786 ( .A(n735), .ZN(n719) );
  XOR2_X1 U787 ( .A(n693), .B(KEYINPUT26), .Z(n695) );
  NAND2_X1 U788 ( .A1(n735), .A2(G1341), .ZN(n694) );
  INV_X1 U789 ( .A(n948), .ZN(n701) );
  NOR2_X1 U790 ( .A1(n719), .A2(G1348), .ZN(n697) );
  NOR2_X1 U791 ( .A1(G2067), .A2(n735), .ZN(n696) );
  NOR2_X1 U792 ( .A1(n697), .A2(n696), .ZN(n702) );
  NAND2_X1 U793 ( .A1(n701), .A2(n702), .ZN(n699) );
  NAND2_X1 U794 ( .A1(n514), .A2(n700), .ZN(n704) );
  OR2_X1 U795 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U797 ( .A(KEYINPUT97), .B(n705), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n719), .A2(G2072), .ZN(n706) );
  XNOR2_X1 U799 ( .A(n706), .B(KEYINPUT27), .ZN(n708) );
  AND2_X1 U800 ( .A1(G1956), .A2(n735), .ZN(n707) );
  NOR2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U802 ( .A1(n712), .A2(n711), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n715) );
  NOR2_X1 U804 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U805 ( .A(n713), .B(KEYINPUT28), .Z(n714) );
  NAND2_X1 U806 ( .A1(n715), .A2(n714), .ZN(n718) );
  XNOR2_X1 U807 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n716) );
  XNOR2_X1 U808 ( .A(n716), .B(KEYINPUT29), .ZN(n717) );
  XOR2_X1 U809 ( .A(n718), .B(n717), .Z(n724) );
  NAND2_X1 U810 ( .A1(G1961), .A2(n735), .ZN(n721) );
  XOR2_X1 U811 ( .A(G2078), .B(KEYINPUT25), .Z(n917) );
  NAND2_X1 U812 ( .A1(n719), .A2(n917), .ZN(n720) );
  NAND2_X1 U813 ( .A1(n721), .A2(n720), .ZN(n726) );
  NOR2_X1 U814 ( .A1(G301), .A2(n726), .ZN(n722) );
  XNOR2_X1 U815 ( .A(KEYINPUT96), .B(n722), .ZN(n723) );
  AND2_X1 U816 ( .A1(G301), .A2(n726), .ZN(n731) );
  NOR2_X1 U817 ( .A1(G1966), .A2(n767), .ZN(n747) );
  NOR2_X1 U818 ( .A1(G2084), .A2(n735), .ZN(n744) );
  NOR2_X1 U819 ( .A1(n747), .A2(n744), .ZN(n727) );
  NAND2_X1 U820 ( .A1(G8), .A2(n727), .ZN(n728) );
  XNOR2_X1 U821 ( .A(KEYINPUT30), .B(n728), .ZN(n729) );
  NOR2_X1 U822 ( .A1(G168), .A2(n729), .ZN(n730) );
  NOR2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U824 ( .A(KEYINPUT31), .B(n732), .ZN(n733) );
  XNOR2_X1 U825 ( .A(n733), .B(KEYINPUT101), .ZN(n734) );
  NAND2_X1 U826 ( .A1(n745), .A2(G286), .ZN(n742) );
  INV_X1 U827 ( .A(G8), .ZN(n740) );
  NOR2_X1 U828 ( .A1(G1971), .A2(n767), .ZN(n737) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U830 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U831 ( .A1(n738), .A2(G303), .ZN(n739) );
  OR2_X1 U832 ( .A1(n740), .A2(n739), .ZN(n741) );
  AND2_X1 U833 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U834 ( .A1(G8), .A2(n744), .ZN(n749) );
  INV_X1 U835 ( .A(n745), .ZN(n746) );
  NOR2_X1 U836 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n749), .A2(n748), .ZN(n763) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n947) );
  INV_X1 U839 ( .A(n767), .ZN(n750) );
  AND2_X1 U840 ( .A1(n947), .A2(n750), .ZN(n752) );
  AND2_X1 U841 ( .A1(n763), .A2(n752), .ZN(n751) );
  NAND2_X1 U842 ( .A1(n762), .A2(n751), .ZN(n756) );
  INV_X1 U843 ( .A(n752), .ZN(n754) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n935) );
  NOR2_X1 U845 ( .A1(G1971), .A2(G303), .ZN(n945) );
  NOR2_X1 U846 ( .A1(n935), .A2(n945), .ZN(n753) );
  OR2_X1 U847 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U848 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U849 ( .A1(KEYINPUT33), .A2(n757), .ZN(n760) );
  NAND2_X1 U850 ( .A1(n935), .A2(KEYINPUT33), .ZN(n758) );
  NOR2_X1 U851 ( .A1(n758), .A2(n767), .ZN(n759) );
  NOR2_X1 U852 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U853 ( .A(G1981), .B(G305), .Z(n932) );
  NAND2_X1 U854 ( .A1(n761), .A2(n932), .ZN(n770) );
  NAND2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n766) );
  NOR2_X1 U856 ( .A1(G2090), .A2(G303), .ZN(n764) );
  NAND2_X1 U857 ( .A1(G8), .A2(n764), .ZN(n765) );
  NAND2_X1 U858 ( .A1(n766), .A2(n765), .ZN(n768) );
  NAND2_X1 U859 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n810) );
  NAND2_X1 U862 ( .A1(G104), .A2(n885), .ZN(n774) );
  NAND2_X1 U863 ( .A1(G140), .A2(n886), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U865 ( .A(KEYINPUT34), .B(n775), .ZN(n781) );
  NAND2_X1 U866 ( .A1(G128), .A2(n890), .ZN(n777) );
  NAND2_X1 U867 ( .A1(G116), .A2(n893), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U869 ( .A(KEYINPUT35), .B(n778), .ZN(n779) );
  XNOR2_X1 U870 ( .A(KEYINPUT91), .B(n779), .ZN(n780) );
  NOR2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U872 ( .A(KEYINPUT36), .B(n782), .Z(n900) );
  XOR2_X1 U873 ( .A(KEYINPUT37), .B(G2067), .Z(n818) );
  AND2_X1 U874 ( .A1(n900), .A2(n818), .ZN(n1001) );
  NOR2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U876 ( .A(KEYINPUT89), .B(n785), .Z(n822) );
  NAND2_X1 U877 ( .A1(n1001), .A2(n822), .ZN(n786) );
  XNOR2_X1 U878 ( .A(n786), .B(KEYINPUT92), .ZN(n816) );
  NOR2_X1 U879 ( .A1(G1986), .A2(G290), .ZN(n811) );
  INV_X1 U880 ( .A(n811), .ZN(n953) );
  NAND2_X1 U881 ( .A1(G1986), .A2(G290), .ZN(n938) );
  NAND2_X1 U882 ( .A1(n953), .A2(n938), .ZN(n787) );
  NAND2_X1 U883 ( .A1(n787), .A2(n822), .ZN(n788) );
  XNOR2_X1 U884 ( .A(n788), .B(KEYINPUT90), .ZN(n808) );
  NAND2_X1 U885 ( .A1(G107), .A2(n893), .ZN(n795) );
  NAND2_X1 U886 ( .A1(G95), .A2(n885), .ZN(n790) );
  NAND2_X1 U887 ( .A1(G119), .A2(n890), .ZN(n789) );
  NAND2_X1 U888 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U889 ( .A1(G131), .A2(n886), .ZN(n791) );
  XNOR2_X1 U890 ( .A(KEYINPUT93), .B(n791), .ZN(n792) );
  NOR2_X1 U891 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U892 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U893 ( .A(n796), .B(KEYINPUT94), .ZN(n870) );
  NAND2_X1 U894 ( .A1(n870), .A2(G1991), .ZN(n806) );
  NAND2_X1 U895 ( .A1(G105), .A2(n885), .ZN(n797) );
  XNOR2_X1 U896 ( .A(n797), .B(KEYINPUT38), .ZN(n804) );
  NAND2_X1 U897 ( .A1(G141), .A2(n886), .ZN(n799) );
  NAND2_X1 U898 ( .A1(G117), .A2(n893), .ZN(n798) );
  NAND2_X1 U899 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U900 ( .A1(G129), .A2(n890), .ZN(n800) );
  XNOR2_X1 U901 ( .A(KEYINPUT95), .B(n800), .ZN(n801) );
  NOR2_X1 U902 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U903 ( .A1(n804), .A2(n803), .ZN(n873) );
  NAND2_X1 U904 ( .A1(G1996), .A2(n873), .ZN(n805) );
  NAND2_X1 U905 ( .A1(n806), .A2(n805), .ZN(n996) );
  NAND2_X1 U906 ( .A1(n996), .A2(n822), .ZN(n807) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n873), .ZN(n992) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n870), .ZN(n997) );
  NOR2_X1 U909 ( .A1(n997), .A2(n811), .ZN(n812) );
  XNOR2_X1 U910 ( .A(n812), .B(KEYINPUT102), .ZN(n813) );
  NOR2_X1 U911 ( .A1(n996), .A2(n813), .ZN(n814) );
  NOR2_X1 U912 ( .A1(n992), .A2(n814), .ZN(n815) );
  XNOR2_X1 U913 ( .A(n815), .B(KEYINPUT39), .ZN(n817) );
  NAND2_X1 U914 ( .A1(n817), .A2(n816), .ZN(n820) );
  NOR2_X1 U915 ( .A1(n818), .A2(n900), .ZN(n819) );
  XNOR2_X1 U916 ( .A(n819), .B(KEYINPUT103), .ZN(n1008) );
  NAND2_X1 U917 ( .A1(n820), .A2(n1008), .ZN(n821) );
  NAND2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U920 ( .A(KEYINPUT40), .B(n825), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U923 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U925 ( .A1(n829), .A2(n828), .ZN(G188) );
  XNOR2_X1 U926 ( .A(G120), .B(KEYINPUT105), .ZN(G236) );
  XOR2_X1 U927 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  INV_X1 U929 ( .A(G108), .ZN(G238) );
  NOR2_X1 U930 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  INV_X1 U932 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U933 ( .A(G171), .B(n948), .ZN(n832) );
  XNOR2_X1 U934 ( .A(n832), .B(G286), .ZN(n834) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n835) );
  NOR2_X1 U936 ( .A1(G37), .A2(n835), .ZN(n836) );
  XOR2_X1 U937 ( .A(KEYINPUT117), .B(n836), .Z(G397) );
  XOR2_X1 U938 ( .A(KEYINPUT41), .B(G1981), .Z(n838) );
  XNOR2_X1 U939 ( .A(G1966), .B(G1956), .ZN(n837) );
  XNOR2_X1 U940 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U941 ( .A(n839), .B(KEYINPUT109), .Z(n841) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n840) );
  XNOR2_X1 U943 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U944 ( .A(G1976), .B(G1971), .Z(n843) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1961), .ZN(n842) );
  XNOR2_X1 U946 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U947 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U948 ( .A(KEYINPUT108), .B(G2474), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(G229) );
  XOR2_X1 U950 ( .A(KEYINPUT42), .B(G2090), .Z(n849) );
  XNOR2_X1 U951 ( .A(G2084), .B(G2078), .ZN(n848) );
  XNOR2_X1 U952 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U953 ( .A(n850), .B(G2100), .Z(n852) );
  XNOR2_X1 U954 ( .A(G2067), .B(G2072), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U956 ( .A(G2096), .B(KEYINPUT43), .Z(n854) );
  XNOR2_X1 U957 ( .A(G2678), .B(KEYINPUT107), .ZN(n853) );
  XNOR2_X1 U958 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U959 ( .A(n856), .B(n855), .Z(G227) );
  NAND2_X1 U960 ( .A1(G112), .A2(n893), .ZN(n857) );
  XNOR2_X1 U961 ( .A(n857), .B(KEYINPUT112), .ZN(n860) );
  NAND2_X1 U962 ( .A1(G136), .A2(n886), .ZN(n858) );
  XOR2_X1 U963 ( .A(KEYINPUT111), .B(n858), .Z(n859) );
  NAND2_X1 U964 ( .A1(n860), .A2(n859), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G124), .A2(n890), .ZN(n861) );
  XNOR2_X1 U966 ( .A(n861), .B(KEYINPUT44), .ZN(n862) );
  XNOR2_X1 U967 ( .A(n862), .B(KEYINPUT110), .ZN(n864) );
  NAND2_X1 U968 ( .A1(G100), .A2(n885), .ZN(n863) );
  NAND2_X1 U969 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U970 ( .A1(n866), .A2(n865), .ZN(G162) );
  XOR2_X1 U971 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n868) );
  XNOR2_X1 U972 ( .A(KEYINPUT116), .B(KEYINPUT115), .ZN(n867) );
  XNOR2_X1 U973 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U974 ( .A(n869), .B(G162), .Z(n872) );
  XNOR2_X1 U975 ( .A(G164), .B(n870), .ZN(n871) );
  XNOR2_X1 U976 ( .A(n872), .B(n871), .ZN(n876) );
  XNOR2_X1 U977 ( .A(G160), .B(n873), .ZN(n874) );
  XNOR2_X1 U978 ( .A(n874), .B(n995), .ZN(n875) );
  XOR2_X1 U979 ( .A(n876), .B(n875), .Z(n899) );
  NAND2_X1 U980 ( .A1(G103), .A2(n885), .ZN(n878) );
  NAND2_X1 U981 ( .A1(G139), .A2(n886), .ZN(n877) );
  NAND2_X1 U982 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U983 ( .A(KEYINPUT114), .B(n879), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G127), .A2(n890), .ZN(n881) );
  NAND2_X1 U985 ( .A1(G115), .A2(n893), .ZN(n880) );
  NAND2_X1 U986 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U987 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  NOR2_X1 U988 ( .A1(n884), .A2(n883), .ZN(n1004) );
  NAND2_X1 U989 ( .A1(G106), .A2(n885), .ZN(n888) );
  NAND2_X1 U990 ( .A1(G142), .A2(n886), .ZN(n887) );
  NAND2_X1 U991 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U992 ( .A(n889), .B(KEYINPUT45), .ZN(n892) );
  NAND2_X1 U993 ( .A1(G130), .A2(n890), .ZN(n891) );
  NAND2_X1 U994 ( .A1(n892), .A2(n891), .ZN(n896) );
  NAND2_X1 U995 ( .A1(G118), .A2(n893), .ZN(n894) );
  XNOR2_X1 U996 ( .A(KEYINPUT113), .B(n894), .ZN(n895) );
  NOR2_X1 U997 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U998 ( .A(n1004), .B(n897), .ZN(n898) );
  XNOR2_X1 U999 ( .A(n899), .B(n898), .ZN(n901) );
  XOR2_X1 U1000 ( .A(n901), .B(n900), .Z(n902) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n902), .ZN(G395) );
  NOR2_X1 U1002 ( .A1(G401), .A2(n909), .ZN(n906) );
  NOR2_X1 U1003 ( .A1(G229), .A2(G227), .ZN(n903) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n903), .ZN(n904) );
  NOR2_X1 U1005 ( .A1(G397), .A2(n904), .ZN(n905) );
  NAND2_X1 U1006 ( .A1(n906), .A2(n905), .ZN(n907) );
  NOR2_X1 U1007 ( .A1(n907), .A2(G395), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(n908), .B(KEYINPUT118), .ZN(G308) );
  INV_X1 U1009 ( .A(G308), .ZN(G225) );
  INV_X1 U1010 ( .A(n909), .ZN(G319) );
  XNOR2_X1 U1011 ( .A(KEYINPUT54), .B(G34), .ZN(n910) );
  XNOR2_X1 U1012 ( .A(n910), .B(KEYINPUT121), .ZN(n911) );
  XNOR2_X1 U1013 ( .A(G2084), .B(n911), .ZN(n928) );
  XNOR2_X1 U1014 ( .A(G2090), .B(G35), .ZN(n926) );
  XOR2_X1 U1015 ( .A(G1991), .B(G25), .Z(n912) );
  NAND2_X1 U1016 ( .A1(n912), .A2(G28), .ZN(n923) );
  XOR2_X1 U1017 ( .A(G2067), .B(G26), .Z(n913) );
  XNOR2_X1 U1018 ( .A(KEYINPUT119), .B(n913), .ZN(n915) );
  XNOR2_X1 U1019 ( .A(G33), .B(G2072), .ZN(n914) );
  NOR2_X1 U1020 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1021 ( .A(KEYINPUT120), .B(n916), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(G1996), .B(G32), .ZN(n919) );
  XNOR2_X1 U1023 ( .A(n917), .B(G27), .ZN(n918) );
  NOR2_X1 U1024 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1025 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1026 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1027 ( .A(KEYINPUT53), .B(n924), .ZN(n925) );
  NOR2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(n929), .B(KEYINPUT122), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(n930), .B(KEYINPUT55), .ZN(n931) );
  NOR2_X1 U1032 ( .A1(G29), .A2(n931), .ZN(n989) );
  XOR2_X1 U1033 ( .A(G16), .B(KEYINPUT56), .Z(n961) );
  XNOR2_X1 U1034 ( .A(G1966), .B(G168), .ZN(n933) );
  NAND2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1036 ( .A(n934), .B(KEYINPUT57), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(G301), .B(G1961), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(n935), .B(KEYINPUT124), .ZN(n936) );
  NOR2_X1 U1039 ( .A1(n937), .A2(n936), .ZN(n939) );
  NAND2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(G1341), .B(n940), .ZN(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n959) );
  INV_X1 U1044 ( .A(n945), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(n948), .B(G1348), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(KEYINPUT123), .B(n949), .ZN(n950) );
  NOR2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n957) );
  NAND2_X1 U1049 ( .A1(G1971), .A2(G303), .ZN(n952) );
  NAND2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(G1956), .B(G299), .ZN(n954) );
  NOR2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n986) );
  XNOR2_X1 U1056 ( .A(G1348), .B(KEYINPUT59), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n962), .B(G4), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(G1956), .B(G20), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(G19), .B(G1341), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1062 ( .A(KEYINPUT125), .B(G1981), .Z(n967) );
  XNOR2_X1 U1063 ( .A(G6), .B(n967), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(KEYINPUT60), .B(n970), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(G1966), .B(G21), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(G5), .B(G1961), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G1986), .B(G24), .ZN(n976) );
  XNOR2_X1 U1071 ( .A(G1971), .B(G22), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n978) );
  XOR2_X1 U1073 ( .A(G1976), .B(G23), .Z(n977) );
  NAND2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1075 ( .A(KEYINPUT58), .B(n979), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1077 ( .A(KEYINPUT61), .B(n982), .Z(n983) );
  NOR2_X1 U1078 ( .A1(G16), .A2(n983), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(KEYINPUT126), .B(n984), .ZN(n985) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(G11), .A2(n987), .ZN(n988) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(n990), .B(KEYINPUT127), .ZN(n1017) );
  INV_X1 U1084 ( .A(G29), .ZN(n1015) );
  XOR2_X1 U1085 ( .A(G2090), .B(G162), .Z(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1087 ( .A(KEYINPUT51), .B(n993), .Z(n1003) );
  XOR2_X1 U1088 ( .A(G160), .B(G2084), .Z(n994) );
  NOR2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1011) );
  XOR2_X1 U1094 ( .A(G2072), .B(n1004), .Z(n1006) );
  XOR2_X1 U1095 ( .A(G164), .B(G2078), .Z(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(KEYINPUT50), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1100 ( .A(KEYINPUT52), .B(n1012), .Z(n1013) );
  NOR2_X1 U1101 ( .A1(KEYINPUT55), .A2(n1013), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1018), .ZN(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
endmodule

