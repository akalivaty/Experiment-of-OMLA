

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772;

  NOR2_X1 U384 ( .A1(n622), .A2(n626), .ZN(n608) );
  INV_X1 U385 ( .A(n623), .ZN(n540) );
  NOR2_X2 U386 ( .A1(n604), .A2(n605), .ZN(n362) );
  NOR2_X1 U387 ( .A1(n383), .A2(n704), .ZN(n523) );
  XNOR2_X1 U388 ( .A(n418), .B(G128), .ZN(n386) );
  XNOR2_X2 U389 ( .A(n445), .B(n444), .ZN(n643) );
  XNOR2_X1 U390 ( .A(n362), .B(KEYINPUT106), .ZN(n607) );
  NAND2_X1 U391 ( .A1(n363), .A2(n633), .ZN(n636) );
  NAND2_X1 U392 ( .A1(n632), .A2(n727), .ZN(n363) );
  NOR2_X1 U393 ( .A1(n688), .A2(n611), .ZN(n617) );
  AND2_X2 U394 ( .A1(n610), .A2(n609), .ZN(n688) );
  AND2_X1 U395 ( .A1(n381), .A2(n379), .ZN(n378) );
  INV_X2 U396 ( .A(G953), .ZN(n480) );
  NAND2_X1 U397 ( .A1(n628), .A2(n677), .ZN(n570) );
  AND2_X1 U398 ( .A1(n391), .A2(n390), .ZN(n364) );
  AND2_X4 U399 ( .A1(n736), .A2(n735), .ZN(n656) );
  NAND2_X2 U400 ( .A1(n640), .A2(n639), .ZN(n736) );
  INV_X2 U401 ( .A(KEYINPUT64), .ZN(n418) );
  XNOR2_X2 U402 ( .A(n570), .B(n569), .ZN(n650) );
  XNOR2_X2 U403 ( .A(KEYINPUT77), .B(G143), .ZN(n385) );
  XNOR2_X2 U404 ( .A(n519), .B(KEYINPUT35), .ZN(n769) );
  NOR2_X1 U405 ( .A1(n681), .A2(n669), .ZN(n547) );
  XNOR2_X2 U406 ( .A(n587), .B(KEYINPUT1), .ZN(n623) );
  XNOR2_X1 U407 ( .A(KEYINPUT4), .B(G146), .ZN(n755) );
  XNOR2_X1 U408 ( .A(KEYINPUT85), .B(KEYINPUT18), .ZN(n414) );
  NOR2_X1 U409 ( .A1(n556), .A2(n380), .ZN(n379) );
  NOR2_X2 U410 ( .A1(n534), .A2(n574), .ZN(n651) );
  AND2_X1 U411 ( .A1(n402), .A2(n401), .ZN(n400) );
  NOR2_X1 U412 ( .A1(n531), .A2(n526), .ZN(n527) );
  OR2_X1 U413 ( .A1(n543), .A2(KEYINPUT34), .ZN(n401) );
  AND2_X1 U414 ( .A1(n566), .A2(n565), .ZN(n614) );
  XNOR2_X1 U415 ( .A(n532), .B(KEYINPUT6), .ZN(n603) );
  NOR2_X2 U416 ( .A1(G902), .A2(n643), .ZN(n446) );
  XNOR2_X1 U417 ( .A(n415), .B(n414), .ZN(n417) );
  XNOR2_X1 U418 ( .A(G113), .B(G122), .ZN(n421) );
  XNOR2_X1 U419 ( .A(G125), .B(G140), .ZN(n447) );
  BUF_X2 U420 ( .A(n656), .Z(n365) );
  XNOR2_X1 U421 ( .A(n376), .B(KEYINPUT45), .ZN(n366) );
  BUF_X1 U422 ( .A(n738), .Z(n367) );
  BUF_X1 U423 ( .A(n770), .Z(n368) );
  XNOR2_X2 U424 ( .A(n524), .B(KEYINPUT22), .ZN(n531) );
  NAND2_X1 U425 ( .A1(n603), .A2(n477), .ZN(n490) );
  XNOR2_X1 U426 ( .A(n479), .B(n478), .ZN(n758) );
  NAND2_X1 U427 ( .A1(n623), .A2(n406), .ZN(n390) );
  NAND2_X1 U428 ( .A1(n392), .A2(KEYINPUT83), .ZN(n639) );
  AND2_X1 U429 ( .A1(n727), .A2(KEYINPUT2), .ZN(n642) );
  NAND2_X1 U430 ( .A1(n399), .A2(n398), .ZN(n397) );
  AND2_X1 U431 ( .A1(n543), .A2(KEYINPUT34), .ZN(n398) );
  OR2_X1 U432 ( .A1(n659), .A2(G902), .ZN(n489) );
  INV_X1 U433 ( .A(n649), .ZN(n380) );
  XNOR2_X1 U434 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U435 ( .A(G122), .B(KEYINPUT9), .Z(n512) );
  NOR2_X1 U436 ( .A1(n623), .A2(n406), .ZN(n404) );
  INV_X1 U437 ( .A(KEYINPUT88), .ZN(n434) );
  NAND2_X1 U438 ( .A1(n656), .A2(G472), .ZN(n644) );
  NAND2_X1 U439 ( .A1(n656), .A2(G475), .ZN(n396) );
  XNOR2_X1 U440 ( .A(G140), .B(G110), .ZN(n483) );
  NAND2_X1 U441 ( .A1(n737), .A2(n736), .ZN(n389) );
  INV_X1 U442 ( .A(n735), .ZN(n382) );
  XNOR2_X1 U443 ( .A(n530), .B(n529), .ZN(n770) );
  XNOR2_X1 U444 ( .A(n370), .B(n542), .ZN(n681) );
  INV_X1 U445 ( .A(KEYINPUT31), .ZN(n542) );
  INV_X1 U446 ( .A(G110), .ZN(n652) );
  XNOR2_X1 U447 ( .A(n557), .B(n384), .ZN(n533) );
  INV_X1 U448 ( .A(KEYINPUT105), .ZN(n384) );
  XOR2_X1 U449 ( .A(n612), .B(n567), .Z(n369) );
  INV_X1 U450 ( .A(n532), .ZN(n708) );
  NOR2_X1 U451 ( .A1(n712), .A2(n383), .ZN(n370) );
  AND2_X1 U452 ( .A1(G210), .A2(n425), .ZN(n371) );
  XNOR2_X1 U453 ( .A(n657), .B(KEYINPUT59), .ZN(n372) );
  XOR2_X1 U454 ( .A(n367), .B(n413), .Z(n373) );
  INV_X1 U455 ( .A(n742), .ZN(n394) );
  XNOR2_X1 U456 ( .A(KEYINPUT56), .B(KEYINPUT123), .ZN(n374) );
  XNOR2_X1 U457 ( .A(KEYINPUT65), .B(KEYINPUT60), .ZN(n375) );
  XNOR2_X2 U458 ( .A(n376), .B(KEYINPUT45), .ZN(n727) );
  NAND2_X2 U459 ( .A1(n378), .A2(n377), .ZN(n376) );
  NAND2_X1 U460 ( .A1(n535), .A2(n538), .ZN(n377) );
  NAND2_X1 U461 ( .A1(n539), .A2(KEYINPUT44), .ZN(n381) );
  NOR2_X1 U462 ( .A1(n731), .A2(n382), .ZN(n732) );
  NAND2_X1 U463 ( .A1(n642), .A2(n763), .ZN(n735) );
  XNOR2_X1 U464 ( .A(n383), .B(n434), .ZN(n543) );
  XNOR2_X2 U465 ( .A(n433), .B(KEYINPUT0), .ZN(n383) );
  NOR2_X2 U466 ( .A1(n531), .A2(n540), .ZN(n557) );
  XNOR2_X2 U467 ( .A(n510), .B(G131), .ZN(n479) );
  XNOR2_X2 U468 ( .A(n435), .B(G134), .ZN(n510) );
  XNOR2_X2 U469 ( .A(n386), .B(n385), .ZN(n435) );
  XNOR2_X1 U470 ( .A(n387), .B(n374), .ZN(G51) );
  NAND2_X1 U471 ( .A1(n388), .A2(n394), .ZN(n387) );
  XNOR2_X1 U472 ( .A(n389), .B(n373), .ZN(n388) );
  NAND2_X1 U473 ( .A1(n490), .A2(n406), .ZN(n391) );
  NAND2_X1 U474 ( .A1(n638), .A2(n727), .ZN(n392) );
  XNOR2_X1 U475 ( .A(n393), .B(n375), .ZN(G60) );
  NAND2_X1 U476 ( .A1(n395), .A2(n394), .ZN(n393) );
  XNOR2_X1 U477 ( .A(n396), .B(n372), .ZN(n395) );
  NAND2_X1 U478 ( .A1(n400), .A2(n397), .ZN(n518) );
  INV_X1 U479 ( .A(n700), .ZN(n399) );
  NAND2_X1 U480 ( .A1(n700), .A2(n407), .ZN(n402) );
  NAND2_X1 U481 ( .A1(n364), .A2(n403), .ZN(n700) );
  NAND2_X1 U482 ( .A1(n405), .A2(n404), .ZN(n403) );
  INV_X1 U483 ( .A(n490), .ZN(n405) );
  INV_X1 U484 ( .A(KEYINPUT33), .ZN(n406) );
  INV_X1 U485 ( .A(KEYINPUT34), .ZN(n407) );
  XNOR2_X2 U486 ( .A(n408), .B(KEYINPUT19), .ZN(n586) );
  NAND2_X1 U487 ( .A1(n612), .A2(n691), .ZN(n408) );
  XNOR2_X2 U488 ( .A(n409), .B(n371), .ZN(n612) );
  NAND2_X1 U489 ( .A1(n738), .A2(n637), .ZN(n409) );
  NOR2_X2 U490 ( .A1(n770), .A2(n651), .ZN(n538) );
  XOR2_X1 U491 ( .A(n643), .B(KEYINPUT62), .Z(n410) );
  AND2_X1 U492 ( .A1(KEYINPUT78), .A2(n594), .ZN(n411) );
  XOR2_X1 U493 ( .A(G472), .B(KEYINPUT71), .Z(n412) );
  XNOR2_X1 U494 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n413) );
  INV_X1 U495 ( .A(KEYINPUT12), .ZN(n496) );
  XNOR2_X1 U496 ( .A(n499), .B(n498), .ZN(n500) );
  INV_X1 U497 ( .A(KEYINPUT32), .ZN(n529) );
  NAND2_X1 U498 ( .A1(G224), .A2(n480), .ZN(n415) );
  XOR2_X1 U499 ( .A(G125), .B(KEYINPUT17), .Z(n416) );
  XNOR2_X1 U500 ( .A(n417), .B(n416), .ZN(n419) );
  XNOR2_X1 U501 ( .A(n435), .B(n419), .ZN(n420) );
  XNOR2_X1 U502 ( .A(n755), .B(G101), .ZN(n486) );
  XNOR2_X1 U503 ( .A(KEYINPUT3), .B(KEYINPUT70), .ZN(n745) );
  XNOR2_X1 U504 ( .A(n486), .B(n745), .ZN(n436) );
  XNOR2_X1 U505 ( .A(n420), .B(n436), .ZN(n424) );
  XNOR2_X1 U506 ( .A(n652), .B(G119), .ZN(n459) );
  XOR2_X1 U507 ( .A(n459), .B(KEYINPUT16), .Z(n423) );
  XOR2_X1 U508 ( .A(G116), .B(G107), .Z(n513) );
  XNOR2_X1 U509 ( .A(n421), .B(G104), .ZN(n501) );
  XNOR2_X1 U510 ( .A(n513), .B(n501), .ZN(n422) );
  XNOR2_X1 U511 ( .A(n423), .B(n422), .ZN(n743) );
  XNOR2_X1 U512 ( .A(n424), .B(n743), .ZN(n738) );
  XNOR2_X1 U513 ( .A(G902), .B(KEYINPUT15), .ZN(n637) );
  OR2_X1 U514 ( .A1(G237), .A2(G902), .ZN(n425) );
  NAND2_X1 U515 ( .A1(G214), .A2(n425), .ZN(n691) );
  NAND2_X1 U516 ( .A1(G234), .A2(G237), .ZN(n426) );
  XNOR2_X1 U517 ( .A(n426), .B(KEYINPUT86), .ZN(n427) );
  XNOR2_X1 U518 ( .A(KEYINPUT14), .B(n427), .ZN(n428) );
  NAND2_X1 U519 ( .A1(G952), .A2(n428), .ZN(n722) );
  NOR2_X1 U520 ( .A1(G953), .A2(n722), .ZN(n563) );
  AND2_X1 U521 ( .A1(n428), .A2(G953), .ZN(n429) );
  NAND2_X1 U522 ( .A1(G902), .A2(n429), .ZN(n561) );
  NOR2_X1 U523 ( .A1(G898), .A2(n561), .ZN(n430) );
  NOR2_X1 U524 ( .A1(n563), .A2(n430), .ZN(n431) );
  XNOR2_X1 U525 ( .A(KEYINPUT87), .B(n431), .ZN(n432) );
  NAND2_X1 U526 ( .A1(n586), .A2(n432), .ZN(n433) );
  XNOR2_X1 U527 ( .A(n479), .B(n436), .ZN(n445) );
  XOR2_X1 U528 ( .A(G116), .B(KEYINPUT73), .Z(n438) );
  NOR2_X1 U529 ( .A1(G953), .A2(G237), .ZN(n491) );
  NAND2_X1 U530 ( .A1(n491), .A2(G210), .ZN(n437) );
  XNOR2_X1 U531 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U532 ( .A(n439), .B(G137), .Z(n443) );
  XOR2_X1 U533 ( .A(KEYINPUT74), .B(KEYINPUT5), .Z(n441) );
  XNOR2_X1 U534 ( .A(G113), .B(G119), .ZN(n440) );
  XNOR2_X1 U535 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U536 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X2 U537 ( .A(n446), .B(n412), .ZN(n532) );
  XNOR2_X1 U538 ( .A(n447), .B(KEYINPUT10), .ZN(n756) );
  XNOR2_X1 U539 ( .A(n756), .B(G146), .ZN(n492) );
  XNOR2_X1 U540 ( .A(KEYINPUT68), .B(KEYINPUT81), .ZN(n449) );
  NAND2_X1 U541 ( .A1(n480), .A2(G234), .ZN(n448) );
  XNOR2_X1 U542 ( .A(n449), .B(n448), .ZN(n452) );
  INV_X1 U543 ( .A(KEYINPUT8), .ZN(n450) );
  XNOR2_X1 U544 ( .A(n450), .B(KEYINPUT67), .ZN(n451) );
  XNOR2_X1 U545 ( .A(n452), .B(n451), .ZN(n508) );
  NAND2_X1 U546 ( .A1(n508), .A2(G221), .ZN(n453) );
  XNOR2_X1 U547 ( .A(n492), .B(n453), .ZN(n463) );
  XNOR2_X1 U548 ( .A(KEYINPUT24), .B(KEYINPUT91), .ZN(n455) );
  XNOR2_X1 U549 ( .A(KEYINPUT23), .B(KEYINPUT80), .ZN(n454) );
  XNOR2_X1 U550 ( .A(n455), .B(n454), .ZN(n458) );
  XNOR2_X1 U551 ( .A(G128), .B(KEYINPUT90), .ZN(n456) );
  XNOR2_X1 U552 ( .A(n456), .B(KEYINPUT89), .ZN(n457) );
  XNOR2_X1 U553 ( .A(n458), .B(n457), .ZN(n461) );
  XNOR2_X1 U554 ( .A(KEYINPUT69), .B(G137), .ZN(n478) );
  XNOR2_X1 U555 ( .A(n459), .B(n478), .ZN(n460) );
  XNOR2_X1 U556 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U557 ( .A(n463), .B(n462), .ZN(n653) );
  OR2_X1 U558 ( .A1(n653), .A2(G902), .ZN(n471) );
  NAND2_X1 U559 ( .A1(n637), .A2(G234), .ZN(n465) );
  INV_X1 U560 ( .A(KEYINPUT20), .ZN(n464) );
  XNOR2_X1 U561 ( .A(n465), .B(n464), .ZN(n473) );
  INV_X1 U562 ( .A(n473), .ZN(n466) );
  NAND2_X1 U563 ( .A1(n466), .A2(G217), .ZN(n469) );
  XNOR2_X1 U564 ( .A(KEYINPUT75), .B(KEYINPUT92), .ZN(n467) );
  XNOR2_X1 U565 ( .A(n467), .B(KEYINPUT25), .ZN(n468) );
  XNOR2_X1 U566 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X2 U567 ( .A(n471), .B(n470), .ZN(n574) );
  INV_X1 U568 ( .A(G221), .ZN(n472) );
  OR2_X1 U569 ( .A1(n473), .A2(n472), .ZN(n476) );
  INV_X1 U570 ( .A(KEYINPUT93), .ZN(n474) );
  XNOR2_X1 U571 ( .A(n474), .B(KEYINPUT21), .ZN(n475) );
  XNOR2_X1 U572 ( .A(n476), .B(n475), .ZN(n704) );
  INV_X1 U573 ( .A(n704), .ZN(n571) );
  NAND2_X1 U574 ( .A1(n574), .A2(n571), .ZN(n702) );
  INV_X1 U575 ( .A(n702), .ZN(n477) );
  XNOR2_X1 U576 ( .A(G107), .B(G104), .ZN(n482) );
  NAND2_X1 U577 ( .A1(n480), .A2(G227), .ZN(n481) );
  XNOR2_X1 U578 ( .A(n482), .B(n481), .ZN(n484) );
  XNOR2_X1 U579 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U580 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U581 ( .A(n758), .B(n487), .ZN(n659) );
  INV_X1 U582 ( .A(G469), .ZN(n488) );
  XNOR2_X2 U583 ( .A(n489), .B(n488), .ZN(n587) );
  NAND2_X1 U584 ( .A1(G214), .A2(n491), .ZN(n493) );
  XOR2_X1 U585 ( .A(n493), .B(n492), .Z(n503) );
  XOR2_X1 U586 ( .A(KEYINPUT96), .B(KEYINPUT98), .Z(n495) );
  XNOR2_X1 U587 ( .A(G131), .B(KEYINPUT97), .ZN(n494) );
  XNOR2_X1 U588 ( .A(n495), .B(n494), .ZN(n499) );
  XNOR2_X1 U589 ( .A(G143), .B(KEYINPUT11), .ZN(n497) );
  XOR2_X1 U590 ( .A(n501), .B(n500), .Z(n502) );
  XNOR2_X1 U591 ( .A(n503), .B(n502), .ZN(n657) );
  NOR2_X1 U592 ( .A1(n657), .A2(G902), .ZN(n507) );
  XOR2_X1 U593 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n505) );
  XNOR2_X1 U594 ( .A(KEYINPUT13), .B(G475), .ZN(n504) );
  XOR2_X1 U595 ( .A(n505), .B(n504), .Z(n506) );
  XNOR2_X1 U596 ( .A(n507), .B(n506), .ZN(n548) );
  NAND2_X1 U597 ( .A1(n508), .A2(G217), .ZN(n509) );
  XNOR2_X1 U598 ( .A(n510), .B(n509), .ZN(n516) );
  XOR2_X1 U599 ( .A(KEYINPUT7), .B(KEYINPUT102), .Z(n511) );
  XOR2_X1 U600 ( .A(n512), .B(n511), .Z(n514) );
  XNOR2_X1 U601 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U602 ( .A(n516), .B(n515), .ZN(n739) );
  NOR2_X1 U603 ( .A1(G902), .A2(n739), .ZN(n517) );
  XNOR2_X1 U604 ( .A(G478), .B(n517), .ZN(n550) );
  NOR2_X1 U605 ( .A1(n548), .A2(n550), .ZN(n613) );
  NAND2_X1 U606 ( .A1(n518), .A2(n613), .ZN(n519) );
  XNOR2_X1 U607 ( .A(n769), .B(KEYINPUT66), .ZN(n520) );
  NOR2_X1 U608 ( .A1(n520), .A2(KEYINPUT44), .ZN(n535) );
  NAND2_X1 U609 ( .A1(n548), .A2(n550), .ZN(n521) );
  XNOR2_X1 U610 ( .A(KEYINPUT104), .B(n521), .ZN(n693) );
  INV_X1 U611 ( .A(n693), .ZN(n522) );
  NAND2_X1 U612 ( .A1(n523), .A2(n522), .ZN(n524) );
  INV_X1 U613 ( .A(n603), .ZN(n525) );
  INV_X1 U614 ( .A(n574), .ZN(n705) );
  NAND2_X1 U615 ( .A1(n525), .A2(n705), .ZN(n526) );
  XNOR2_X1 U616 ( .A(n540), .B(KEYINPUT84), .ZN(n609) );
  NAND2_X1 U617 ( .A1(n527), .A2(n609), .ZN(n528) );
  XNOR2_X1 U618 ( .A(n528), .B(KEYINPUT76), .ZN(n530) );
  NAND2_X1 U619 ( .A1(n533), .A2(n532), .ZN(n534) );
  INV_X1 U620 ( .A(KEYINPUT66), .ZN(n536) );
  NOR2_X1 U621 ( .A1(n769), .A2(n536), .ZN(n537) );
  NAND2_X1 U622 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U623 ( .A1(n532), .A2(n702), .ZN(n541) );
  NAND2_X1 U624 ( .A1(n541), .A2(n540), .ZN(n712) );
  AND2_X1 U625 ( .A1(n532), .A2(n543), .ZN(n546) );
  OR2_X1 U626 ( .A1(n587), .A2(n702), .ZN(n545) );
  INV_X1 U627 ( .A(KEYINPUT94), .ZN(n544) );
  XNOR2_X1 U628 ( .A(n545), .B(n544), .ZN(n566) );
  AND2_X1 U629 ( .A1(n546), .A2(n566), .ZN(n669) );
  XNOR2_X1 U630 ( .A(n547), .B(KEYINPUT95), .ZN(n554) );
  XNOR2_X1 U631 ( .A(n548), .B(KEYINPUT101), .ZN(n549) );
  AND2_X2 U632 ( .A1(n549), .A2(n550), .ZN(n677) );
  INV_X1 U633 ( .A(n677), .ZN(n553) );
  INV_X1 U634 ( .A(n549), .ZN(n552) );
  INV_X1 U635 ( .A(n550), .ZN(n551) );
  NAND2_X1 U636 ( .A1(n552), .A2(n551), .ZN(n668) );
  NAND2_X1 U637 ( .A1(n553), .A2(n668), .ZN(n695) );
  NAND2_X1 U638 ( .A1(n554), .A2(n695), .ZN(n555) );
  XNOR2_X1 U639 ( .A(n555), .B(KEYINPUT103), .ZN(n556) );
  NOR2_X1 U640 ( .A1(n603), .A2(n705), .ZN(n558) );
  NAND2_X1 U641 ( .A1(n558), .A2(n557), .ZN(n649) );
  NAND2_X1 U642 ( .A1(n708), .A2(n691), .ZN(n560) );
  INV_X1 U643 ( .A(KEYINPUT30), .ZN(n559) );
  XNOR2_X1 U644 ( .A(n560), .B(n559), .ZN(n564) );
  NOR2_X1 U645 ( .A1(G900), .A2(n561), .ZN(n562) );
  OR2_X1 U646 ( .A1(n563), .A2(n562), .ZN(n572) );
  AND2_X1 U647 ( .A1(n564), .A2(n572), .ZN(n565) );
  XNOR2_X1 U648 ( .A(KEYINPUT72), .B(KEYINPUT38), .ZN(n567) );
  NAND2_X1 U649 ( .A1(n614), .A2(n369), .ZN(n568) );
  XNOR2_X2 U650 ( .A(n568), .B(KEYINPUT39), .ZN(n628) );
  INV_X1 U651 ( .A(KEYINPUT40), .ZN(n569) );
  INV_X1 U652 ( .A(n650), .ZN(n583) );
  XOR2_X1 U653 ( .A(KEYINPUT109), .B(KEYINPUT28), .Z(n577) );
  NAND2_X1 U654 ( .A1(n572), .A2(n571), .ZN(n573) );
  OR2_X1 U655 ( .A1(n574), .A2(n573), .ZN(n605) );
  INV_X1 U656 ( .A(n605), .ZN(n575) );
  NAND2_X1 U657 ( .A1(n708), .A2(n575), .ZN(n576) );
  XNOR2_X1 U658 ( .A(n577), .B(n576), .ZN(n590) );
  NOR2_X1 U659 ( .A1(n590), .A2(n587), .ZN(n579) );
  NAND2_X1 U660 ( .A1(n691), .A2(n369), .ZN(n697) );
  NOR2_X1 U661 ( .A1(n693), .A2(n697), .ZN(n578) );
  XOR2_X1 U662 ( .A(KEYINPUT41), .B(n578), .Z(n716) );
  NAND2_X1 U663 ( .A1(n579), .A2(n716), .ZN(n581) );
  INV_X1 U664 ( .A(KEYINPUT42), .ZN(n580) );
  XNOR2_X1 U665 ( .A(n581), .B(n580), .ZN(n772) );
  INV_X1 U666 ( .A(n772), .ZN(n582) );
  NAND2_X1 U667 ( .A1(n583), .A2(n582), .ZN(n585) );
  INV_X1 U668 ( .A(KEYINPUT46), .ZN(n584) );
  XNOR2_X1 U669 ( .A(n585), .B(n584), .ZN(n619) );
  INV_X1 U670 ( .A(n587), .ZN(n588) );
  NAND2_X1 U671 ( .A1(n586), .A2(n588), .ZN(n589) );
  NOR2_X1 U672 ( .A1(n590), .A2(n589), .ZN(n674) );
  INV_X1 U673 ( .A(KEYINPUT78), .ZN(n598) );
  OR2_X1 U674 ( .A1(n674), .A2(n598), .ZN(n593) );
  OR2_X1 U675 ( .A1(n695), .A2(KEYINPUT79), .ZN(n591) );
  AND2_X1 U676 ( .A1(n591), .A2(KEYINPUT47), .ZN(n592) );
  NAND2_X1 U677 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U678 ( .A1(n674), .A2(n695), .ZN(n594) );
  NOR2_X1 U679 ( .A1(KEYINPUT79), .A2(KEYINPUT47), .ZN(n595) );
  NAND2_X1 U680 ( .A1(n411), .A2(n595), .ZN(n596) );
  NAND2_X1 U681 ( .A1(n597), .A2(n596), .ZN(n602) );
  NAND2_X1 U682 ( .A1(n674), .A2(n598), .ZN(n600) );
  NAND2_X1 U683 ( .A1(KEYINPUT79), .A2(n695), .ZN(n599) );
  AND2_X1 U684 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U685 ( .A1(n602), .A2(n601), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n677), .A2(n603), .ZN(n604) );
  NAND2_X1 U687 ( .A1(n607), .A2(n691), .ZN(n622) );
  INV_X1 U688 ( .A(n612), .ZN(n626) );
  XNOR2_X1 U689 ( .A(n608), .B(KEYINPUT36), .ZN(n610) );
  AND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n616), .B(KEYINPUT108), .ZN(n771) );
  AND2_X1 U693 ( .A1(n617), .A2(n771), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n621) );
  INV_X1 U695 ( .A(KEYINPUT48), .ZN(n620) );
  XNOR2_X1 U696 ( .A(n621), .B(n620), .ZN(n631) );
  XNOR2_X1 U697 ( .A(KEYINPUT107), .B(n622), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U699 ( .A(n625), .B(KEYINPUT43), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n627), .A2(n626), .ZN(n690) );
  INV_X1 U701 ( .A(n628), .ZN(n629) );
  OR2_X1 U702 ( .A1(n629), .A2(n668), .ZN(n648) );
  AND2_X1 U703 ( .A1(n690), .A2(n648), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n631), .A2(n630), .ZN(n641) );
  NOR2_X1 U705 ( .A1(KEYINPUT83), .A2(n641), .ZN(n632) );
  INV_X1 U706 ( .A(KEYINPUT2), .ZN(n633) );
  INV_X1 U707 ( .A(n637), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n636), .A2(n635), .ZN(n640) );
  NOR2_X1 U709 ( .A1(n641), .A2(n637), .ZN(n638) );
  INV_X1 U710 ( .A(n641), .ZN(n763) );
  XNOR2_X1 U711 ( .A(n644), .B(n410), .ZN(n646) );
  INV_X1 U712 ( .A(G952), .ZN(n645) );
  AND2_X1 U713 ( .A1(n645), .A2(G953), .ZN(n742) );
  NAND2_X1 U714 ( .A1(n646), .A2(n394), .ZN(n647) );
  XNOR2_X1 U715 ( .A(n647), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U716 ( .A(n648), .B(G134), .ZN(G36) );
  XNOR2_X1 U717 ( .A(n649), .B(G101), .ZN(G3) );
  XOR2_X1 U718 ( .A(G131), .B(n650), .Z(G33) );
  XNOR2_X1 U719 ( .A(n651), .B(n652), .ZN(G12) );
  NAND2_X1 U720 ( .A1(n365), .A2(G217), .ZN(n654) );
  XNOR2_X1 U721 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X1 U722 ( .A1(n655), .A2(n742), .ZN(G66) );
  NAND2_X1 U723 ( .A1(n365), .A2(G469), .ZN(n661) );
  XOR2_X1 U724 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n658) );
  XNOR2_X1 U725 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U726 ( .A(n661), .B(n660), .ZN(n662) );
  NOR2_X1 U727 ( .A1(n662), .A2(n742), .ZN(G54) );
  NAND2_X1 U728 ( .A1(n669), .A2(n677), .ZN(n663) );
  XNOR2_X1 U729 ( .A(n663), .B(KEYINPUT110), .ZN(n664) );
  XNOR2_X1 U730 ( .A(G104), .B(n664), .ZN(G6) );
  XOR2_X1 U731 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n666) );
  XNOR2_X1 U732 ( .A(G107), .B(KEYINPUT111), .ZN(n665) );
  XNOR2_X1 U733 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U734 ( .A(KEYINPUT26), .B(n667), .Z(n671) );
  INV_X1 U735 ( .A(n668), .ZN(n680) );
  NAND2_X1 U736 ( .A1(n669), .A2(n680), .ZN(n670) );
  XNOR2_X1 U737 ( .A(n671), .B(n670), .ZN(G9) );
  XOR2_X1 U738 ( .A(G128), .B(KEYINPUT29), .Z(n673) );
  NAND2_X1 U739 ( .A1(n674), .A2(n680), .ZN(n672) );
  XNOR2_X1 U740 ( .A(n673), .B(n672), .ZN(G30) );
  XOR2_X1 U741 ( .A(G146), .B(KEYINPUT113), .Z(n676) );
  NAND2_X1 U742 ( .A1(n674), .A2(n677), .ZN(n675) );
  XNOR2_X1 U743 ( .A(n676), .B(n675), .ZN(G48) );
  NAND2_X1 U744 ( .A1(n681), .A2(n677), .ZN(n678) );
  XNOR2_X1 U745 ( .A(n678), .B(KEYINPUT114), .ZN(n679) );
  XNOR2_X1 U746 ( .A(G113), .B(n679), .ZN(G15) );
  XOR2_X1 U747 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n683) );
  NAND2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U749 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U750 ( .A(G116), .B(n684), .ZN(G18) );
  XOR2_X1 U751 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n686) );
  XNOR2_X1 U752 ( .A(G125), .B(KEYINPUT37), .ZN(n685) );
  XNOR2_X1 U753 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U754 ( .A(n688), .B(n687), .ZN(G27) );
  XOR2_X1 U755 ( .A(G140), .B(KEYINPUT119), .Z(n689) );
  XNOR2_X1 U756 ( .A(n690), .B(n689), .ZN(G42) );
  NOR2_X1 U757 ( .A1(n369), .A2(n691), .ZN(n692) );
  NOR2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U759 ( .A(n694), .B(KEYINPUT122), .ZN(n699) );
  INV_X1 U760 ( .A(n695), .ZN(n696) );
  NOR2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U762 ( .A1(n699), .A2(n698), .ZN(n701) );
  NOR2_X1 U763 ( .A1(n701), .A2(n700), .ZN(n719) );
  NAND2_X1 U764 ( .A1(n623), .A2(n702), .ZN(n703) );
  XNOR2_X1 U765 ( .A(n703), .B(KEYINPUT50), .ZN(n710) );
  NAND2_X1 U766 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U767 ( .A(n706), .B(KEYINPUT49), .ZN(n707) );
  NOR2_X1 U768 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U770 ( .A(n711), .B(KEYINPUT120), .ZN(n713) );
  NAND2_X1 U771 ( .A1(n713), .A2(n712), .ZN(n715) );
  XOR2_X1 U772 ( .A(KEYINPUT51), .B(KEYINPUT121), .Z(n714) );
  XNOR2_X1 U773 ( .A(n715), .B(n714), .ZN(n717) );
  INV_X1 U774 ( .A(n716), .ZN(n723) );
  NOR2_X1 U775 ( .A1(n717), .A2(n723), .ZN(n718) );
  NOR2_X1 U776 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U777 ( .A(n720), .B(KEYINPUT52), .ZN(n721) );
  NOR2_X1 U778 ( .A1(n722), .A2(n721), .ZN(n725) );
  NOR2_X1 U779 ( .A1(n700), .A2(n723), .ZN(n724) );
  NOR2_X1 U780 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U781 ( .A1(n726), .A2(n480), .ZN(n733) );
  OR2_X1 U782 ( .A1(KEYINPUT2), .A2(n366), .ZN(n728) );
  XNOR2_X1 U783 ( .A(n728), .B(KEYINPUT82), .ZN(n730) );
  NAND2_X1 U784 ( .A1(n641), .A2(n633), .ZN(n729) );
  NAND2_X1 U785 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U786 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U787 ( .A(KEYINPUT53), .B(n734), .ZN(G75) );
  AND2_X1 U788 ( .A1(G210), .A2(n735), .ZN(n737) );
  NAND2_X1 U789 ( .A1(n365), .A2(G478), .ZN(n740) );
  XNOR2_X1 U790 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U791 ( .A1(n742), .A2(n741), .ZN(G63) );
  XOR2_X1 U792 ( .A(G101), .B(n743), .Z(n744) );
  XNOR2_X1 U793 ( .A(n745), .B(n744), .ZN(n747) );
  NOR2_X1 U794 ( .A1(G898), .A2(n480), .ZN(n746) );
  NOR2_X1 U795 ( .A1(n747), .A2(n746), .ZN(n754) );
  NAND2_X1 U796 ( .A1(G224), .A2(G953), .ZN(n748) );
  XNOR2_X1 U797 ( .A(n748), .B(KEYINPUT61), .ZN(n749) );
  XNOR2_X1 U798 ( .A(KEYINPUT124), .B(n749), .ZN(n750) );
  NAND2_X1 U799 ( .A1(G898), .A2(n750), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n366), .A2(n480), .ZN(n751) );
  NAND2_X1 U801 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U802 ( .A(n754), .B(n753), .ZN(G69) );
  XNOR2_X1 U803 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U804 ( .A(n758), .B(n757), .ZN(n762) );
  XNOR2_X1 U805 ( .A(KEYINPUT126), .B(n762), .ZN(n759) );
  XNOR2_X1 U806 ( .A(G227), .B(n759), .ZN(n760) );
  NAND2_X1 U807 ( .A1(n760), .A2(G900), .ZN(n761) );
  NAND2_X1 U808 ( .A1(n761), .A2(G953), .ZN(n767) );
  XNOR2_X1 U809 ( .A(n763), .B(n762), .ZN(n764) );
  NOR2_X1 U810 ( .A1(n764), .A2(G953), .ZN(n765) );
  XNOR2_X1 U811 ( .A(KEYINPUT125), .B(n765), .ZN(n766) );
  NAND2_X1 U812 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U813 ( .A(KEYINPUT127), .B(n768), .Z(G72) );
  XOR2_X1 U814 ( .A(n769), .B(G122), .Z(G24) );
  XOR2_X1 U815 ( .A(G119), .B(n368), .Z(G21) );
  XNOR2_X1 U816 ( .A(G143), .B(n771), .ZN(G45) );
  XOR2_X1 U817 ( .A(G137), .B(n772), .Z(G39) );
endmodule

