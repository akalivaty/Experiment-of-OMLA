//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1261, new_n1262;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT66), .B(KEYINPUT67), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n453), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND3_X1  g034(.A1(new_n453), .A2(KEYINPUT68), .A3(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(G2106), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n462), .B1(new_n452), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n460), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  XNOR2_X1  g043(.A(new_n467), .B(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OR2_X1    g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(G2105), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n476), .A2(G137), .ZN(new_n477));
  INV_X1    g052(.A(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n475), .A2(new_n477), .B1(G101), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n475), .A2(KEYINPUT70), .ZN(new_n488));
  AOI21_X1  g063(.A(G2105), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n476), .B1(new_n487), .B2(new_n488), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n476), .A2(G112), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n490), .B(new_n492), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  XOR2_X1   g070(.A(new_n495), .B(KEYINPUT71), .Z(G162));
  NAND2_X1  g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n471), .B2(new_n472), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(new_n483), .B2(new_n484), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n500), .B(new_n503), .C1(new_n484), .C2(new_n483), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n498), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n506));
  OAI21_X1  g081(.A(G2105), .B1(KEYINPUT72), .B2(G114), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT72), .A2(G114), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n510), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n512), .B(KEYINPUT73), .C1(new_n508), .C2(new_n507), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G50), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n524), .A2(new_n530), .ZN(G166));
  OR2_X1    g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT6), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n518), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n537));
  AOI22_X1  g112(.A1(G51), .A2(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n521), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n525), .A2(G89), .ZN(new_n541));
  NAND2_X1  g116(.A1(G63), .A2(G651), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n539), .A2(new_n543), .ZN(G168));
  NAND2_X1  g119(.A1(new_n534), .A2(G52), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT74), .B(G90), .Z(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n545), .B1(new_n547), .B2(new_n526), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n523), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n548), .A2(new_n550), .ZN(G171));
  NAND2_X1  g126(.A1(new_n534), .A2(G43), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n526), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n521), .A2(G56), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n523), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n540), .B2(new_n565), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n521), .A2(new_n525), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n566), .A2(G651), .B1(new_n567), .B2(G91), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n534), .A2(new_n569), .A3(G53), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  AND2_X1   g146(.A1(KEYINPUT6), .A2(G651), .ZN(new_n572));
  NOR2_X1   g147(.A1(KEYINPUT6), .A2(G651), .ZN(new_n573));
  OAI211_X1 g148(.A(G53), .B(G543), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n575));
  AND3_X1   g150(.A1(new_n570), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n571), .B1(new_n570), .B2(new_n575), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n568), .B1(new_n576), .B2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  INV_X1    g154(.A(G168), .ZN(G286));
  OR2_X1    g155(.A1(new_n524), .A2(new_n530), .ZN(G303));
  NAND2_X1  g156(.A1(new_n567), .A2(G87), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n534), .A2(G49), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n519), .B2(new_n520), .ZN(new_n587));
  AND2_X1   g162(.A1(G73), .A2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n521), .A2(new_n525), .A3(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI211_X1 g167(.A(G48), .B(G543), .C1(new_n572), .C2(new_n573), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT76), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT76), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n525), .A2(new_n595), .A3(G48), .A4(G543), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n592), .A2(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n523), .ZN(new_n600));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT77), .B(G47), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n526), .A2(new_n601), .B1(new_n528), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n534), .A2(G54), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n521), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n523), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n526), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n567), .A2(KEYINPUT10), .A3(G92), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n606), .B1(G868), .B2(new_n614), .ZN(G284));
  OAI21_X1  g190(.A(new_n606), .B1(G868), .B2(new_n614), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G91), .ZN(new_n619));
  OAI22_X1  g194(.A1(new_n618), .A2(new_n523), .B1(new_n619), .B2(new_n526), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n570), .A2(new_n575), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(KEYINPUT75), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n570), .A2(new_n575), .A3(new_n571), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G868), .ZN(G297));
  OAI21_X1  g200(.A(new_n617), .B1(new_n624), .B2(G868), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n614), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n614), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n475), .A2(new_n479), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT13), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2100), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n489), .A2(G135), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n491), .A2(G123), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT78), .ZN(new_n640));
  INV_X1    g215(.A(G111), .ZN(new_n641));
  AOI22_X1  g216(.A1(new_n639), .A2(new_n640), .B1(new_n641), .B2(G2105), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n640), .B2(new_n639), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n637), .A2(new_n638), .A3(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(G2096), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n636), .A2(new_n645), .A3(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(KEYINPUT14), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n653), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  OAI21_X1  g234(.A(G14), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n661), .A2(KEYINPUT79), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(KEYINPUT79), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(KEYINPUT17), .ZN(new_n671));
  INV_X1    g246(.A(new_n665), .ZN(new_n672));
  INV_X1    g247(.A(new_n666), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n668), .A3(new_n673), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(new_n667), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n670), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2096), .B(G2100), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n688));
  INV_X1    g263(.A(new_n685), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n683), .A2(new_n684), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n687), .B(new_n688), .C1(new_n682), .C2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT81), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT82), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n697), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n695), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n699), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n700), .A2(new_n704), .ZN(G229));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G5), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G171), .B2(new_n706), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1961), .ZN(new_n709));
  NOR2_X1   g284(.A1(G16), .A2(G21), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G168), .B2(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G1966), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n713));
  INV_X1    g288(.A(G34), .ZN(new_n714));
  AOI21_X1  g289(.A(G29), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT91), .ZN(new_n717));
  OAI22_X1  g292(.A1(new_n716), .A2(new_n717), .B1(new_n714), .B2(new_n713), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n715), .A2(KEYINPUT91), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  OAI22_X1  g295(.A1(new_n718), .A2(new_n719), .B1(new_n481), .B2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G2084), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n712), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G16), .A2(G19), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n558), .B2(G16), .ZN(new_n725));
  OAI22_X1  g300(.A1(new_n725), .A2(G1341), .B1(new_n644), .B2(new_n720), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  AOI211_X1 g302(.A(new_n709), .B(new_n727), .C1(G1341), .C2(new_n725), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n720), .A2(G26), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT28), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n489), .A2(G140), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n487), .A2(new_n488), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n732), .A2(G128), .A3(G2105), .ZN(new_n733));
  OAI21_X1  g308(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n734));
  INV_X1    g309(.A(G116), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(G2105), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n731), .A2(new_n733), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n730), .B1(new_n738), .B2(G29), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G2067), .ZN(new_n740));
  NAND2_X1  g315(.A1(G164), .A2(G29), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G27), .B2(G29), .ZN(new_n742));
  INV_X1    g317(.A(G2078), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT31), .B(G11), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT93), .ZN(new_n748));
  AND3_X1   g323(.A1(new_n748), .A2(new_n747), .A3(G28), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n747), .B2(G28), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n720), .B1(new_n747), .B2(G28), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n746), .B(new_n751), .C1(new_n711), .C2(G1966), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n744), .A2(new_n745), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g328(.A1(new_n728), .A2(new_n740), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n720), .A2(G33), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n489), .A2(G139), .ZN(new_n756));
  NAND2_X1  g331(.A1(G115), .A2(G2104), .ZN(new_n757));
  INV_X1    g332(.A(G127), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n485), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G2105), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT88), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT25), .Z(new_n764));
  NAND3_X1  g339(.A1(new_n759), .A2(KEYINPUT88), .A3(G2105), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n756), .A2(new_n762), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n755), .B1(new_n767), .B2(new_n720), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT89), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G2072), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT92), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n706), .A2(G20), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT23), .Z(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G299), .B2(G16), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT95), .B(G1956), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(G162), .A2(G29), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G29), .B2(G35), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT29), .B(G2090), .Z(new_n779));
  OAI21_X1  g354(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n778), .B2(new_n779), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n769), .A2(G2072), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n706), .A2(G4), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n614), .B2(new_n706), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1348), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n720), .A2(G32), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n489), .A2(G141), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n491), .A2(G129), .ZN(new_n788));
  NAND3_X1  g363(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT26), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n791), .A2(new_n792), .B1(G105), .B2(new_n479), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n787), .A2(new_n788), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n786), .B1(new_n795), .B2(new_n720), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT27), .B(G1996), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n721), .A2(new_n722), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT94), .ZN(new_n800));
  NOR4_X1   g375(.A1(new_n782), .A2(new_n785), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n754), .A2(new_n771), .A3(new_n781), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n706), .A2(G23), .ZN(new_n803));
  INV_X1    g378(.A(G288), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n706), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT33), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1976), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n706), .A2(G22), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G166), .B2(new_n706), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT87), .Z(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(G1971), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(G1971), .ZN(new_n812));
  NOR2_X1   g387(.A1(G6), .A2(G16), .ZN(new_n813));
  INV_X1    g388(.A(new_n597), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(new_n591), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n813), .B1(new_n815), .B2(G16), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT32), .B(G1981), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT86), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n816), .B(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n807), .A2(new_n811), .A3(new_n812), .A4(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT85), .B(KEYINPUT34), .Z(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n489), .A2(G131), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n491), .A2(G119), .ZN(new_n825));
  NOR2_X1   g400(.A1(G95), .A2(G2105), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT83), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT84), .ZN(new_n828));
  INV_X1    g403(.A(G107), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n478), .B1(new_n829), .B2(G2105), .ZN(new_n830));
  AND3_X1   g405(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n828), .B1(new_n827), .B2(new_n830), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n824), .B(new_n825), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G29), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(G25), .B2(G29), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT35), .B(G1991), .Z(new_n837));
  AND2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n706), .A2(G24), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n604), .B2(new_n706), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G1986), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n838), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n822), .A2(new_n823), .A3(new_n843), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(KEYINPUT36), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(KEYINPUT36), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n802), .B1(new_n845), .B2(new_n846), .ZN(G311));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  INV_X1    g423(.A(new_n802), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(G150));
  NAND3_X1  g425(.A1(new_n521), .A2(new_n525), .A3(G93), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n525), .A2(G55), .A3(G543), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n520), .ZN(new_n854));
  NOR2_X1   g429(.A1(KEYINPUT5), .A2(G543), .ZN(new_n855));
  OAI21_X1  g430(.A(G67), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n523), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(KEYINPUT97), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n853), .A2(new_n858), .A3(KEYINPUT97), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(G860), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n613), .A2(new_n612), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n608), .A2(new_n523), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n607), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(new_n627), .ZN(new_n869));
  XOR2_X1   g444(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  AOI22_X1  g446(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n872));
  OAI221_X1 g447(.A(new_n552), .B1(new_n526), .B2(new_n553), .C1(new_n872), .C2(new_n523), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n860), .B2(new_n861), .ZN(new_n874));
  INV_X1    g449(.A(new_n858), .ZN(new_n875));
  INV_X1    g450(.A(new_n853), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n558), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n871), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n880), .A2(KEYINPUT39), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n863), .B1(new_n880), .B2(KEYINPUT39), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n865), .B1(new_n881), .B2(new_n882), .ZN(G145));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n491), .A2(G130), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n491), .A2(KEYINPUT98), .A3(G130), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  INV_X1    g465(.A(G118), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n891), .B2(G2105), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n489), .A2(G142), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n889), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n833), .A2(new_n634), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n833), .A2(new_n634), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n895), .B1(new_n901), .B2(new_n897), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n738), .A2(new_n515), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n736), .B1(new_n491), .B2(G128), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n907), .A2(new_n731), .B1(new_n514), .B2(new_n505), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n767), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n738), .A2(new_n515), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n907), .A2(new_n514), .A3(new_n505), .A4(new_n731), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n911), .A3(new_n766), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(new_n795), .A3(new_n912), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n910), .A2(new_n911), .A3(new_n766), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n766), .B1(new_n910), .B2(new_n911), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n794), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n904), .A2(new_n905), .A3(new_n913), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n913), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT100), .B1(new_n918), .B2(new_n903), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n918), .A2(KEYINPUT99), .A3(new_n903), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT99), .B1(new_n918), .B2(new_n903), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n917), .B(new_n919), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n644), .B(new_n481), .ZN(new_n923));
  XNOR2_X1  g498(.A(G162), .B(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n918), .A2(new_n903), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n924), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n914), .A2(new_n915), .A3(new_n794), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n795), .B1(new_n909), .B2(new_n912), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT101), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n916), .A2(new_n933), .A3(new_n913), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n934), .A3(new_n904), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT102), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n932), .A2(new_n904), .A3(new_n937), .A4(new_n934), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n929), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n926), .B(new_n927), .C1(new_n939), .C2(KEYINPUT103), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n939), .A2(KEYINPUT103), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n884), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n939), .A2(KEYINPUT103), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n939), .A2(KEYINPUT103), .ZN(new_n944));
  AOI21_X1  g519(.A(G37), .B1(new_n922), .B2(new_n925), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n943), .A2(KEYINPUT40), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n942), .A2(new_n946), .ZN(G395));
  XNOR2_X1  g522(.A(new_n629), .B(KEYINPUT104), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(new_n878), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n624), .A2(new_n614), .ZN(new_n950));
  NAND2_X1  g525(.A1(G299), .A2(new_n868), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT41), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT41), .B1(new_n950), .B2(new_n951), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n953), .B1(new_n949), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(G290), .A2(new_n815), .ZN(new_n958));
  NAND2_X1  g533(.A1(G305), .A2(new_n604), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(G303), .A2(new_n804), .ZN(new_n961));
  NAND2_X1  g536(.A1(G166), .A2(G288), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n958), .A2(new_n961), .A3(new_n959), .A4(new_n962), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(KEYINPUT105), .B2(KEYINPUT42), .ZN(new_n967));
  NOR2_X1   g542(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n967), .B(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n957), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(G868), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(G868), .B2(new_n862), .ZN(G295));
  OAI21_X1  g547(.A(new_n971), .B1(G868), .B2(new_n862), .ZN(G331));
  OR2_X1    g548(.A1(new_n549), .A2(new_n523), .ZN(new_n974));
  AOI22_X1  g549(.A1(new_n567), .A2(new_n546), .B1(G52), .B2(new_n534), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n974), .B(new_n975), .C1(new_n539), .C2(new_n543), .ZN(new_n976));
  INV_X1    g551(.A(new_n543), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n977), .B(new_n538), .C1(new_n550), .C2(new_n548), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n874), .A2(new_n877), .A3(new_n976), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n978), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT97), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n876), .A2(new_n981), .A3(new_n875), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n558), .B1(new_n982), .B2(new_n859), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n873), .A2(new_n858), .A3(new_n853), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n952), .B1(new_n979), .B2(new_n985), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n980), .A2(new_n983), .A3(new_n984), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n874), .A2(new_n877), .B1(new_n976), .B2(new_n978), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n986), .B1(new_n956), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(G37), .B1(new_n990), .B2(new_n966), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT41), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n952), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT41), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n993), .A2(new_n994), .A3(new_n979), .A4(new_n985), .ZN(new_n995));
  INV_X1    g570(.A(new_n952), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n987), .B2(new_n988), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n966), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n991), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n995), .A2(new_n997), .A3(new_n966), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n927), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT106), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n990), .B2(new_n966), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n998), .A2(KEYINPUT106), .A3(new_n999), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT43), .ZN(new_n1008));
  MUX2_X1   g583(.A(new_n1001), .B(new_n1007), .S(new_n1008), .Z(new_n1009));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT107), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT106), .B1(new_n998), .B2(new_n999), .ZN(new_n1013));
  AOI211_X1 g588(.A(new_n1004), .B(new_n966), .C1(new_n995), .C2(new_n997), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n991), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n1016), .A3(KEYINPUT43), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n991), .A2(new_n1008), .A3(new_n1000), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT44), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT108), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT108), .ZN(new_n1023));
  AOI211_X1 g598(.A(new_n1023), .B(new_n1020), .C1(new_n1012), .C2(new_n1017), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1011), .B1(new_n1022), .B2(new_n1024), .ZN(G397));
  INV_X1    g600(.A(G1981), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n592), .B2(new_n597), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n597), .A2(new_n1026), .A3(new_n590), .A4(new_n589), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n815), .A2(new_n1029), .A3(new_n1026), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT49), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G8), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1384), .B1(new_n505), .B2(new_n514), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n474), .A2(G40), .A3(new_n480), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1038));
  OAI21_X1  g613(.A(G1981), .B1(new_n814), .B2(new_n591), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(new_n1029), .A3(new_n1028), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT49), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1033), .A2(new_n1037), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n804), .A2(G1976), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT52), .B1(G288), .B2(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1037), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1048), .B1(new_n1037), .B2(new_n1044), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1035), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT114), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n474), .A2(G40), .A3(new_n480), .ZN(new_n1054));
  INV_X1    g629(.A(G1384), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n511), .A2(new_n513), .ZN(new_n1056));
  INV_X1    g631(.A(new_n498), .ZN(new_n1057));
  INV_X1    g632(.A(new_n504), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n503), .B1(new_n475), .B2(new_n500), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1055), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1054), .B1(new_n1061), .B2(KEYINPUT50), .ZN(new_n1062));
  AOI211_X1 g637(.A(KEYINPUT50), .B(G1384), .C1(new_n505), .C2(new_n514), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G2090), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1053), .A2(new_n1062), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G1971), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT45), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(G1384), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n1036), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1035), .A2(KEYINPUT45), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1068), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1034), .B1(new_n1067), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(G303), .A2(G8), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1076), .B(new_n1077), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1043), .B(new_n1050), .C1(new_n1075), .C2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT111), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1036), .B1(new_n1035), .B2(new_n1051), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1081), .A2(G2090), .A3(new_n1063), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1061), .A2(new_n1069), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1054), .B1(new_n515), .B2(new_n1070), .ZN(new_n1084));
  AOI21_X1  g659(.A(G1971), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1080), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1061), .A2(KEYINPUT50), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1087), .A2(new_n1066), .A3(new_n1036), .A4(new_n1052), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1074), .A2(new_n1088), .A3(KEYINPUT111), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1086), .A2(G8), .A3(new_n1089), .A4(new_n1078), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT112), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1074), .A2(new_n1088), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1034), .B1(new_n1093), .B2(new_n1080), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1094), .A2(KEYINPUT112), .A3(new_n1078), .A4(new_n1089), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1079), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1071), .B(new_n1036), .C1(KEYINPUT45), .C2(new_n1035), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(G2078), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT53), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1097), .B(new_n1101), .C1(new_n1098), .C2(G2078), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1961), .B1(new_n1062), .B2(new_n1052), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1100), .A2(G301), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT124), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1100), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(G171), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1103), .B1(new_n1099), .B2(KEYINPUT53), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1109), .A2(new_n1110), .A3(G301), .A4(new_n1102), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1106), .A2(new_n1108), .A3(KEYINPUT54), .A4(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G1966), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1098), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1087), .A2(new_n722), .A3(new_n1036), .A4(new_n1052), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(new_n1115), .A3(G168), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT51), .ZN(new_n1118));
  AOI21_X1  g693(.A(G168), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1120), .A2(KEYINPUT51), .ZN(new_n1121));
  OAI211_X1 g696(.A(G8), .B(new_n1116), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1105), .ZN(new_n1125));
  AOI21_X1  g700(.A(G301), .B1(new_n1109), .B2(new_n1102), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1124), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AND4_X1   g702(.A1(new_n1096), .A2(new_n1112), .A3(new_n1123), .A4(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1129), .A2(G2067), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1062), .A2(new_n1052), .ZN(new_n1131));
  INV_X1    g706(.A(G1348), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OR3_X1    g708(.A1(new_n1133), .A2(KEYINPUT118), .A3(new_n868), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n624), .A2(KEYINPUT57), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n621), .A2(KEYINPUT116), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n621), .A2(KEYINPUT116), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n620), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1135), .B1(new_n1138), .B2(KEYINPUT57), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1064), .B1(new_n1035), .B2(new_n1051), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1081), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(G1956), .B1(new_n1142), .B2(new_n1065), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT56), .B(G2072), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1140), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT118), .B1(new_n1133), .B2(new_n868), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1134), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1053), .A2(new_n1062), .A3(new_n1065), .ZN(new_n1150));
  INV_X1    g725(.A(G1956), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(new_n1139), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1152), .A2(KEYINPUT117), .A3(new_n1139), .A4(new_n1153), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1149), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT61), .B1(new_n1158), .B2(new_n1147), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1147), .A2(KEYINPUT61), .A3(new_n1154), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1132), .B1(new_n1081), .B2(new_n1063), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n614), .A2(KEYINPUT60), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1162), .B(new_n1163), .C1(G2067), .C2(new_n1129), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n614), .A2(KEYINPUT60), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT120), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1164), .B(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(KEYINPUT58), .B(G1341), .Z(new_n1168));
  NAND2_X1  g743(.A1(new_n1129), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(new_n1098), .B2(G1996), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT119), .B1(new_n1170), .B2(new_n558), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1170), .A2(KEYINPUT119), .A3(new_n558), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1171), .B1(KEYINPUT59), .B2(new_n1172), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1171), .A2(KEYINPUT59), .A3(new_n1172), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1161), .B(new_n1167), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1159), .B1(new_n1160), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1128), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1079), .ZN(new_n1179));
  NAND2_X1  g754(.A1(G168), .A2(G8), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1180), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1178), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1043), .A2(new_n1181), .A3(new_n1050), .A4(KEYINPUT63), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1078), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1086), .A2(G8), .A3(new_n1089), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1178), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(KEYINPUT115), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT115), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1178), .A2(new_n1188), .A3(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1184), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1043), .A2(new_n1045), .A3(new_n804), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1028), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1037), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1043), .A2(new_n1050), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1196), .B1(new_n1178), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1118), .A2(new_n1199), .A3(new_n1122), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(new_n1126), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1199), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1198), .B1(new_n1203), .B2(new_n1096), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1177), .A2(new_n1193), .A3(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT110), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT109), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1207), .B1(new_n1083), .B2(new_n1054), .ZN(new_n1208));
  NOR4_X1   g783(.A1(new_n1035), .A2(new_n1207), .A3(new_n1054), .A4(KEYINPUT45), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1206), .B1(new_n1211), .B2(G1996), .ZN(new_n1212));
  AOI21_X1  g787(.A(KEYINPUT109), .B1(new_n1073), .B2(new_n1036), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1213), .A2(new_n1209), .ZN(new_n1214));
  INV_X1    g789(.A(G1996), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1214), .A2(KEYINPUT110), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n794), .B1(new_n1212), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1217), .ZN(new_n1218));
  INV_X1    g793(.A(G2067), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n738), .B(new_n1219), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1220), .B1(new_n1215), .B2(new_n795), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1221), .A2(new_n1214), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n833), .B(new_n837), .ZN(new_n1223));
  OR2_X1    g798(.A1(new_n1211), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1218), .A2(new_n1222), .A3(new_n1224), .ZN(new_n1225));
  XOR2_X1   g800(.A(new_n604), .B(G1986), .Z(new_n1226));
  AOI21_X1  g801(.A(new_n1225), .B1(new_n1214), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1205), .A2(new_n1227), .ZN(new_n1228));
  NOR3_X1   g803(.A1(new_n1211), .A2(G1986), .A3(G290), .ZN(new_n1229));
  XNOR2_X1  g804(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1230));
  XNOR2_X1  g805(.A(new_n1229), .B(new_n1230), .ZN(new_n1231));
  NAND4_X1  g806(.A1(new_n1231), .A2(new_n1218), .A3(new_n1222), .A4(new_n1224), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1220), .A2(new_n795), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1233), .A2(new_n1214), .ZN(new_n1234));
  INV_X1    g809(.A(new_n1234), .ZN(new_n1235));
  INV_X1    g810(.A(KEYINPUT46), .ZN(new_n1236));
  NOR3_X1   g811(.A1(new_n1211), .A2(new_n1206), .A3(G1996), .ZN(new_n1237));
  AOI21_X1  g812(.A(KEYINPUT110), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1238));
  OAI21_X1  g813(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g814(.A1(new_n1212), .A2(KEYINPUT46), .A3(new_n1216), .ZN(new_n1240));
  AOI21_X1  g815(.A(new_n1235), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g816(.A(KEYINPUT47), .ZN(new_n1242));
  NOR2_X1   g817(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  AOI211_X1 g818(.A(KEYINPUT47), .B(new_n1235), .C1(new_n1239), .C2(new_n1240), .ZN(new_n1244));
  OAI21_X1  g819(.A(new_n1232), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g820(.A(new_n1222), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n834), .A2(new_n837), .ZN(new_n1247));
  XNOR2_X1  g822(.A(new_n1247), .B(KEYINPUT125), .ZN(new_n1248));
  NOR3_X1   g823(.A1(new_n1217), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1249));
  NAND3_X1  g824(.A1(new_n907), .A2(new_n1219), .A3(new_n731), .ZN(new_n1250));
  INV_X1    g825(.A(new_n1250), .ZN(new_n1251));
  OAI21_X1  g826(.A(new_n1214), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g827(.A(new_n1252), .ZN(new_n1253));
  OAI21_X1  g828(.A(KEYINPUT127), .B1(new_n1245), .B2(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g829(.A(new_n1241), .B(new_n1242), .ZN(new_n1255));
  INV_X1    g830(.A(KEYINPUT127), .ZN(new_n1256));
  NAND4_X1  g831(.A1(new_n1255), .A2(new_n1256), .A3(new_n1252), .A4(new_n1232), .ZN(new_n1257));
  NAND2_X1  g832(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g833(.A1(new_n1228), .A2(new_n1258), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g834(.A1(G227), .A2(new_n465), .ZN(new_n1261));
  NOR3_X1   g835(.A1(G229), .A2(G401), .A3(new_n1261), .ZN(new_n1262));
  OAI211_X1 g836(.A(new_n1262), .B(new_n1009), .C1(new_n940), .C2(new_n941), .ZN(G225));
  INV_X1    g837(.A(G225), .ZN(G308));
endmodule


