//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024;
  INV_X1    g000(.A(KEYINPUT16), .ZN(new_n202));
  AND2_X1   g001(.A1(G15gat), .A2(G22gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G15gat), .A2(G22gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G1gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT86), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n210), .B(new_n208), .C1(new_n203), .C2(new_n204), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n207), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n210), .B1(new_n203), .B2(new_n204), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G8gat), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n216), .A2(new_n206), .A3(new_n205), .A4(new_n212), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G71gat), .A2(G78gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT93), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT9), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G57gat), .B(G64gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n220), .B1(new_n219), .B2(new_n221), .ZN(new_n225));
  NOR3_X1   g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G71gat), .ZN(new_n227));
  INV_X1    g026(.A(G78gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(new_n219), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(new_n224), .B2(KEYINPUT94), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G64gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G57gat), .ZN(new_n234));
  INV_X1    g033(.A(G57gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G64gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT94), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n237), .A2(new_n238), .B1(new_n219), .B2(new_n229), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n221), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT93), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(new_n237), .A3(new_n222), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n232), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n218), .B1(KEYINPUT21), .B2(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(G127gat), .B(G155gat), .Z(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n244), .A2(KEYINPUT21), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n248), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n252), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n249), .A2(new_n254), .A3(new_n250), .ZN(new_n255));
  XOR2_X1   g054(.A(G183gat), .B(G211gat), .Z(new_n256));
  NAND2_X1  g055(.A1(G231gat), .A2(G233gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT95), .B(KEYINPUT96), .Z(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n253), .A2(new_n255), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n260), .B1(new_n253), .B2(new_n255), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(G232gat), .A2(G233gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(KEYINPUT41), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(G162gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(G99gat), .A2(G106gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(G99gat), .A2(G106gat), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT97), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G99gat), .ZN(new_n271));
  INV_X1    g070(.A(G106gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT97), .ZN(new_n274));
  NAND2_X1  g073(.A1(G99gat), .A2(G106gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G85gat), .A2(G92gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT7), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT7), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n280), .A2(G85gat), .A3(G92gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G85gat), .ZN(new_n283));
  INV_X1    g082(.A(G92gat), .ZN(new_n284));
  AOI22_X1  g083(.A1(KEYINPUT8), .A2(new_n275), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n277), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n270), .A2(new_n276), .A3(new_n282), .A4(new_n285), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G29gat), .A2(G36gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT14), .ZN(new_n292));
  INV_X1    g091(.A(G29gat), .ZN(new_n293));
  INV_X1    g092(.A(G36gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n294), .A3(KEYINPUT14), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G50gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G43gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT15), .ZN(new_n301));
  INV_X1    g100(.A(G43gat), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n301), .B1(new_n302), .B2(G50gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n298), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT17), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT85), .B1(new_n299), .B2(G43gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT85), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(new_n302), .A3(G50gat), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n302), .A2(KEYINPUT84), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT84), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G43gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n312), .A3(new_n299), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT15), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n302), .A2(G50gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n300), .A2(new_n315), .A3(KEYINPUT15), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(new_n296), .A3(new_n297), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n304), .B(new_n305), .C1(new_n314), .C2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n310), .A2(new_n312), .A3(new_n299), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n306), .A2(new_n308), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n301), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n316), .A2(new_n296), .A3(new_n297), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n305), .B1(new_n324), .B2(new_n304), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n290), .B1(new_n319), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n316), .B1(new_n297), .B2(new_n296), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n327), .B1(new_n322), .B2(new_n323), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n290), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n264), .A2(KEYINPUT41), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n326), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT98), .B(G134gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n326), .A2(new_n330), .A3(new_n331), .A4(new_n333), .ZN(new_n336));
  XNOR2_X1  g135(.A(G190gat), .B(G218gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n338), .B1(new_n335), .B2(new_n336), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n267), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n335), .A2(new_n336), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n337), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n266), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G230gat), .A2(G233gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n226), .A2(new_n231), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n239), .A2(new_n242), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n289), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT99), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n232), .A2(new_n243), .A3(new_n288), .A4(new_n287), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n290), .A2(KEYINPUT99), .A3(new_n232), .A4(new_n243), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT10), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n347), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT100), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g159(.A(KEYINPUT100), .B(new_n347), .C1(new_n355), .C2(new_n357), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G120gat), .B(G148gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT101), .ZN(new_n364));
  INV_X1    g163(.A(G176gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n366), .B(G204gat), .Z(new_n367));
  NAND2_X1  g166(.A1(new_n353), .A2(new_n354), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n362), .B(new_n367), .C1(new_n347), .C2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n367), .ZN(new_n370));
  INV_X1    g169(.A(new_n358), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n368), .A2(new_n347), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n263), .A2(new_n346), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G15gat), .B(G43gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT68), .ZN(new_n378));
  OR2_X1    g177(.A1(new_n378), .A2(new_n227), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n227), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n379), .A2(new_n380), .A3(G99gat), .ZN(new_n381));
  AOI21_X1  g180(.A(G99gat), .B1(new_n379), .B2(new_n380), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT26), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n387));
  INV_X1    g186(.A(G169gat), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n386), .B(new_n387), .C1(new_n388), .C2(new_n365), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT27), .B(G183gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT28), .ZN(new_n391));
  INV_X1    g190(.A(G190gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G183gat), .A2(G190gat), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n389), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  XOR2_X1   g194(.A(KEYINPUT27), .B(G183gat), .Z(new_n396));
  INV_X1    g195(.A(KEYINPUT65), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n390), .A2(KEYINPUT65), .ZN(new_n399));
  AOI21_X1  g198(.A(G190gat), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n395), .B1(new_n400), .B2(new_n391), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT23), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n384), .B(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n394), .A2(KEYINPUT24), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n365), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OR2_X1    g205(.A1(G183gat), .A2(G190gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT24), .A3(new_n394), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n403), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT25), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n403), .A2(new_n406), .A3(KEYINPUT25), .A4(new_n408), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n401), .A2(new_n413), .ZN(new_n414));
  XOR2_X1   g213(.A(G127gat), .B(G134gat), .Z(new_n415));
  XNOR2_X1  g214(.A(G113gat), .B(G120gat), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n416), .A2(KEYINPUT66), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT1), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(new_n416), .B2(KEYINPUT66), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n415), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT67), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT1), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n415), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n422), .B(new_n423), .C1(new_n421), .C2(new_n416), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n414), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(G227gat), .A2(G233gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT64), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n420), .A2(new_n424), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n401), .A2(new_n413), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n426), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT32), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT33), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n383), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT33), .B1(new_n381), .B2(new_n382), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n432), .A2(new_n436), .A3(KEYINPUT32), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT69), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n432), .A2(new_n436), .A3(KEYINPUT69), .A4(KEYINPUT32), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n431), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n427), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT34), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT34), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n442), .A2(new_n445), .A3(new_n428), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT70), .B1(new_n441), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n441), .A2(new_n448), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT36), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n439), .A2(new_n440), .ZN(new_n453));
  INV_X1    g252(.A(new_n435), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(new_n447), .ZN(new_n456));
  OR3_X1    g255(.A1(new_n456), .A2(KEYINPUT36), .A3(new_n450), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G22gat), .B(G50gat), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(G228gat), .A2(G233gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(G197gat), .B(G204gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT22), .ZN(new_n463));
  NAND2_X1  g262(.A1(G211gat), .A2(G218gat), .ZN(new_n464));
  INV_X1    g263(.A(G211gat), .ZN(new_n465));
  INV_X1    g264(.A(G218gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT71), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT22), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n464), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n462), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT71), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n463), .A2(new_n473), .A3(new_n464), .A4(new_n467), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT29), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT2), .ZN(new_n480));
  INV_X1    g279(.A(G148gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(G141gat), .ZN(new_n482));
  INV_X1    g281(.A(G141gat), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(G148gat), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n480), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G155gat), .A2(G162gat), .ZN(new_n486));
  INV_X1    g285(.A(G155gat), .ZN(new_n487));
  INV_X1    g286(.A(G162gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n486), .B1(new_n489), .B2(KEYINPUT2), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT76), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n492), .B1(new_n483), .B2(G148gat), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n481), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n491), .B1(new_n495), .B2(new_n482), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n479), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n478), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n476), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT72), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n475), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n469), .A2(KEYINPUT72), .A3(new_n472), .A4(new_n474), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n501), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n461), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n468), .A2(new_n472), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n478), .B1(new_n507), .B2(KEYINPUT29), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n508), .A2(new_n498), .B1(G228gat), .B2(G233gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT31), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT31), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n501), .A2(new_n503), .A3(new_n504), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n497), .B1(new_n477), .B2(new_n478), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n513), .B(new_n510), .C1(new_n516), .C2(new_n461), .ZN(new_n517));
  XOR2_X1   g316(.A(G78gat), .B(G106gat), .Z(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n512), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n512), .B2(new_n517), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n460), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n512), .A2(new_n517), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n518), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n512), .A2(new_n517), .A3(new_n519), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n459), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G8gat), .B(G36gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT75), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(G64gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(new_n284), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT74), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n401), .A2(new_n413), .ZN(new_n535));
  NAND2_X1  g334(.A1(G226gat), .A2(G233gat), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n536), .B(KEYINPUT73), .Z(new_n537));
  OAI21_X1  g336(.A(new_n534), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n536), .B1(new_n535), .B2(KEYINPUT29), .ZN(new_n539));
  INV_X1    g338(.A(new_n537), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n414), .A2(KEYINPUT74), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n503), .A2(new_n504), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n535), .A2(new_n536), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n540), .B1(new_n414), .B2(new_n476), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(new_n543), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n533), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n547), .A2(new_n543), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n542), .A2(new_n543), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n551), .A3(new_n532), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n549), .A2(new_n552), .A3(KEYINPUT30), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n551), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n555), .A3(new_n533), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G225gat), .A2(G233gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n425), .A2(new_n497), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n559), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n498), .A2(KEYINPUT3), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n430), .A2(KEYINPUT77), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT77), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n566), .B1(new_n420), .B2(new_n424), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n500), .B(new_n564), .C1(new_n565), .C2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT4), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n563), .B(new_n568), .C1(new_n569), .C2(new_n560), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n498), .A2(new_n430), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n430), .B(KEYINPUT77), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(new_n498), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n570), .B(new_n571), .C1(new_n558), .C2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n571), .A2(new_n559), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n569), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n561), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n568), .A2(new_n576), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT80), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n575), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G1gat), .B(G29gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT0), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G57gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(new_n283), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n568), .A2(new_n577), .A3(new_n578), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n559), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n558), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(new_n593), .A3(KEYINPUT39), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n594), .B(new_n587), .C1(KEYINPUT39), .C2(new_n592), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT40), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n557), .A2(new_n590), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n596), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n528), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT6), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n575), .B(new_n587), .C1(new_n581), .C2(new_n582), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n589), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n532), .B1(new_n550), .B2(new_n551), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n605));
  OAI211_X1 g404(.A(KEYINPUT37), .B(new_n605), .C1(new_n542), .C2(new_n543), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT38), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n606), .A2(new_n607), .A3(new_n532), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT81), .B(KEYINPUT37), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n544), .B2(new_n548), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n604), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n583), .A2(KEYINPUT6), .A3(new_n588), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n603), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT82), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n611), .B1(new_n554), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT38), .B1(new_n617), .B2(new_n533), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT82), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n603), .A2(new_n612), .A3(new_n619), .A4(new_n613), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n615), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n458), .B1(new_n600), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n603), .A2(new_n613), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n557), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n528), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n455), .A2(new_n447), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n449), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n455), .A2(KEYINPUT70), .A3(new_n447), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT83), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n630), .A2(new_n527), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(new_n630), .B2(new_n527), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n623), .A2(KEYINPUT35), .A3(new_n557), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT35), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n456), .A2(new_n450), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n527), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n636), .B1(new_n624), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n214), .A2(new_n217), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT87), .B1(new_n643), .B2(new_n328), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n304), .B1(new_n314), .B2(new_n317), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT87), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n645), .A2(new_n646), .A3(new_n217), .A4(new_n214), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n648), .B1(new_n218), .B2(new_n645), .ZN(new_n649));
  NAND2_X1  g448(.A1(G229gat), .A2(G233gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n650), .B(KEYINPUT13), .Z(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n643), .B1(new_n319), .B2(new_n325), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT88), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n648), .A2(new_n653), .A3(new_n654), .A4(new_n650), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT18), .B1(new_n655), .B2(KEYINPUT89), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT88), .B1(KEYINPUT89), .B2(KEYINPUT18), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n645), .A2(KEYINPUT17), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n318), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n659), .A2(new_n643), .B1(new_n644), .B2(new_n647), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n657), .B1(new_n660), .B2(new_n650), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n652), .B1(new_n656), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G113gat), .B(G141gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G197gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT11), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n665), .A2(G169gat), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(G169gat), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(KEYINPUT12), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n665), .B(G169gat), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT12), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n662), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n668), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n652), .B(new_n673), .C1(new_n656), .C2(new_n661), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT90), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT91), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n656), .A2(new_n661), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n681), .A2(KEYINPUT90), .A3(new_n652), .A4(new_n673), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n674), .A2(new_n675), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(KEYINPUT91), .A3(new_n672), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n642), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT92), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n642), .A2(KEYINPUT92), .A3(new_n687), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n376), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n623), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G1gat), .ZN(G1324gat));
  INV_X1    g494(.A(new_n557), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n202), .A2(new_n208), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n208), .B1(new_n692), .B2(new_n696), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT42), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(KEYINPUT42), .B2(new_n700), .ZN(G1325gat));
  AOI21_X1  g502(.A(G15gat), .B1(new_n692), .B2(new_n637), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n458), .A2(G15gat), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n692), .B2(new_n705), .ZN(G1326gat));
  NAND2_X1  g505(.A1(new_n692), .A2(new_n528), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT43), .B(G22gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1327gat));
  INV_X1    g508(.A(new_n263), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n374), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT92), .B1(new_n642), .B2(new_n687), .ZN(new_n712));
  AOI211_X1 g511(.A(new_n689), .B(new_n686), .C1(new_n626), .C2(new_n641), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n346), .B(new_n711), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n293), .A3(new_n693), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT45), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  INV_X1    g517(.A(new_n346), .ZN(new_n719));
  AOI211_X1 g518(.A(new_n718), .B(new_n719), .C1(new_n626), .C2(new_n641), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n635), .B2(new_n640), .ZN(new_n722));
  INV_X1    g521(.A(new_n633), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n630), .A2(new_n527), .A3(new_n631), .ZN(new_n724));
  INV_X1    g523(.A(new_n634), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(KEYINPUT104), .A3(new_n639), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n621), .A2(new_n600), .ZN(new_n729));
  INV_X1    g528(.A(new_n458), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT102), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n624), .A2(new_n731), .A3(new_n528), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n603), .A2(new_n613), .B1(new_n556), .B2(new_n553), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT102), .B1(new_n733), .B2(new_n527), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n729), .A2(new_n730), .A3(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n622), .A2(KEYINPUT103), .A3(new_n735), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n728), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n346), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n720), .B1(new_n741), .B2(new_n718), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n711), .A2(new_n678), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G29gat), .B1(new_n745), .B2(new_n623), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n717), .A2(new_n746), .ZN(G1328gat));
  NAND3_X1  g546(.A1(new_n715), .A2(new_n294), .A3(new_n696), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n748), .A2(KEYINPUT46), .ZN(new_n749));
  OAI21_X1  g548(.A(G36gat), .B1(new_n745), .B2(new_n557), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(KEYINPUT46), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(G1329gat));
  NAND2_X1  g551(.A1(new_n310), .A2(new_n312), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n715), .A2(new_n637), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT44), .B1(new_n740), .B2(new_n346), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n755), .A2(new_n730), .A3(new_n743), .A4(new_n720), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT47), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT105), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n756), .B2(new_n753), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  OAI221_X1 g560(.A(new_n754), .B1(new_n759), .B2(KEYINPUT47), .C1(new_n753), .C2(new_n756), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1330gat));
  OAI21_X1  g562(.A(new_n299), .B1(new_n714), .B2(new_n527), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT48), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n528), .A2(G50gat), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n764), .B(new_n766), .C1(new_n745), .C2(new_n767), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n765), .A2(KEYINPUT48), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1331gat));
  INV_X1    g569(.A(new_n678), .ZN(new_n771));
  INV_X1    g570(.A(new_n374), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n263), .A2(new_n346), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n740), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n623), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(new_n235), .ZN(G1332gat));
  NOR2_X1   g575(.A1(new_n774), .A2(new_n557), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  AND2_X1   g577(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n777), .B2(new_n778), .ZN(G1333gat));
  INV_X1    g580(.A(new_n637), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n227), .B1(new_n774), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n458), .A2(G71gat), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n774), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g585(.A1(new_n774), .A2(new_n527), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(new_n228), .ZN(G1335gat));
  NAND2_X1  g587(.A1(new_n263), .A2(new_n771), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT107), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n742), .A2(new_n374), .A3(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n792), .A2(new_n283), .A3(new_n623), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n740), .A2(new_n346), .A3(new_n791), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n795), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n799), .A2(new_n693), .A3(new_n374), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n793), .B1(new_n800), .B2(new_n283), .ZN(G1336gat));
  NAND3_X1  g600(.A1(new_n696), .A2(new_n284), .A3(new_n374), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT109), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n794), .A2(new_n795), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n796), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT108), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR4_X1   g607(.A1(new_n755), .A2(new_n772), .A3(new_n720), .A4(new_n790), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n284), .B1(new_n809), .B2(new_n696), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n803), .B1(new_n797), .B2(new_n798), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n808), .B(KEYINPUT52), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G92gat), .B1(new_n792), .B2(new_n557), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n813), .B(new_n806), .C1(new_n807), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n815), .ZN(G1337gat));
  XOR2_X1   g615(.A(KEYINPUT110), .B(G99gat), .Z(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n792), .B2(new_n730), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n799), .A2(new_n374), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n782), .A2(new_n817), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(G1338gat));
  NAND4_X1  g620(.A1(new_n742), .A2(new_n528), .A3(new_n374), .A4(new_n791), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G106gat), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n527), .A2(G106gat), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n374), .B(new_n824), .C1(new_n805), .C2(new_n796), .ZN(new_n825));
  XNOR2_X1  g624(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n823), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n826), .B1(new_n823), .B2(new_n825), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(G1339gat));
  NOR2_X1   g628(.A1(new_n376), .A2(new_n678), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n832));
  AOI211_X1 g631(.A(new_n372), .B(new_n370), .C1(new_n360), .C2(new_n361), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n368), .A2(new_n356), .ZN(new_n834));
  INV_X1    g633(.A(new_n347), .ZN(new_n835));
  INV_X1    g634(.A(new_n357), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(KEYINPUT54), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n362), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n840), .B(new_n347), .C1(new_n355), .C2(new_n357), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n370), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n833), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n837), .A2(KEYINPUT54), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n847), .B1(new_n360), .B2(new_n361), .ZN(new_n848));
  NOR4_X1   g647(.A1(new_n848), .A2(KEYINPUT112), .A3(new_n845), .A4(new_n842), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT112), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n842), .B1(new_n362), .B2(new_n838), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n851), .B2(KEYINPUT55), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n846), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n649), .A2(new_n651), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n660), .A2(new_n650), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n669), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n684), .A2(new_n346), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n832), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n369), .B1(new_n851), .B2(KEYINPUT55), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n839), .A2(KEYINPUT55), .A3(new_n843), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT112), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n851), .A2(new_n850), .A3(KEYINPUT55), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n860), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI221_X4 g663(.A(new_n856), .B1(new_n341), .B2(new_n345), .C1(new_n682), .C2(new_n683), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT113), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n859), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n678), .B(new_n846), .C1(new_n852), .C2(new_n849), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n684), .A2(new_n374), .A3(new_n857), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n719), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n867), .A2(new_n871), .A3(KEYINPUT114), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n263), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT114), .B1(new_n867), .B2(new_n871), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n831), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n638), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n696), .A2(new_n623), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G113gat), .B1(new_n878), .B2(new_n686), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n877), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n723), .A2(new_n724), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n771), .A2(G113gat), .ZN(new_n883));
  XOR2_X1   g682(.A(new_n883), .B(KEYINPUT115), .Z(new_n884));
  OAI21_X1  g683(.A(new_n879), .B1(new_n882), .B2(new_n884), .ZN(G1340gat));
  OAI21_X1  g684(.A(G120gat), .B1(new_n878), .B2(new_n772), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n772), .A2(G120gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n882), .B2(new_n887), .ZN(G1341gat));
  INV_X1    g687(.A(new_n878), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(G127gat), .A3(new_n710), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(G127gat), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n893), .B1(new_n882), .B2(new_n263), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n889), .A2(KEYINPUT116), .A3(G127gat), .A4(new_n710), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT117), .ZN(G1342gat));
  NOR2_X1   g696(.A1(new_n880), .A2(new_n881), .ZN(new_n898));
  INV_X1    g697(.A(G134gat), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n899), .A3(new_n346), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT56), .ZN(new_n901));
  OAI21_X1  g700(.A(G134gat), .B1(new_n878), .B2(new_n719), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT56), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n898), .A2(new_n903), .A3(new_n899), .A4(new_n346), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n905), .B(new_n906), .ZN(G1343gat));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n875), .A2(new_n910), .A3(new_n528), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n730), .A2(new_n877), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n853), .A2(new_n832), .A3(new_n858), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT113), .B1(new_n864), .B2(new_n865), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n864), .A2(new_n680), .A3(new_n685), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n346), .B1(new_n917), .B2(new_n869), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n263), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT119), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n830), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g720(.A(KEYINPUT119), .B(new_n263), .C1(new_n916), .C2(new_n918), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n527), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n911), .B(new_n913), .C1(new_n923), .C2(new_n910), .ZN(new_n924));
  OAI21_X1  g723(.A(G141gat), .B1(new_n924), .B2(new_n771), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n458), .A2(new_n527), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT120), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n875), .A2(new_n687), .A3(new_n877), .A4(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n928), .A2(G141gat), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n909), .B1(new_n925), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n909), .B1(new_n928), .B2(G141gat), .ZN(new_n932));
  INV_X1    g731(.A(new_n874), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n263), .A3(new_n872), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n527), .B1(new_n934), .B2(new_n831), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n912), .B1(new_n935), .B2(new_n910), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n922), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n528), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT57), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n936), .A2(new_n939), .A3(new_n687), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n932), .B1(new_n940), .B2(G141gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n908), .B1(new_n931), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(G141gat), .B1(new_n924), .B2(new_n686), .ZN(new_n943));
  INV_X1    g742(.A(new_n932), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n936), .A2(new_n939), .A3(new_n678), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n929), .B1(new_n946), .B2(G141gat), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n945), .B(KEYINPUT121), .C1(new_n947), .C2(new_n909), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n942), .A2(new_n948), .ZN(G1344gat));
  NAND2_X1  g748(.A1(new_n875), .A2(new_n528), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT57), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n375), .A2(new_n686), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT122), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n918), .B1(new_n864), .B2(new_n865), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n954), .A2(new_n710), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n910), .B(new_n528), .C1(new_n953), .C2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n951), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n913), .A2(new_n374), .ZN(new_n958));
  OAI211_X1 g757(.A(KEYINPUT59), .B(G148gat), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n875), .A2(new_n877), .A3(new_n927), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(new_n481), .A3(new_n374), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n936), .A2(new_n939), .A3(new_n374), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT59), .B1(new_n963), .B2(G148gat), .ZN(new_n964));
  OAI21_X1  g763(.A(KEYINPUT123), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(G148gat), .B1(new_n924), .B2(new_n772), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT59), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n968), .A2(new_n969), .A3(new_n959), .A4(new_n961), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n965), .A2(new_n970), .ZN(G1345gat));
  NOR3_X1   g770(.A1(new_n924), .A2(new_n487), .A3(new_n263), .ZN(new_n972));
  AOI21_X1  g771(.A(G155gat), .B1(new_n960), .B2(new_n710), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n972), .A2(new_n973), .ZN(G1346gat));
  OAI21_X1  g773(.A(G162gat), .B1(new_n924), .B2(new_n719), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n960), .A2(new_n488), .A3(new_n346), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1347gat));
  NOR2_X1   g776(.A1(new_n693), .A2(new_n557), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n875), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(new_n876), .ZN(new_n980));
  OAI21_X1  g779(.A(G169gat), .B1(new_n980), .B2(new_n686), .ZN(new_n981));
  AND4_X1   g780(.A1(new_n723), .A2(new_n875), .A3(new_n724), .A4(new_n978), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n982), .A2(new_n388), .A3(new_n678), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n981), .A2(new_n983), .ZN(G1348gat));
  OAI21_X1  g783(.A(G176gat), .B1(new_n980), .B2(new_n772), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n982), .A2(new_n365), .A3(new_n374), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g786(.A(new_n987), .B(KEYINPUT124), .Z(G1349gat));
  OAI21_X1  g787(.A(G183gat), .B1(new_n980), .B2(new_n263), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n263), .B1(new_n399), .B2(new_n398), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n982), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g792(.A1(new_n982), .A2(new_n392), .A3(new_n346), .ZN(new_n994));
  OAI21_X1  g793(.A(G190gat), .B1(new_n980), .B2(new_n719), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n995), .A2(KEYINPUT61), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n995), .A2(KEYINPUT61), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(G1351gat));
  AND2_X1   g797(.A1(new_n951), .A2(new_n956), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n730), .A2(new_n978), .ZN(new_n1000));
  XOR2_X1   g799(.A(new_n1000), .B(KEYINPUT125), .Z(new_n1001));
  NAND2_X1  g800(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g801(.A(G197gat), .B1(new_n1002), .B2(new_n686), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n979), .A2(new_n926), .ZN(new_n1004));
  OR2_X1    g803(.A1(new_n771), .A2(G197gat), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(G1352gat));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1007), .B1(new_n1002), .B2(new_n772), .ZN(new_n1008));
  NAND4_X1  g807(.A1(new_n999), .A2(KEYINPUT126), .A3(new_n374), .A4(new_n1001), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n1008), .A2(G204gat), .A3(new_n1009), .ZN(new_n1010));
  NOR3_X1   g809(.A1(new_n1004), .A2(G204gat), .A3(new_n772), .ZN(new_n1011));
  XNOR2_X1  g810(.A(new_n1011), .B(KEYINPUT62), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1010), .A2(new_n1012), .ZN(G1353gat));
  NAND4_X1  g812(.A1(new_n979), .A2(new_n465), .A3(new_n710), .A4(new_n926), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n999), .A2(new_n710), .A3(new_n1001), .ZN(new_n1015));
  AND3_X1   g814(.A1(new_n1015), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1016));
  AOI21_X1  g815(.A(KEYINPUT63), .B1(new_n1015), .B2(G211gat), .ZN(new_n1017));
  OAI21_X1  g816(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(G1354gat));
  OAI21_X1  g817(.A(new_n466), .B1(new_n1004), .B2(new_n719), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n346), .A2(G218gat), .ZN(new_n1020));
  OAI21_X1  g819(.A(new_n1019), .B1(new_n1002), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1021), .A2(KEYINPUT127), .ZN(new_n1022));
  INV_X1    g821(.A(KEYINPUT127), .ZN(new_n1023));
  OAI211_X1 g822(.A(new_n1023), .B(new_n1019), .C1(new_n1002), .C2(new_n1020), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1022), .A2(new_n1024), .ZN(G1355gat));
endmodule


