//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G128), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT24), .B(G110), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT76), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT74), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n190), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n190), .A2(new_n196), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n189), .A2(KEYINPUT74), .A3(KEYINPUT23), .A4(G119), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n197), .A2(new_n188), .A3(new_n198), .A4(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n194), .B1(G110), .B2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G125), .B(G140), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NOR3_X1   g019(.A1(new_n205), .A2(KEYINPUT16), .A3(G140), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n206), .B1(new_n202), .B2(KEYINPUT16), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n201), .A2(new_n204), .A3(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n191), .A2(new_n192), .ZN(new_n210));
  OR2_X1    g024(.A1(new_n207), .A2(G146), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(new_n208), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n200), .B(KEYINPUT75), .ZN(new_n213));
  INV_X1    g027(.A(G110), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT69), .B(G953), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(G221), .A3(G234), .ZN(new_n218));
  XOR2_X1   g032(.A(new_n218), .B(KEYINPUT22), .Z(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(G137), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G137), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n219), .B(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n209), .A3(new_n215), .ZN(new_n224));
  INV_X1    g038(.A(G902), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT77), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT25), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT25), .B1(new_n226), .B2(new_n227), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G217), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(G234), .B2(new_n225), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(G902), .ZN(new_n233));
  XOR2_X1   g047(.A(new_n233), .B(KEYINPUT78), .Z(new_n234));
  NAND2_X1  g048(.A1(new_n221), .A2(new_n224), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n230), .A2(new_n232), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT72), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT28), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n222), .A2(G134), .ZN(new_n240));
  AND2_X1   g054(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n240), .B(KEYINPUT65), .C1(new_n241), .C2(new_n242), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n222), .A2(G134), .ZN(new_n247));
  INV_X1    g061(.A(G134), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(G137), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n247), .B1(KEYINPUT11), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n245), .A2(new_n246), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G131), .ZN(new_n252));
  INV_X1    g066(.A(G131), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n245), .A2(new_n246), .A3(new_n253), .A4(new_n250), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n203), .A2(G143), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G146), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT0), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n256), .B(new_n258), .C1(new_n259), .C2(new_n189), .ZN(new_n260));
  XOR2_X1   g074(.A(KEYINPUT0), .B(G128), .Z(new_n261));
  XNOR2_X1  g075(.A(G143), .B(G146), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n265), .B1(new_n187), .B2(G116), .ZN(new_n266));
  INV_X1    g080(.A(G116), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT67), .A3(G119), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n187), .A2(G116), .ZN(new_n270));
  INV_X1    g084(.A(G113), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT2), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT2), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G113), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n269), .A2(new_n270), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n275), .B1(new_n269), .B2(new_n270), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n278));
  NOR3_X1   g092(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n267), .A2(KEYINPUT67), .A3(G119), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT67), .B1(new_n267), .B2(G119), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n270), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n275), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n269), .A2(new_n270), .A3(new_n275), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT68), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n256), .A3(new_n258), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT66), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n257), .A2(G146), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n203), .A2(G143), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G128), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n189), .A2(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n288), .A2(new_n256), .A3(new_n258), .A4(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n290), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G131), .B1(new_n247), .B2(new_n249), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n254), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n264), .A2(new_n287), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n278), .B1(new_n276), .B2(new_n277), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n284), .A2(KEYINPUT68), .A3(new_n285), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n263), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n305), .B1(new_n252), .B2(new_n254), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n254), .A2(new_n298), .A3(new_n299), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n239), .B1(new_n301), .B2(new_n308), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n306), .A2(new_n304), .A3(new_n307), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(KEYINPUT28), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(G101), .ZN(new_n313));
  INV_X1    g127(.A(G237), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n217), .A2(G210), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n313), .B(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n309), .A2(new_n311), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT30), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n264), .A2(new_n319), .A3(new_n300), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT30), .B1(new_n306), .B2(new_n307), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n287), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n317), .B1(new_n322), .B2(new_n310), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n318), .B1(KEYINPUT71), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n309), .ZN(new_n325));
  INV_X1    g139(.A(new_n311), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n325), .A2(KEYINPUT71), .A3(new_n326), .A4(new_n316), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n238), .B1(new_n324), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT29), .B1(new_n318), .B2(KEYINPUT71), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n323), .A2(KEYINPUT71), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n331), .B(KEYINPUT72), .C1(new_n332), .C2(new_n318), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n309), .A2(KEYINPUT73), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n325), .A2(new_n326), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n334), .B1(new_n335), .B2(KEYINPUT73), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n317), .A2(new_n328), .ZN(new_n337));
  AOI21_X1  g151(.A(G902), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n330), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n339), .A2(G472), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n309), .A2(new_n311), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(new_n316), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n319), .B1(new_n264), .B2(new_n300), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT30), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n304), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT70), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n301), .A4(new_n316), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT31), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n320), .A2(new_n321), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n310), .B1(new_n350), .B2(new_n304), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n351), .A2(new_n346), .A3(KEYINPUT31), .A4(new_n316), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n342), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT32), .ZN(new_n354));
  NOR2_X1   g168(.A1(G472), .A2(G902), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n354), .B1(new_n353), .B2(new_n356), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n237), .B1(new_n340), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT79), .ZN(new_n362));
  INV_X1    g176(.A(new_n237), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n349), .A2(new_n352), .ZN(new_n364));
  INV_X1    g178(.A(new_n342), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT32), .B1(new_n366), .B2(new_n355), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(new_n357), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n339), .A2(G472), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n363), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT79), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n362), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT9), .B(G234), .ZN(new_n374));
  OAI21_X1  g188(.A(G221), .B1(new_n374), .B2(G902), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n375), .B(KEYINPUT80), .Z(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G469), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(new_n225), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT86), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n381));
  XNOR2_X1  g195(.A(G104), .B(G107), .ZN(new_n382));
  INV_X1    g196(.A(G101), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT82), .B(G101), .ZN(new_n385));
  INV_X1    g199(.A(G104), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G107), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n388));
  INV_X1    g202(.A(G107), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(G104), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT3), .B1(new_n386), .B2(G107), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n385), .A2(new_n387), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(G104), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n387), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(KEYINPUT83), .A3(G101), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n384), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n380), .B1(new_n396), .B2(new_n298), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n298), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n290), .A2(new_n297), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n384), .A2(new_n392), .A3(new_n395), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n399), .A2(new_n400), .A3(KEYINPUT86), .A4(new_n295), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT85), .B1(new_n252), .B2(new_n254), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT12), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n406));
  OR2_X1    g220(.A1(new_n406), .A2(KEYINPUT10), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n396), .A2(new_n298), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(KEYINPUT10), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n255), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n391), .A2(new_n390), .A3(new_n387), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n412), .A2(new_n413), .A3(G101), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n391), .A2(new_n390), .A3(new_n387), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n413), .B1(new_n415), .B2(new_n385), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(G101), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n263), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n396), .A2(new_n406), .A3(KEYINPUT10), .A4(new_n298), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n410), .A2(new_n411), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT12), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n402), .A2(new_n422), .A3(new_n403), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n405), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G110), .B(G140), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT81), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n217), .A2(G227), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n408), .A2(new_n409), .B1(new_n418), .B2(new_n263), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n420), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n255), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n421), .A2(new_n428), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n424), .A2(new_n429), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n379), .B1(new_n434), .B2(G469), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n433), .A2(new_n405), .A3(new_n423), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n428), .B1(new_n432), .B2(new_n421), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n378), .B(new_n225), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n377), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G214), .B1(G237), .B2(G902), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT90), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n290), .A2(new_n295), .A3(new_n205), .A4(new_n297), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n260), .B(G125), .C1(new_n261), .C2(new_n262), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n441), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G224), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n447), .B1(new_n448), .B2(G953), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(G953), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n444), .B2(new_n446), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G122), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT88), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT87), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n304), .A2(new_n458), .A3(new_n418), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n458), .B1(new_n304), .B2(new_n418), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g275(.A(KEYINPUT5), .B(new_n270), .C1(new_n280), .C2(new_n281), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n270), .A2(KEYINPUT5), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(G113), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n285), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(new_n400), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n457), .B1(new_n461), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n418), .B1(new_n279), .B2(new_n286), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT87), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n304), .A2(new_n458), .A3(new_n418), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n470), .A2(new_n457), .A3(new_n467), .A4(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n456), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n461), .A2(new_n475), .A3(new_n455), .A4(new_n467), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n470), .A2(new_n455), .A3(new_n467), .A4(new_n471), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT89), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n454), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n470), .A2(new_n467), .A3(new_n471), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT88), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n455), .B1(new_n482), .B2(new_n472), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(KEYINPUT6), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n453), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT93), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n442), .A2(new_n443), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT90), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n450), .A2(KEYINPUT91), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT7), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(new_n450), .B2(KEYINPUT91), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n488), .A2(new_n445), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT92), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n447), .A2(KEYINPUT92), .A3(new_n489), .A4(new_n491), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n455), .B(KEYINPUT8), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n383), .B1(new_n387), .B2(new_n393), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n415), .A2(new_n385), .B1(KEYINPUT83), .B2(new_n498), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n384), .A2(new_n499), .B1(new_n464), .B2(new_n285), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n497), .B1(new_n466), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n490), .B1(new_n444), .B2(new_n446), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n501), .A2(new_n451), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(new_n476), .B2(new_n478), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n486), .B1(new_n505), .B2(G902), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n496), .A2(new_n503), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n479), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(KEYINPUT93), .A3(new_n225), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G210), .B1(G237), .B2(G902), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n485), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n511), .B1(new_n485), .B2(new_n510), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n439), .B(new_n440), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n217), .A2(G214), .A3(new_n314), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n515), .A2(new_n257), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n257), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G131), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(new_n253), .A3(new_n517), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n211), .A2(new_n208), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n518), .A2(KEYINPUT17), .A3(G131), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n202), .B(new_n203), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(new_n253), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n526), .B1(new_n518), .B2(new_n528), .ZN(new_n529));
  AOI211_X1 g343(.A(new_n527), .B(new_n253), .C1(new_n516), .C2(new_n517), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(G113), .B(G122), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(new_n386), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n532), .B(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(G475), .B1(new_n535), .B2(G902), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n525), .A2(new_n531), .A3(new_n534), .ZN(new_n537));
  INV_X1    g351(.A(new_n534), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT19), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n202), .B1(KEYINPUT94), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(KEYINPUT94), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n208), .B1(new_n542), .B2(G146), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n543), .B1(new_n519), .B2(new_n521), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n529), .A2(new_n530), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n538), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n537), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT97), .ZN(new_n548));
  NOR2_X1   g362(.A1(G475), .A2(G902), .ZN(new_n549));
  XOR2_X1   g363(.A(new_n549), .B(KEYINPUT95), .Z(new_n550));
  OR2_X1    g364(.A1(new_n550), .A2(KEYINPUT96), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT20), .B1(new_n550), .B2(KEYINPUT96), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n547), .A2(new_n548), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT20), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n550), .B1(new_n537), .B2(new_n546), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n552), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n537), .B2(new_n546), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n548), .B1(new_n558), .B2(new_n551), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n536), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(G128), .B(G143), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT13), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n257), .A2(G128), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n562), .B(G134), .C1(KEYINPUT13), .C2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(G116), .B(G122), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(new_n389), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n561), .A2(new_n248), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n561), .B(new_n248), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n267), .A2(KEYINPUT14), .A3(G122), .ZN(new_n570));
  INV_X1    g384(.A(new_n565), .ZN(new_n571));
  OAI211_X1 g385(.A(G107), .B(new_n570), .C1(new_n571), .C2(KEYINPUT14), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n569), .B(new_n572), .C1(G107), .C2(new_n571), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n374), .A2(new_n231), .A3(G953), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n568), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n573), .B2(new_n568), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(KEYINPUT98), .A3(new_n225), .ZN(new_n578));
  INV_X1    g392(.A(G478), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(KEYINPUT15), .ZN(new_n580));
  XOR2_X1   g394(.A(new_n578), .B(new_n580), .Z(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G952), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(G953), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(G234), .B2(G237), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI211_X1 g401(.A(new_n225), .B(new_n217), .C1(G234), .C2(G237), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT21), .B(G898), .Z(new_n590));
  OAI21_X1  g404(.A(new_n587), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n591), .B(KEYINPUT99), .Z(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n560), .A2(new_n582), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n514), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n373), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n597), .B(new_n385), .Z(G3));
  INV_X1    g412(.A(new_n440), .ZN(new_n599));
  INV_X1    g413(.A(new_n511), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT93), .B1(new_n508), .B2(new_n225), .ZN(new_n601));
  AOI211_X1 g415(.A(new_n486), .B(G902), .C1(new_n479), .C2(new_n507), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n477), .B(new_n475), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT6), .B1(new_n604), .B2(new_n483), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n474), .A2(new_n454), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n452), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n600), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n485), .A2(new_n510), .A3(new_n511), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n599), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n353), .A2(new_n356), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n366), .A2(new_n225), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n611), .B1(new_n612), .B2(G472), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n613), .A2(KEYINPUT100), .A3(new_n439), .A4(new_n237), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n366), .A2(new_n355), .ZN(new_n615));
  OAI21_X1  g429(.A(G472), .B1(new_n353), .B2(G902), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n237), .A2(new_n615), .A3(new_n616), .A4(new_n439), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n610), .A2(new_n614), .A3(new_n619), .A4(new_n592), .ZN(new_n620));
  INV_X1    g434(.A(new_n560), .ZN(new_n621));
  AOI21_X1  g435(.A(G478), .B1(new_n577), .B2(new_n225), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT101), .B1(new_n575), .B2(new_n576), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT33), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(G902), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n622), .B1(new_n628), .B2(G478), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n620), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT34), .B(G104), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  NOR2_X1   g448(.A1(new_n555), .A2(new_n554), .ZN(new_n635));
  INV_X1    g449(.A(new_n550), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n547), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(KEYINPUT20), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n536), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n620), .A2(new_n581), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT35), .B(G107), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  INV_X1    g456(.A(new_n613), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n514), .A2(new_n595), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n229), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT25), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n232), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n220), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(new_n216), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n234), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n644), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT37), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(new_n214), .ZN(G12));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n586), .B1(new_n588), .B2(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n639), .A2(new_n581), .A3(new_n656), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n440), .B(new_n657), .C1(new_n512), .C2(new_n513), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT102), .ZN(new_n659));
  INV_X1    g473(.A(new_n439), .ZN(new_n660));
  INV_X1    g474(.A(new_n651), .ZN(new_n661));
  AOI211_X1 g475(.A(new_n660), .B(new_n661), .C1(new_n368), .C2(new_n369), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n608), .A2(new_n609), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n663), .A2(new_n664), .A3(new_n440), .A4(new_n657), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n659), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  NAND2_X1  g481(.A1(new_n560), .A2(new_n582), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n656), .B(KEYINPUT104), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT39), .Z(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n439), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n669), .B1(KEYINPUT40), .B2(new_n673), .ZN(new_n674));
  AOI211_X1 g488(.A(new_n599), .B(new_n674), .C1(KEYINPUT40), .C2(new_n673), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n351), .A2(new_n316), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n301), .A2(new_n308), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(KEYINPUT103), .A3(new_n317), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT103), .B1(new_n677), .B2(new_n317), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n225), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(G472), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n368), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n663), .B(KEYINPUT38), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n675), .A2(new_n661), .A3(new_n683), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT105), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  NAND3_X1  g501(.A1(new_n547), .A2(new_n551), .A3(new_n552), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT97), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n637), .A2(KEYINPUT20), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n690), .A3(new_n553), .ZN(new_n691));
  AOI211_X1 g505(.A(new_n629), .B(new_n656), .C1(new_n691), .C2(new_n536), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n440), .B(new_n692), .C1(new_n512), .C2(new_n513), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n662), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  AOI211_X1 g510(.A(new_n599), .B(new_n593), .C1(new_n608), .C2(new_n609), .ZN(new_n697));
  INV_X1    g511(.A(new_n375), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n405), .A2(new_n423), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n432), .A2(new_n421), .ZN(new_n700));
  AOI22_X1  g514(.A1(new_n699), .A2(new_n433), .B1(new_n700), .B2(new_n429), .ZN(new_n701));
  OAI21_X1  g515(.A(G469), .B1(new_n701), .B2(G902), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(KEYINPUT106), .A3(new_n438), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n704), .B(G469), .C1(new_n701), .C2(G902), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n698), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n697), .A2(new_n370), .A3(new_n630), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NOR2_X1   g523(.A1(new_n639), .A2(new_n581), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n697), .A2(new_n370), .A3(new_n710), .A4(new_n706), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  AOI21_X1  g526(.A(new_n661), .B1(new_n368), .B2(new_n369), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n713), .A2(new_n610), .A3(new_n594), .A4(new_n706), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  OAI21_X1  g529(.A(new_n364), .B1(new_n316), .B2(new_n336), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n355), .ZN(new_n717));
  AND4_X1   g531(.A1(new_n592), .A2(new_n717), .A3(new_n237), .A4(new_n616), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n610), .A2(new_n669), .A3(new_n706), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G122), .ZN(G24));
  NAND4_X1  g534(.A1(new_n706), .A2(new_n616), .A3(new_n651), .A4(new_n717), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT107), .B1(new_n693), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n438), .A2(KEYINPUT106), .ZN(new_n723));
  INV_X1    g537(.A(new_n437), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n433), .A2(new_n405), .A3(new_n423), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n378), .B1(new_n726), .B2(new_n225), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n705), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n375), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n717), .A2(new_n616), .A3(new_n651), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n610), .A3(new_n733), .A4(new_n692), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n722), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  NAND4_X1  g550(.A1(new_n608), .A2(new_n375), .A3(new_n440), .A4(new_n609), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n435), .A2(new_n438), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n738), .A2(new_n739), .A3(new_n370), .A4(new_n692), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT42), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT108), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n359), .A2(new_n742), .ZN(new_n743));
  OAI211_X1 g557(.A(KEYINPUT108), .B(new_n354), .C1(new_n353), .C2(new_n356), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n357), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI211_X1 g559(.A(new_n741), .B(new_n363), .C1(new_n745), .C2(new_n369), .ZN(new_n746));
  INV_X1    g560(.A(new_n739), .ZN(new_n747));
  INV_X1    g561(.A(new_n629), .ZN(new_n748));
  INV_X1    g562(.A(new_n656), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n560), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n737), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n740), .A2(new_n741), .B1(new_n746), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n253), .ZN(G33));
  NOR2_X1   g567(.A1(new_n737), .A2(new_n747), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n370), .A3(new_n657), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n434), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(G469), .ZN(new_n759));
  INV_X1    g573(.A(new_n379), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(KEYINPUT46), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n762), .B(G469), .C1(new_n758), .C2(G902), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(new_n438), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n375), .A3(new_n672), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n629), .B(KEYINPUT109), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n621), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n621), .A2(KEYINPUT110), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n560), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n629), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n768), .B(new_n643), .C1(new_n772), .C2(new_n767), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n773), .A2(new_n661), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n765), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n773), .A2(new_n661), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n608), .A2(new_n440), .A3(new_n609), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n779), .A2(KEYINPUT111), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(KEYINPUT111), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n777), .A2(KEYINPUT44), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  NAND3_X1  g598(.A1(new_n368), .A2(new_n692), .A3(new_n369), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n764), .A2(new_n375), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT47), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n764), .A2(KEYINPUT47), .A3(new_n375), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n785), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n779), .A2(new_n237), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT112), .Z(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  NOR2_X1   g608(.A1(new_n728), .A2(new_n729), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT49), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n684), .A2(new_n377), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n683), .A2(new_n363), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n440), .A3(new_n772), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n711), .A2(new_n714), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n630), .B1(new_n582), .B2(new_n621), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n719), .B1(new_n620), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n373), .A2(new_n596), .B1(new_n644), .B2(new_n651), .ZN(new_n805));
  INV_X1    g619(.A(new_n731), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n751), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n804), .A2(new_n805), .A3(new_n707), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n809));
  INV_X1    g623(.A(new_n639), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n582), .A2(new_n656), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n778), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n608), .A2(new_n810), .A3(new_n440), .A4(new_n609), .ZN(new_n813));
  INV_X1    g627(.A(new_n811), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT113), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n662), .A3(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n740), .A2(new_n741), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n746), .A2(new_n751), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n755), .B(new_n816), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n808), .A2(new_n819), .ZN(new_n820));
  AOI211_X1 g634(.A(new_n599), .B(new_n668), .C1(new_n608), .C2(new_n609), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n651), .A2(new_n656), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n375), .A3(new_n739), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT114), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n822), .A2(new_n825), .A3(new_n375), .A4(new_n739), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n821), .A2(new_n683), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n735), .A2(new_n666), .A3(new_n695), .A4(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n722), .A2(new_n734), .B1(new_n694), .B2(new_n662), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(KEYINPUT52), .A3(new_n666), .A4(new_n827), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n831), .B1(new_n830), .B2(new_n833), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n820), .B(KEYINPUT53), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n812), .A2(new_n662), .A3(new_n815), .ZN(new_n838));
  INV_X1    g652(.A(new_n755), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n752), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n707), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n801), .A2(new_n803), .A3(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n840), .A2(new_n807), .A3(new_n842), .A4(new_n805), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n830), .A2(new_n833), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n837), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n800), .B1(new_n836), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n820), .A2(KEYINPUT53), .A3(new_n844), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n844), .A2(KEYINPUT115), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n843), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n800), .B(new_n848), .C1(new_n851), .C2(KEYINPUT53), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n847), .B1(new_n852), .B2(KEYINPUT116), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n847), .A2(KEYINPUT116), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n768), .B1(new_n772), .B2(new_n767), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n717), .A2(new_n616), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n855), .A2(new_n587), .A3(new_n363), .A4(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(KEYINPUT118), .A3(new_n610), .A4(new_n706), .ZN(new_n858));
  OR3_X1    g672(.A1(new_n737), .A2(new_n587), .A3(new_n795), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n859), .A2(new_n363), .A3(new_n683), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n585), .B1(new_n860), .B2(new_n630), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n862));
  INV_X1    g676(.A(new_n855), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n856), .A2(new_n363), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n586), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n610), .A2(new_n706), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n858), .A2(new_n861), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n859), .A2(new_n855), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n363), .B1(new_n745), .B2(new_n369), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(KEYINPUT120), .B2(KEYINPUT48), .ZN(new_n875));
  XNOR2_X1  g689(.A(KEYINPUT120), .B(KEYINPUT48), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n875), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n870), .A2(new_n871), .A3(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n859), .A2(new_n855), .A3(new_n731), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n860), .A2(new_n621), .A3(new_n629), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n788), .B(new_n789), .C1(new_n376), .C2(new_n795), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n865), .B1(new_n781), .B2(new_n780), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n879), .B(new_n880), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n684), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n706), .A2(new_n599), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT117), .Z(new_n886));
  NAND3_X1  g700(.A1(new_n857), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT50), .Z(new_n888));
  INV_X1    g702(.A(KEYINPUT51), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n883), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n889), .B1(new_n883), .B2(new_n888), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n878), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n853), .A2(new_n854), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(G952), .A2(G953), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n799), .B1(new_n893), .B2(new_n894), .ZN(G75));
  OAI21_X1  g709(.A(new_n820), .B1(new_n834), .B2(new_n835), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n837), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n848), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(G210), .A3(G902), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT56), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n480), .A2(new_n453), .A3(new_n484), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(new_n607), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT55), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n899), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n903), .B1(new_n899), .B2(new_n900), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n217), .A2(G952), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(G51));
  NAND2_X1  g721(.A1(new_n760), .A2(KEYINPUT57), .ZN(new_n908));
  INV_X1    g722(.A(new_n852), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n800), .B1(new_n897), .B2(new_n848), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n760), .A2(KEYINPUT57), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n726), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n898), .A2(G469), .A3(G902), .A4(new_n758), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n906), .B1(new_n913), .B2(new_n914), .ZN(G54));
  AND2_X1   g729(.A1(KEYINPUT58), .A2(G475), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(KEYINPUT121), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(KEYINPUT121), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n898), .A2(G902), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n547), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n921), .A2(new_n922), .A3(new_n906), .ZN(G60));
  INV_X1    g737(.A(new_n625), .ZN(new_n924));
  INV_X1    g738(.A(new_n627), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT59), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n927), .B(new_n929), .C1(new_n909), .C2(new_n910), .ZN(new_n930));
  INV_X1    g744(.A(new_n906), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n929), .B1(new_n853), .B2(new_n854), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n926), .B2(new_n933), .ZN(G63));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n935));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT122), .Z(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT60), .Z(new_n938));
  NAND3_X1  g752(.A1(new_n898), .A2(new_n649), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n931), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n236), .B1(new_n898), .B2(new_n938), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n935), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n941), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n943), .A2(KEYINPUT61), .A3(new_n931), .A4(new_n939), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(G66));
  INV_X1    g759(.A(new_n590), .ZN(new_n946));
  OAI21_X1  g760(.A(G953), .B1(new_n946), .B2(new_n448), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n842), .A2(new_n805), .ZN(new_n948));
  INV_X1    g762(.A(new_n217), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n605), .B(new_n606), .C1(G898), .C2(new_n217), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G69));
  AOI22_X1  g766(.A1(new_n776), .A2(new_n782), .B1(new_n791), .B2(new_n790), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n752), .A2(new_n839), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n832), .A2(new_n666), .ZN(new_n955));
  INV_X1    g769(.A(new_n765), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(new_n873), .A3(new_n821), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n953), .A2(new_n954), .A3(new_n955), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n217), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n949), .A2(KEYINPUT125), .A3(new_n655), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n949), .A2(new_n655), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n959), .A2(new_n960), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT126), .ZN(new_n965));
  AOI22_X1  g779(.A1(new_n958), .A2(new_n217), .B1(new_n962), .B2(new_n961), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n966), .A2(new_n967), .A3(new_n960), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n350), .B(new_n542), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n217), .B1(G227), .B2(G900), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n955), .A2(new_n685), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT62), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n783), .A2(new_n792), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n673), .B1(new_n362), .B2(new_n372), .ZN(new_n978));
  INV_X1    g792(.A(new_n802), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n779), .B1(new_n979), .B2(KEYINPUT123), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n978), .B(new_n980), .C1(KEYINPUT123), .C2(new_n979), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT124), .Z(new_n982));
  NOR3_X1   g796(.A1(new_n976), .A2(new_n977), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n970), .B1(new_n983), .B2(new_n949), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n972), .A2(new_n974), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n970), .B1(new_n965), .B2(new_n968), .ZN(new_n986));
  INV_X1    g800(.A(new_n984), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n973), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n985), .A2(new_n988), .ZN(G72));
  NAND2_X1  g803(.A1(new_n676), .A2(new_n323), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n958), .A2(new_n317), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n948), .B(new_n991), .C1(new_n983), .C2(new_n351), .ZN(new_n992));
  XOR2_X1   g806(.A(KEYINPUT127), .B(KEYINPUT63), .Z(new_n993));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n990), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n990), .A2(new_n995), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n997), .B1(new_n836), .B2(new_n846), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n996), .A2(new_n906), .A3(new_n998), .ZN(G57));
endmodule


