//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT22), .ZN(new_n207));
  INV_X1    g006(.A(G211gat), .ZN(new_n208));
  INV_X1    g007(.A(G218gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT72), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(new_n206), .A3(new_n210), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n211), .A2(KEYINPUT72), .A3(new_n213), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT27), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT27), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(G190gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT68), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(KEYINPUT28), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n222), .A2(G183gat), .ZN(new_n233));
  INV_X1    g032(.A(G183gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT27), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n233), .A2(new_n235), .A3(KEYINPUT69), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT69), .B1(new_n233), .B2(new_n235), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n232), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n228), .A2(new_n230), .A3(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT26), .ZN(new_n242));
  NAND2_X1  g041(.A1(G169gat), .A2(G176gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n240), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n239), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT64), .B1(new_n241), .B2(KEYINPUT23), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT23), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n249), .B(new_n250), .C1(G169gat), .C2(G176gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n224), .A2(G183gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n234), .A2(G190gat), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT24), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT24), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n256), .A2(new_n240), .B1(new_n241), .B2(KEYINPUT23), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n252), .A2(new_n255), .A3(new_n245), .A4(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT25), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n241), .A2(KEYINPUT23), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n256), .A2(G183gat), .A3(G190gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n243), .A2(new_n244), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n261), .B(new_n262), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n266), .A2(KEYINPUT25), .A3(new_n252), .A4(new_n255), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G226gat), .A2(G233gat), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n247), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n269), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(KEYINPUT29), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n272), .B1(new_n247), .B2(new_n268), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n219), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n247), .A2(new_n268), .A3(new_n269), .ZN(new_n275));
  INV_X1    g074(.A(new_n219), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n239), .A2(new_n246), .B1(new_n260), .B2(new_n267), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n275), .B(new_n276), .C1(new_n277), .C2(new_n272), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n274), .A2(KEYINPUT73), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n280), .B(new_n219), .C1(new_n270), .C2(new_n273), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n205), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(KEYINPUT86), .B(KEYINPUT37), .Z(new_n283));
  AOI21_X1  g082(.A(new_n283), .B1(new_n279), .B2(new_n281), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT87), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n204), .A2(KEYINPUT38), .ZN(new_n287));
  INV_X1    g086(.A(new_n274), .ZN(new_n288));
  INV_X1    g087(.A(new_n278), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT37), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT85), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT85), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n292), .B(KEYINPUT37), .C1(new_n288), .C2(new_n289), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n287), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n282), .B1(new_n286), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G1gat), .B(G29gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT0), .ZN(new_n297));
  XNOR2_X1  g096(.A(G57gat), .B(G85gat), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n297), .B(new_n298), .Z(new_n299));
  XOR2_X1   g098(.A(KEYINPUT79), .B(KEYINPUT6), .Z(new_n300));
  INV_X1    g099(.A(KEYINPUT1), .ZN(new_n301));
  AND2_X1   g100(.A1(G113gat), .A2(G120gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(G113gat), .A2(G120gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(G127gat), .A2(G134gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(G127gat), .A2(G134gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n301), .B(new_n304), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G113gat), .ZN(new_n310));
  INV_X1    g109(.A(G120gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G113gat), .A2(G120gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(new_n301), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n308), .A3(new_n313), .ZN(new_n315));
  XNOR2_X1  g114(.A(G127gat), .B(G134gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n309), .A2(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G141gat), .B(G148gat), .Z(new_n319));
  XNOR2_X1  g118(.A(G155gat), .B(G162gat), .ZN(new_n320));
  INV_X1    g119(.A(G155gat), .ZN(new_n321));
  INV_X1    g120(.A(G162gat), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT2), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n322), .ZN(new_n326));
  XNOR2_X1  g125(.A(G141gat), .B(G148gat), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n325), .B(new_n326), .C1(new_n327), .C2(KEYINPUT2), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT75), .B(KEYINPUT3), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n324), .A2(new_n328), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n318), .B(new_n330), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n309), .A2(new_n317), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT4), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n328), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT76), .B1(new_n318), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n331), .A2(new_n336), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n338), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n318), .A2(new_n341), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n342), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n334), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT77), .B1(new_n350), .B2(KEYINPUT5), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT5), .ZN(new_n353));
  AOI211_X1 g152(.A(new_n352), .B(new_n353), .C1(new_n348), .C2(new_n349), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n346), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n342), .A2(KEYINPUT4), .A3(new_n344), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n356), .B(new_n357), .C1(KEYINPUT4), .C2(new_n337), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n342), .A2(new_n344), .A3(KEYINPUT78), .A4(KEYINPUT4), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n335), .A2(KEYINPUT5), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI211_X1 g160(.A(new_n299), .B(new_n300), .C1(new_n355), .C2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n345), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n363), .A2(new_n335), .A3(new_n339), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n350), .A2(KEYINPUT5), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n352), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n350), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n361), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT84), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n299), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT84), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n372), .A3(new_n361), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n355), .A2(new_n361), .A3(new_n299), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n300), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n362), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n279), .A2(KEYINPUT37), .A3(new_n281), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n279), .A2(new_n281), .ZN(new_n380));
  INV_X1    g179(.A(new_n283), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n285), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AOI211_X1 g181(.A(KEYINPUT87), .B(new_n283), .C1(new_n279), .C2(new_n281), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n205), .B(new_n379), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT38), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n295), .A2(new_n378), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n330), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n219), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G228gat), .A2(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n217), .A2(new_n387), .A3(new_n218), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n331), .B1(new_n393), .B2(new_n332), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n390), .B(KEYINPUT80), .Z(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT29), .B1(new_n214), .B2(new_n216), .ZN(new_n398));
  INV_X1    g197(.A(new_n329), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n341), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n397), .B1(new_n389), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(G22gat), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n214), .A2(new_n216), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n387), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n331), .B1(new_n405), .B2(new_n329), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n217), .A2(new_n218), .B1(new_n330), .B2(new_n387), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n396), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(G22gat), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n408), .B(new_n409), .C1(new_n394), .C2(new_n392), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n402), .A2(new_n403), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT82), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n402), .A2(new_n403), .A3(new_n410), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n402), .A2(new_n410), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT81), .ZN(new_n417));
  XNOR2_X1  g216(.A(G78gat), .B(G106gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT31), .B(G50gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n412), .A2(new_n417), .A3(new_n420), .A4(new_n414), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n355), .A2(new_n361), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n299), .B1(new_n425), .B2(KEYINPUT84), .ZN(new_n426));
  INV_X1    g225(.A(new_n356), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n357), .B1(new_n337), .B2(KEYINPUT4), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n359), .B(new_n333), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT39), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n430), .A3(new_n349), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n299), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n348), .A2(new_n349), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT39), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n434), .B1(new_n349), .B2(new_n429), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT40), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n429), .A2(new_n349), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(KEYINPUT39), .A3(new_n433), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT40), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n299), .A4(new_n431), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n426), .A2(new_n373), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n380), .A2(KEYINPUT30), .A3(new_n204), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n279), .A2(new_n281), .A3(new_n205), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT74), .B(KEYINPUT30), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n442), .B(new_n443), .C1(new_n282), .C2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n424), .B1(new_n441), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n386), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT83), .ZN(new_n449));
  INV_X1    g248(.A(new_n300), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n425), .A2(new_n371), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n299), .B1(new_n355), .B2(new_n361), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n451), .B1(new_n376), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n282), .A2(new_n445), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT30), .ZN(new_n455));
  AOI211_X1 g254(.A(new_n455), .B(new_n205), .C1(new_n279), .C2(new_n281), .ZN(new_n456));
  INV_X1    g255(.A(new_n443), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n454), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n453), .A2(new_n458), .B1(new_n423), .B2(new_n422), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n260), .A2(new_n267), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n242), .A2(new_n245), .ZN(new_n462));
  INV_X1    g261(.A(new_n240), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT69), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n234), .A2(KEYINPUT27), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n222), .A2(G183gat), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n233), .A2(new_n235), .A3(KEYINPUT69), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n231), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n229), .B1(new_n225), .B2(new_n226), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n464), .B1(new_n472), .B2(new_n230), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n336), .B1(new_n461), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G227gat), .ZN(new_n475));
  INV_X1    g274(.A(G233gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n247), .A2(new_n268), .A3(new_n318), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n474), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT32), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT33), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(G15gat), .B(G43gat), .Z(new_n483));
  XNOR2_X1  g282(.A(G71gat), .B(G99gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n480), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n485), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n479), .B(KEYINPUT32), .C1(new_n481), .C2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n477), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT34), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(KEYINPUT71), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n277), .A2(new_n318), .ZN(new_n492));
  INV_X1    g291(.A(new_n478), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n489), .B(new_n491), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n477), .B1(new_n474), .B2(new_n478), .ZN(new_n495));
  XOR2_X1   g294(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n486), .A2(new_n488), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n497), .B1(new_n486), .B2(new_n488), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n460), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n486), .A2(new_n488), .ZN(new_n501));
  INV_X1    g300(.A(new_n497), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n497), .A3(new_n488), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(KEYINPUT36), .A3(new_n504), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n449), .B1(new_n459), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n500), .A2(new_n505), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n425), .A2(new_n371), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n509), .A2(new_n300), .A3(new_n375), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n446), .B1(new_n510), .B2(new_n451), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n422), .A2(new_n423), .ZN(new_n512));
  OAI211_X1 g311(.A(KEYINPUT83), .B(new_n508), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n448), .A2(new_n507), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n515), .A2(new_n423), .A3(new_n422), .ZN(new_n516));
  INV_X1    g315(.A(new_n454), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT35), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n517), .A2(new_n518), .A3(new_n443), .A4(new_n442), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n378), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n453), .A2(new_n458), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT35), .B1(new_n523), .B2(new_n516), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n514), .A2(KEYINPUT88), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT88), .B1(new_n514), .B2(new_n525), .ZN(new_n527));
  XNOR2_X1  g326(.A(G43gat), .B(G50gat), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n528), .A2(KEYINPUT15), .ZN(new_n529));
  NOR2_X1   g328(.A1(G29gat), .A2(G36gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT14), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT14), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(G29gat), .B2(G36gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(KEYINPUT91), .B(G36gat), .Z(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT90), .B(G29gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n535), .B(new_n538), .C1(KEYINPUT15), .C2(new_n528), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(KEYINPUT89), .B2(new_n534), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n534), .A2(KEYINPUT89), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n529), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT17), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT92), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(new_n542), .A3(KEYINPUT17), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT93), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G15gat), .B(G22gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT16), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n549), .B1(new_n550), .B2(G1gat), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(G1gat), .B2(new_n549), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(G8gat), .Z(new_n553));
  NAND3_X1  g352(.A1(new_n545), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555));
  INV_X1    g354(.A(new_n553), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n542), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n554), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT18), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n554), .A2(KEYINPUT18), .A3(new_n555), .A4(new_n558), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n553), .B(new_n557), .Z(new_n563));
  XOR2_X1   g362(.A(new_n555), .B(KEYINPUT13), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n561), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G197gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT11), .B(G169gat), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n568), .B(new_n569), .Z(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT12), .Z(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT94), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT94), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n566), .A2(new_n574), .A3(new_n571), .ZN(new_n575));
  INV_X1    g374(.A(new_n571), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n561), .A2(new_n576), .A3(new_n562), .A4(new_n565), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT95), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n559), .A2(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT95), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n576), .A4(new_n562), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n573), .A2(new_n575), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n526), .A2(new_n527), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  NAND2_X1  g385(.A1(G99gat), .A2(G106gat), .ZN(new_n587));
  INV_X1    g386(.A(G85gat), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  AOI22_X1  g388(.A1(KEYINPUT8), .A2(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT102), .ZN(new_n592));
  XOR2_X1   g391(.A(G99gat), .B(G106gat), .Z(new_n593));
  INV_X1    g392(.A(KEYINPUT102), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n586), .A2(new_n594), .A3(new_n590), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n593), .ZN(new_n597));
  INV_X1    g396(.A(new_n595), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n594), .B1(new_n586), .B2(new_n590), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n545), .A2(new_n548), .A3(new_n596), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n596), .ZN(new_n602));
  AND2_X1   g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603));
  AOI22_X1  g402(.A1(new_n602), .A2(new_n557), .B1(KEYINPUT41), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G190gat), .B(G218gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n603), .A2(KEYINPUT41), .ZN(new_n608));
  XNOR2_X1  g407(.A(G134gat), .B(G162gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G71gat), .B(G78gat), .Z(new_n615));
  XOR2_X1   g414(.A(G57gat), .B(G64gat), .Z(new_n616));
  AOI21_X1  g415(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI22_X1  g417(.A1(KEYINPUT96), .A2(new_n615), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(KEYINPUT96), .B2(new_n615), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n616), .A2(new_n621), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n615), .A2(new_n617), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT98), .ZN(new_n629));
  XOR2_X1   g428(.A(G127gat), .B(G155gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT20), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n629), .B(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n553), .B1(new_n626), .B2(new_n627), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT100), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n632), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT99), .B(KEYINPUT19), .Z(new_n636));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G183gat), .B(G211gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n635), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n614), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT103), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G230gat), .A2(G233gat), .ZN(new_n645));
  INV_X1    g444(.A(new_n626), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n598), .A2(new_n597), .A3(new_n599), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n593), .B1(new_n592), .B2(new_n595), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n600), .A2(new_n626), .A3(new_n596), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n652), .A2(KEYINPUT104), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n649), .A2(new_n654), .A3(new_n650), .A4(new_n651), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n602), .A2(KEYINPUT10), .A3(new_n646), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n645), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n649), .A2(new_n651), .ZN(new_n659));
  INV_X1    g458(.A(new_n645), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n658), .A2(new_n661), .A3(new_n665), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n644), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n583), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n453), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(G1gat), .Z(G1324gat));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n583), .A2(new_n446), .A3(new_n672), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n676), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n680), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n677), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(KEYINPUT42), .B2(new_n680), .ZN(G1325gat));
  OAI21_X1  g481(.A(G15gat), .B1(new_n673), .B2(new_n508), .ZN(new_n683));
  INV_X1    g482(.A(new_n515), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n684), .A2(G15gat), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n683), .B1(new_n673), .B2(new_n685), .ZN(G1326gat));
  NOR2_X1   g485(.A1(new_n673), .A2(new_n512), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT43), .B(G22gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  INV_X1    g488(.A(new_n641), .ZN(new_n690));
  INV_X1    g489(.A(new_n614), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n583), .A2(new_n690), .A3(new_n691), .A4(new_n670), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n693));
  INV_X1    g492(.A(new_n453), .ZN(new_n694));
  INV_X1    g493(.A(new_n537), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OR3_X1    g495(.A1(new_n692), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n693), .B1(new_n692), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n514), .A2(new_n525), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT88), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n514), .A2(KEYINPUT88), .A3(new_n525), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n702), .A3(new_n691), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n704), .B1(new_n386), .B2(new_n447), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n511), .A2(new_n512), .A3(new_n515), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n706), .A2(KEYINPUT35), .B1(new_n520), .B2(new_n521), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT108), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n709));
  INV_X1    g508(.A(new_n448), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n525), .B(new_n709), .C1(new_n710), .C2(new_n704), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n614), .A2(KEYINPUT44), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n703), .A2(KEYINPUT44), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n578), .A2(new_n581), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n574), .B1(new_n566), .B2(new_n571), .ZN(new_n716));
  AOI211_X1 g515(.A(KEYINPUT94), .B(new_n576), .C1(new_n579), .C2(new_n562), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n715), .B(KEYINPUT106), .C1(new_n716), .C2(new_n717), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n669), .B(KEYINPUT107), .Z(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n723), .A2(new_n690), .A3(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n714), .A2(new_n453), .A3(new_n726), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n697), .B(new_n698), .C1(new_n727), .C2(new_n695), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT109), .Z(G1328gat));
  NOR3_X1   g528(.A1(new_n692), .A2(new_n458), .A3(new_n536), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(KEYINPUT110), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n536), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n714), .A2(new_n458), .A3(new_n726), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT110), .B(KEYINPUT46), .ZN(new_n735));
  OAI221_X1 g534(.A(new_n732), .B1(new_n733), .B2(new_n734), .C1(new_n730), .C2(new_n735), .ZN(G1329gat));
  NOR2_X1   g535(.A1(new_n714), .A2(new_n726), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n737), .A2(G43gat), .A3(new_n506), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n692), .A2(new_n684), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(G43gat), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g540(.A1(new_n692), .A2(G50gat), .A3(new_n512), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n737), .A2(new_n424), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G50gat), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n745), .A2(new_n746), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n744), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n745), .A2(G50gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n743), .B1(new_n751), .B2(new_n742), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1331gat));
  AND3_X1   g552(.A1(new_n644), .A2(new_n722), .A3(new_n724), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n712), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n694), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g557(.A(new_n458), .B(KEYINPUT112), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  AND2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n760), .B2(new_n761), .ZN(G1333gat));
  NAND3_X1  g563(.A1(new_n756), .A2(G71gat), .A3(new_n506), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n515), .B(KEYINPUT113), .Z(new_n766));
  AND2_X1   g565(.A1(new_n756), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n767), .B2(G71gat), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g568(.A1(new_n756), .A2(new_n424), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G78gat), .ZN(G1335gat));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n722), .A2(new_n690), .A3(new_n669), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n714), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n708), .A2(new_n711), .A3(new_n713), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n526), .A2(new_n527), .A3(new_n614), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n773), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(KEYINPUT114), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n774), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(G85gat), .B1(new_n781), .B2(new_n453), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n722), .A2(new_n690), .A3(new_n691), .A4(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n705), .A2(new_n707), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n783), .B2(new_n784), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT115), .B(KEYINPUT51), .C1(new_n786), .C2(new_n787), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n669), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n694), .A2(new_n588), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n782), .B1(new_n792), .B2(new_n793), .ZN(G1336gat));
  NOR2_X1   g593(.A1(new_n759), .A2(G92gat), .ZN(new_n795));
  AND4_X1   g594(.A1(new_n724), .A2(new_n789), .A3(new_n790), .A4(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n714), .A2(new_n759), .A3(new_n773), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n589), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n774), .A2(new_n780), .A3(new_n446), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G92gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n797), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT116), .B1(new_n803), .B2(KEYINPUT52), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n796), .B1(new_n801), .B2(G92gat), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n805), .A2(new_n806), .A3(new_n798), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n800), .B1(new_n804), .B2(new_n807), .ZN(G1337gat));
  OAI21_X1  g607(.A(G99gat), .B1(new_n781), .B2(new_n508), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n684), .A2(G99gat), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n792), .B2(new_n810), .ZN(G1338gat));
  NOR2_X1   g610(.A1(new_n512), .A2(G106gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n791), .A2(new_n724), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814));
  XNOR2_X1  g613(.A(KEYINPUT117), .B(G106gat), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n714), .A2(new_n512), .A3(new_n773), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n813), .B(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n815), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n781), .B2(new_n512), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(new_n813), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n817), .B1(new_n820), .B2(new_n814), .ZN(G1339gat));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n652), .A2(KEYINPUT104), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n823), .A2(new_n660), .A3(new_n656), .A4(new_n655), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n658), .A2(KEYINPUT54), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n826), .B(new_n645), .C1(new_n653), .C2(new_n657), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n666), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n822), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n668), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n827), .A2(new_n666), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n658), .A2(KEYINPUT54), .A3(new_n824), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(KEYINPUT55), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT118), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n831), .A2(new_n835), .A3(KEYINPUT55), .A4(new_n832), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n830), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n720), .A2(new_n721), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n555), .B1(new_n554), .B2(new_n558), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n563), .A2(new_n564), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n570), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT119), .Z(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n715), .A3(new_n669), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n691), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n837), .A2(new_n691), .A3(new_n715), .A4(new_n842), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n690), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n644), .A2(new_n670), .A3(new_n722), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n424), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n759), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n694), .A2(new_n515), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n310), .A3(new_n723), .ZN(new_n855));
  OAI21_X1  g654(.A(G113gat), .B1(new_n853), .B2(new_n582), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(G1340gat));
  NOR3_X1   g659(.A1(new_n853), .A2(new_n311), .A3(new_n725), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n854), .A2(new_n669), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n311), .B2(new_n862), .ZN(G1341gat));
  NAND2_X1  g662(.A1(new_n854), .A2(new_n641), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(G127gat), .ZN(G1342gat));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(KEYINPUT56), .ZN(new_n867));
  NOR4_X1   g666(.A1(new_n614), .A2(new_n851), .A3(G134gat), .A4(new_n446), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n849), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(KEYINPUT56), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n869), .B(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(G134gat), .B1(new_n853), .B2(new_n614), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(G1343gat));
  NAND2_X1  g675(.A1(new_n834), .A2(new_n836), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n829), .A2(new_n668), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n843), .B1(new_n879), .B2(new_n582), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(KEYINPUT123), .B(new_n843), .C1(new_n879), .C2(new_n582), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n614), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n641), .B1(new_n884), .B2(new_n845), .ZN(new_n885));
  INV_X1    g684(.A(new_n848), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n424), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT57), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n512), .B1(new_n847), .B2(new_n848), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n508), .A2(new_n694), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n850), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n888), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n723), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n889), .A2(new_n893), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n582), .A2(G141gat), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n895), .A2(G141gat), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT58), .ZN(new_n899));
  INV_X1    g698(.A(G141gat), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n900), .B1(new_n894), .B2(new_n718), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n896), .A2(new_n897), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n899), .ZN(new_n903));
  OAI22_X1  g702(.A1(new_n898), .A2(new_n899), .B1(new_n901), .B2(new_n903), .ZN(G1344gat));
  INV_X1    g703(.A(G148gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n896), .A2(new_n905), .A3(new_n669), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n847), .A2(new_n848), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(KEYINPUT57), .A3(new_n424), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT124), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n889), .A2(new_n911), .A3(KEYINPUT57), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n671), .A2(new_n718), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n424), .B1(new_n885), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n890), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n910), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n669), .A3(new_n893), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n907), .B1(new_n917), .B2(G148gat), .ZN(new_n918));
  AOI211_X1 g717(.A(KEYINPUT59), .B(new_n905), .C1(new_n894), .C2(new_n669), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n906), .B1(new_n918), .B2(new_n919), .ZN(G1345gat));
  NAND3_X1  g719(.A1(new_n896), .A2(new_n321), .A3(new_n641), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n894), .A2(new_n641), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n321), .ZN(G1346gat));
  NOR4_X1   g722(.A1(new_n614), .A2(new_n892), .A3(G162gat), .A4(new_n446), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n889), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n894), .A2(new_n691), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n322), .ZN(G1347gat));
  AOI21_X1  g726(.A(new_n694), .B1(new_n847), .B2(new_n848), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n759), .A2(new_n516), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n723), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n694), .A2(new_n458), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n849), .A2(new_n766), .A3(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(G169gat), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n934), .A2(new_n935), .A3(new_n582), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n932), .A2(new_n936), .ZN(G1348gat));
  OAI21_X1  g736(.A(G176gat), .B1(new_n934), .B2(new_n725), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n670), .A2(G176gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n930), .B2(new_n939), .ZN(G1349gat));
  AOI211_X1 g739(.A(new_n690), .B(new_n930), .C1(new_n469), .C2(new_n468), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n934), .A2(new_n690), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n942), .A2(new_n234), .ZN(new_n943));
  OR3_X1    g742(.A1(new_n941), .A2(new_n943), .A3(KEYINPUT60), .ZN(new_n944));
  OAI21_X1  g743(.A(KEYINPUT60), .B1(new_n941), .B2(new_n943), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n934), .B2(new_n614), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n947), .A2(KEYINPUT125), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(KEYINPUT125), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(KEYINPUT61), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n931), .A2(new_n224), .A3(new_n691), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n950), .B(new_n951), .C1(KEYINPUT61), .C2(new_n949), .ZN(G1351gat));
  AND4_X1   g751(.A1(new_n424), .A2(new_n928), .A3(new_n508), .A4(new_n850), .ZN(new_n953));
  AOI21_X1  g752(.A(G197gat), .B1(new_n953), .B2(new_n723), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n506), .A2(new_n694), .A3(new_n458), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n916), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n718), .A2(G197gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(G1352gat));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n724), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(G204gat), .ZN(new_n960));
  INV_X1    g759(.A(G204gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n953), .A2(new_n961), .A3(new_n669), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n960), .A2(new_n964), .ZN(G1353gat));
  NAND3_X1  g764(.A1(new_n953), .A2(new_n208), .A3(new_n641), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n916), .A2(new_n641), .A3(new_n955), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n967), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT63), .B1(new_n967), .B2(G211gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(G1354gat));
  AOI21_X1  g769(.A(G218gat), .B1(new_n953), .B2(new_n691), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n691), .A2(G218gat), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT126), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n971), .B1(new_n956), .B2(new_n973), .ZN(G1355gat));
endmodule


