//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1214, new_n1215, new_n1216, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT64), .Z(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n210), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n202), .A2(new_n203), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G50), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n213), .B1(KEYINPUT1), .B2(new_n220), .C1(new_n222), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  XNOR2_X1  g0042(.A(KEYINPUT8), .B(G58), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n208), .A2(G33), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g0045(.A1(G20), .A2(G33), .ZN(new_n246));
  AOI21_X1  g0046(.A(new_n245), .B1(G150), .B2(new_n246), .ZN(new_n247));
  AOI22_X1  g0047(.A1(new_n247), .A2(KEYINPUT67), .B1(G20), .B2(new_n204), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n248), .B1(KEYINPUT67), .B2(new_n247), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G1), .A2(G13), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n252), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n201), .B1(new_n207), .B2(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n255), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n257), .A2(new_n258), .B1(new_n201), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT9), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n263), .B1(new_n221), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n221), .A2(new_n264), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(new_n268), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n272), .A2(G226), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  OR2_X1    g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n277), .A2(G223), .B1(new_n280), .B2(G77), .ZN(new_n281));
  INV_X1    g0081(.A(G222), .ZN(new_n282));
  OR2_X1    g0082(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n283), .B(new_n284), .C1(new_n278), .C2(new_n279), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n281), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  AOI211_X1 g0086(.A(new_n269), .B(new_n273), .C1(new_n286), .C2(new_n271), .ZN(new_n287));
  INV_X1    g0087(.A(G200), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n289), .B1(G190), .B2(new_n287), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n262), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT10), .ZN(new_n292));
  INV_X1    g0092(.A(G179), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n261), .B(new_n294), .C1(G169), .C2(new_n287), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n246), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(new_n201), .ZN(new_n298));
  INV_X1    g0098(.A(G77), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n244), .A2(new_n299), .B1(new_n208), .B2(G68), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n252), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT11), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT69), .B1(new_n255), .B2(G68), .ZN(new_n304));
  XOR2_X1   g0104(.A(new_n304), .B(KEYINPUT12), .Z(new_n305));
  NAND2_X1  g0105(.A1(new_n207), .A2(G20), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n257), .A2(G68), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n301), .A2(new_n302), .ZN(new_n308));
  AND4_X1   g0108(.A1(new_n303), .A2(new_n305), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT14), .ZN(new_n311));
  AND2_X1   g0111(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n312));
  NOR2_X1   g0112(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G226), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G232), .A2(G1698), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n280), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AND3_X1   g0117(.A1(KEYINPUT68), .A2(G33), .A3(G97), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT68), .B1(G33), .B2(G97), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n271), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT13), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n269), .B1(G238), .B2(new_n272), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n322), .B1(new_n321), .B2(new_n323), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n311), .B(G169), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n326), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(G179), .A3(new_n324), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n324), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n311), .B1(new_n331), .B2(G169), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n310), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(G200), .ZN(new_n334));
  INV_X1    g0134(.A(G190), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n334), .B(new_n309), .C1(new_n335), .C2(new_n331), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n243), .A2(new_n297), .B1(new_n208), .B2(new_n299), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT15), .B(G87), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n244), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n252), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n306), .A2(G77), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n341), .B1(G77), .B2(new_n255), .C1(new_n256), .C2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n269), .B1(G244), .B2(new_n272), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n280), .A2(G107), .ZN(new_n345));
  INV_X1    g0145(.A(G232), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n285), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(G238), .B2(new_n277), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n344), .B1(new_n348), .B2(new_n270), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n343), .B1(new_n349), .B2(G200), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n335), .B2(new_n349), .ZN(new_n351));
  INV_X1    g0151(.A(G169), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n353), .B(new_n343), .C1(G179), .C2(new_n349), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  OR3_X1    g0155(.A1(new_n296), .A2(new_n337), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n275), .A2(new_n276), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  NOR3_X1   g0158(.A1(new_n357), .A2(new_n358), .A3(G20), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT7), .B1(new_n280), .B2(new_n208), .ZN(new_n360));
  OAI21_X1  g0160(.A(G68), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  XNOR2_X1  g0161(.A(G58), .B(G68), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(G20), .B1(G159), .B2(new_n246), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT16), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n361), .A2(KEYINPUT16), .A3(new_n363), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(new_n252), .ZN(new_n368));
  XOR2_X1   g0168(.A(KEYINPUT8), .B(G58), .Z(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n306), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n370), .A2(KEYINPUT70), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n256), .B1(new_n370), .B2(KEYINPUT70), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n255), .B2(new_n369), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n368), .A2(new_n375), .A3(KEYINPUT71), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT71), .B1(new_n368), .B2(new_n375), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT18), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n357), .A2(G226), .A3(G1698), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G87), .ZN(new_n381));
  INV_X1    g0181(.A(G223), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n380), .B(new_n381), .C1(new_n382), .C2(new_n285), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n271), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n269), .B1(G232), .B2(new_n272), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G169), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n293), .B2(new_n386), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n378), .A2(new_n379), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n368), .A2(new_n375), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT71), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n254), .B1(new_n364), .B2(new_n365), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n374), .B1(new_n393), .B2(new_n367), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT71), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(new_n395), .A3(new_n388), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT18), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n384), .A2(G190), .A3(new_n385), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n386), .A2(G200), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n368), .A2(new_n375), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n398), .B1(new_n401), .B2(KEYINPUT72), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n400), .A2(new_n399), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT72), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n403), .A2(new_n394), .A3(new_n404), .A4(KEYINPUT17), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n389), .A2(new_n397), .A3(new_n402), .A4(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n356), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n266), .A2(KEYINPUT5), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n207), .A2(G45), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT73), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT5), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G41), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT73), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(new_n207), .A4(G45), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n266), .A2(KEYINPUT5), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n411), .A2(new_n415), .A3(new_n265), .A4(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT74), .ZN(new_n418));
  AND2_X1   g0218(.A1(G33), .A2(G41), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n416), .B(G274), .C1(new_n419), .C2(new_n251), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT74), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(new_n415), .A4(new_n411), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n409), .A2(new_n410), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n271), .B1(new_n425), .B2(new_n416), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G264), .A2(G1698), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n283), .A2(new_n284), .ZN(new_n428));
  INV_X1    g0228(.A(G257), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n357), .B(new_n427), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G303), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n270), .B1(new_n280), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n426), .A2(G270), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n424), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G283), .ZN(new_n435));
  INV_X1    g0235(.A(G97), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n435), .B(new_n208), .C1(G33), .C2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(G116), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G20), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n252), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT20), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n437), .A2(KEYINPUT20), .A3(new_n252), .A4(new_n439), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n207), .A2(G33), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n255), .A2(new_n445), .A3(new_n251), .A4(new_n250), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G116), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n259), .A2(new_n438), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n444), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n434), .A2(G169), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT78), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT21), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n451), .A2(KEYINPUT78), .A3(KEYINPUT21), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n424), .A2(new_n433), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n457), .A2(KEYINPUT77), .A3(G179), .A4(new_n450), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n450), .A2(new_n424), .A3(G179), .A4(new_n433), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT77), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n450), .B1(new_n434), .B2(G200), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(KEYINPUT79), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(KEYINPUT79), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n457), .A2(G190), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n456), .B(new_n462), .C1(new_n464), .C2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n435), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n277), .B2(G250), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT4), .ZN(new_n471));
  OAI21_X1  g0271(.A(G244), .B1(new_n278), .B2(new_n279), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n471), .B1(new_n472), .B2(new_n428), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n357), .A2(new_n314), .A3(KEYINPUT4), .A4(G244), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n470), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n271), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n426), .A2(G257), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n476), .A2(new_n424), .A3(G190), .A4(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT75), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(new_n424), .A3(new_n477), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G200), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n259), .A2(new_n436), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n446), .B2(new_n436), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT6), .ZN(new_n485));
  INV_X1    g0285(.A(G107), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n436), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(G97), .A2(G107), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n486), .A2(KEYINPUT6), .A3(G97), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(G20), .B1(G77), .B2(new_n246), .ZN(new_n492));
  OAI21_X1  g0292(.A(G107), .B1(new_n359), .B2(new_n360), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n484), .B1(new_n494), .B2(new_n252), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n418), .A2(new_n423), .B1(G257), .B2(new_n426), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n496), .A2(KEYINPUT75), .A3(new_n476), .A4(G190), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n480), .A2(new_n482), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(G257), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT83), .ZN(new_n500));
  XNOR2_X1  g0300(.A(new_n499), .B(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G250), .ZN(new_n502));
  INV_X1    g0302(.A(G33), .ZN(new_n503));
  INV_X1    g0303(.A(G294), .ZN(new_n504));
  OAI22_X1  g0304(.A1(new_n285), .A2(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n271), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n426), .A2(G264), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(new_n424), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G200), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT81), .B1(new_n208), .B2(G107), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT23), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT23), .ZN(new_n512));
  OAI211_X1 g0312(.A(KEYINPUT81), .B(new_n512), .C1(new_n208), .C2(G107), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n503), .A2(new_n438), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n511), .A2(new_n513), .B1(new_n208), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n208), .B(G87), .C1(new_n278), .C2(new_n279), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT22), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(KEYINPUT80), .A3(new_n517), .ZN(new_n518));
  XNOR2_X1  g0318(.A(KEYINPUT80), .B(KEYINPUT22), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n357), .A2(new_n519), .A3(new_n208), .A4(G87), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n515), .A2(new_n518), .A3(KEYINPUT24), .A4(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n515), .A2(new_n518), .A3(new_n520), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT24), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n254), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OR3_X1    g0324(.A1(new_n255), .A2(KEYINPUT25), .A3(G107), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT25), .B1(new_n255), .B2(G107), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n525), .B(new_n526), .C1(new_n486), .C2(new_n446), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n527), .A2(KEYINPUT82), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(KEYINPUT82), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n521), .A2(new_n524), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n506), .A2(G190), .A3(new_n424), .A4(new_n507), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n509), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n481), .A2(new_n352), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n494), .A2(new_n252), .ZN(new_n534));
  INV_X1    g0334(.A(new_n484), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n496), .A2(new_n293), .A3(new_n476), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n533), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n498), .A2(new_n532), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n410), .A2(new_n502), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n207), .A2(new_n263), .A3(G45), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n270), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n357), .A2(new_n314), .A3(G238), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n357), .A2(G244), .A3(G1698), .ZN(new_n545));
  INV_X1    g0345(.A(new_n514), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n547), .B2(new_n271), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G190), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n288), .B2(new_n548), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n357), .A2(new_n208), .A3(G68), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT19), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n244), .B2(new_n436), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NOR3_X1   g0354(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT19), .B1(new_n318), .B2(new_n319), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n555), .B1(new_n556), .B2(new_n208), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n252), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n339), .A2(new_n259), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n447), .A2(G87), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n550), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT76), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n548), .A2(new_n352), .ZN(new_n564));
  AOI211_X1 g0364(.A(new_n293), .B(new_n543), .C1(new_n547), .C2(new_n271), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n472), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n514), .B1(new_n567), .B2(G1698), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n270), .B1(new_n568), .B2(new_n544), .ZN(new_n569));
  OAI21_X1  g0369(.A(G169), .B1(new_n569), .B2(new_n543), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n548), .A2(G179), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(KEYINPUT76), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n558), .A2(new_n559), .ZN(new_n574));
  INV_X1    g0374(.A(new_n339), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n447), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n562), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n508), .A2(new_n352), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n524), .A2(new_n521), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n528), .A2(new_n529), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n506), .A2(new_n293), .A3(new_n424), .A4(new_n507), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  NOR4_X1   g0385(.A1(new_n408), .A2(new_n468), .A3(new_n539), .A4(new_n585), .ZN(G372));
  AND2_X1   g0386(.A1(new_n498), .A2(new_n538), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT86), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n570), .A2(new_n571), .B1(new_n574), .B2(new_n576), .ZN(new_n589));
  OAI211_X1 g0389(.A(KEYINPUT84), .B(G200), .C1(new_n569), .C2(new_n543), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT84), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n548), .B2(new_n288), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n592), .A3(new_n549), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n561), .A2(KEYINPUT85), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT85), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n558), .A2(new_n596), .A3(new_n559), .A4(new_n560), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n589), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n587), .A2(new_n588), .A3(new_n532), .A4(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n577), .B1(new_n564), .B2(new_n565), .ZN(new_n601));
  INV_X1    g0401(.A(new_n598), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(new_n593), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT86), .B1(new_n539), .B2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n451), .A2(KEYINPUT78), .A3(KEYINPUT21), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT21), .B1(new_n451), .B2(KEYINPUT78), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n584), .B(new_n462), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT87), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n456), .A2(KEYINPUT87), .A3(new_n462), .A4(new_n584), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n600), .A2(new_n604), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n598), .A2(new_n549), .A3(new_n590), .A4(new_n592), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n533), .A2(new_n536), .A3(new_n537), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT26), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .A4(new_n601), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n601), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n614), .B1(new_n578), .B2(new_n613), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n407), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n402), .A2(new_n405), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n354), .B(KEYINPUT88), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n336), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n621), .B1(new_n624), .B2(new_n333), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n390), .A2(new_n379), .A3(new_n388), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n379), .B1(new_n390), .B2(new_n388), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n292), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n295), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n631), .B(KEYINPUT89), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n620), .A2(new_n632), .ZN(G369));
  NAND2_X1  g0433(.A1(new_n456), .A2(new_n462), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n636), .A2(G213), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G343), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n640), .A2(new_n450), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n468), .B2(new_n641), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n643), .A2(G330), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n532), .B1(new_n530), .B2(new_n639), .ZN(new_n645));
  INV_X1    g0445(.A(new_n584), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n584), .B2(new_n639), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n640), .B1(new_n456), .B2(new_n462), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n651), .A2(new_n647), .B1(new_n646), .B2(new_n639), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(G399));
  INV_X1    g0453(.A(new_n211), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(G41), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n555), .A2(new_n438), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n655), .A2(new_n656), .A3(new_n207), .ZN(new_n657));
  INV_X1    g0457(.A(new_n224), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n657), .B1(new_n658), .B2(new_n655), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT90), .ZN(new_n660));
  XOR2_X1   g0460(.A(new_n660), .B(KEYINPUT28), .Z(new_n661));
  NAND2_X1  g0461(.A1(new_n619), .A2(new_n639), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT91), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT29), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n619), .A2(new_n665), .A3(new_n639), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  OR4_X1    g0467(.A1(new_n468), .A2(new_n585), .A3(new_n539), .A4(new_n640), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n506), .A2(new_n507), .A3(new_n548), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n434), .A2(new_n293), .ZN(new_n670));
  INV_X1    g0470(.A(new_n481), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT30), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n669), .A2(new_n670), .A3(new_n671), .A4(KEYINPUT30), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n548), .A2(G179), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n508), .A2(new_n676), .A3(new_n481), .A4(new_n434), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n674), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n640), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT31), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n678), .A2(KEYINPUT31), .A3(new_n640), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n668), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  INV_X1    g0485(.A(new_n607), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n686), .A2(new_n539), .A3(new_n603), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT26), .B1(new_n603), .B2(new_n538), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n578), .A2(new_n614), .A3(new_n613), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n601), .B(KEYINPUT92), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n639), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT29), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n667), .A2(new_n685), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT93), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n667), .A2(KEYINPUT93), .A3(new_n685), .A4(new_n693), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n661), .B1(new_n698), .B2(G1), .ZN(G364));
  AND2_X1   g0499(.A1(new_n208), .A2(G13), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n207), .B1(new_n700), .B2(G45), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n655), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n654), .A2(new_n280), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G355), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(G116), .B2(new_n211), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n654), .A2(new_n357), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n267), .B2(new_n658), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n241), .A2(G45), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n706), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G13), .A2(G33), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G20), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n251), .B1(G20), .B2(new_n352), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n703), .B1(new_n711), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n288), .A2(G190), .ZN(new_n719));
  OAI21_X1  g0519(.A(G20), .B1(new_n719), .B2(G179), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT95), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n720), .A2(new_n721), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G294), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n208), .A2(new_n293), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G190), .A2(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G311), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n719), .A2(new_n208), .A3(new_n293), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G322), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n280), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n208), .A2(G179), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n729), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n732), .B(new_n736), .C1(G329), .C2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(G190), .A3(G200), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n737), .A2(new_n335), .A3(G200), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n742), .A2(G303), .B1(new_n744), .B2(G283), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n728), .A2(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n335), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(G190), .ZN(new_n748));
  XNOR2_X1  g0548(.A(KEYINPUT33), .B(G317), .ZN(new_n749));
  AOI22_X1  g0549(.A1(G326), .A2(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n727), .A2(new_n740), .A3(new_n745), .A4(new_n750), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT96), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n743), .A2(new_n486), .ZN(new_n753));
  INV_X1    g0553(.A(new_n747), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n357), .B1(new_n202), .B2(new_n734), .C1(new_n754), .C2(new_n201), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n753), .B(new_n755), .C1(G87), .C2(new_n742), .ZN(new_n756));
  INV_X1    g0556(.A(new_n730), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT94), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n757), .A2(KEYINPUT94), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G77), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n726), .A2(G97), .ZN(new_n764));
  INV_X1    g0564(.A(new_n748), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT32), .ZN(new_n766));
  INV_X1    g0566(.A(G159), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n738), .A2(new_n767), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n765), .A2(new_n203), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(new_n766), .B2(new_n768), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n756), .A2(new_n763), .A3(new_n764), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n751), .A2(KEYINPUT96), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n752), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n718), .B1(new_n773), .B2(new_n715), .ZN(new_n774));
  INV_X1    g0574(.A(new_n714), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n774), .B1(new_n643), .B2(new_n775), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT97), .Z(new_n777));
  NOR2_X1   g0577(.A1(new_n643), .A2(G330), .ZN(new_n778));
  INV_X1    g0578(.A(new_n655), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n778), .B(new_n644), .C1(new_n779), .C2(new_n701), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(G396));
  AND2_X1   g0582(.A1(new_n663), .A2(new_n666), .ZN(new_n783));
  INV_X1    g0583(.A(new_n355), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n343), .A2(new_n640), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n622), .B2(new_n785), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n355), .A2(new_n640), .ZN(new_n788));
  AOI21_X1  g0588(.A(KEYINPUT100), .B1(new_n619), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT100), .ZN(new_n790));
  INV_X1    g0590(.A(new_n788), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n790), .B(new_n791), .C1(new_n611), .C2(new_n618), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n783), .A2(new_n787), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n703), .B1(new_n793), .B2(new_n685), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n685), .B2(new_n793), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n715), .A2(new_n712), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT98), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n703), .B1(new_n797), .B2(G77), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n744), .A2(G87), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n765), .A2(new_n800), .B1(new_n741), .B2(new_n486), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n799), .B(new_n801), .C1(G303), .C2(new_n747), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n762), .A2(G116), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n280), .B1(new_n738), .B2(new_n731), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G294), .B2(new_n733), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n802), .A2(new_n764), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n743), .A2(new_n203), .ZN(new_n807));
  INV_X1    g0607(.A(G132), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n357), .B1(new_n738), .B2(new_n808), .C1(new_n201), .C2(new_n741), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n807), .B(new_n809), .C1(new_n726), .C2(G58), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n747), .A2(G137), .B1(G143), .B2(new_n733), .ZN(new_n811));
  INV_X1    g0611(.A(G150), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n811), .B1(new_n812), .B2(new_n765), .C1(new_n761), .C2(new_n767), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n810), .B1(new_n814), .B2(KEYINPUT34), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT34), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n806), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT99), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n715), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n818), .B2(new_n819), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n798), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n713), .B2(new_n787), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n795), .A2(new_n824), .ZN(G384));
  NAND2_X1  g0625(.A1(new_n491), .A2(KEYINPUT35), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n222), .A2(new_n438), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n491), .B2(KEYINPUT35), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT101), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n829), .B2(new_n828), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT36), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n658), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n201), .A2(G68), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n207), .B(G13), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT104), .ZN(new_n837));
  NOR4_X1   g0637(.A1(new_n468), .A2(new_n585), .A3(new_n539), .A4(new_n640), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n681), .A2(new_n682), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n787), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT102), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n330), .A2(new_n332), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n336), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n309), .A2(new_n639), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n844), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n333), .A2(new_n336), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AND4_X1   g0648(.A1(new_n841), .A2(new_n333), .A3(new_n336), .A4(new_n846), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n837), .B1(new_n840), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n392), .A2(new_n395), .A3(new_n638), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n396), .A2(new_n853), .A3(new_n854), .A4(new_n401), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n390), .A2(new_n388), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n401), .ZN(new_n857));
  INV_X1    g0657(.A(new_n638), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n394), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT37), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n379), .B1(new_n378), .B2(new_n388), .ZN(new_n862));
  AND4_X1   g0662(.A1(new_n379), .A2(new_n392), .A3(new_n395), .A4(new_n388), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n862), .A2(new_n863), .A3(new_n621), .ZN(new_n864));
  INV_X1    g0664(.A(new_n859), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(KEYINPUT38), .B(new_n861), .C1(new_n864), .C2(new_n865), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n849), .B1(new_n847), .B2(new_n845), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n684), .A2(new_n871), .A3(KEYINPUT104), .A4(new_n787), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n852), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT40), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n840), .A2(new_n851), .A3(new_n874), .ZN(new_n876));
  AOI221_X4 g0676(.A(new_n867), .B1(new_n855), .B2(new_n860), .C1(new_n406), .C2(new_n859), .ZN(new_n877));
  INV_X1    g0677(.A(new_n853), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n402), .A2(new_n405), .A3(KEYINPUT103), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n628), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT103), .B1(new_n402), .B2(new_n405), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n878), .B2(new_n857), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n855), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT38), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT105), .B1(new_n877), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n885), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT105), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(new_n888), .A3(new_n869), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n876), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n875), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n407), .A3(new_n684), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(G330), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n891), .B1(new_n407), .B2(new_n684), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n667), .A2(new_n693), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n407), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n897), .A2(new_n632), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n877), .B2(new_n885), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n868), .A2(KEYINPUT39), .A3(new_n869), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n333), .A2(new_n640), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n902), .A2(new_n903), .B1(new_n628), .B2(new_n638), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n354), .A2(new_n640), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n789), .B2(new_n792), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n907), .A2(new_n870), .A3(new_n871), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n898), .B(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n895), .A2(KEYINPUT106), .A3(new_n910), .ZN(new_n911));
  OAI221_X1 g0711(.A(new_n911), .B1(new_n207), .B2(new_n700), .C1(new_n910), .C2(new_n895), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT106), .B1(new_n895), .B2(new_n910), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n836), .B1(new_n912), .B2(new_n913), .ZN(G367));
  AOI21_X1  g0714(.A(new_n717), .B1(new_n654), .B2(new_n575), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n707), .A2(new_n233), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n655), .B(new_n702), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n599), .B1(new_n598), .B2(new_n639), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n602), .A2(new_n589), .A3(new_n640), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n743), .A2(new_n299), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n747), .A2(G143), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n765), .B2(new_n767), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n921), .B(new_n923), .C1(G58), .C2(new_n742), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n726), .A2(G68), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n762), .A2(G50), .ZN(new_n926));
  INV_X1    g0726(.A(G137), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n357), .B1(new_n738), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(G150), .B2(new_n733), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n924), .A2(new_n925), .A3(new_n926), .A4(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n743), .A2(new_n436), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(G294), .B2(new_n748), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n731), .B2(new_n754), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(G107), .B2(new_n726), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n739), .A2(G317), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n935), .B(new_n280), .C1(new_n431), .C2(new_n734), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n741), .A2(new_n438), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(KEYINPUT46), .B2(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n934), .B(new_n938), .C1(new_n800), .C2(new_n761), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n937), .A2(KEYINPUT46), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT112), .Z(new_n941));
  OAI21_X1  g0741(.A(new_n930), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT47), .Z(new_n943));
  OAI221_X1 g0743(.A(new_n917), .B1(new_n775), .B2(new_n920), .C1(new_n943), .C2(new_n821), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n701), .B(KEYINPUT111), .Z(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n651), .A2(new_n647), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n649), .B2(new_n651), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(new_n644), .Z(new_n949));
  INV_X1    g0749(.A(KEYINPUT45), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT110), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n536), .A2(new_n640), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n498), .A2(new_n538), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(KEYINPUT108), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n613), .A2(new_n640), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT108), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n498), .A2(new_n956), .A3(new_n538), .A4(new_n952), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n652), .A2(new_n951), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n951), .B1(new_n652), .B2(new_n958), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n950), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n961), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n963), .A2(new_n959), .A3(KEYINPUT45), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT44), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n652), .A2(new_n965), .A3(new_n958), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n965), .B1(new_n652), .B2(new_n958), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n962), .A2(new_n964), .A3(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n650), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n962), .A2(new_n650), .A3(new_n964), .A4(new_n968), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n698), .B1(new_n949), .B2(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n655), .B(KEYINPUT41), .Z(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n946), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n958), .B(KEYINPUT109), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n978), .A2(new_n646), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n639), .B1(new_n979), .B2(new_n613), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n958), .A2(new_n647), .A3(new_n651), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT42), .Z(new_n982));
  INV_X1    g0782(.A(KEYINPUT43), .ZN(new_n983));
  INV_X1    g0783(.A(new_n920), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT107), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n920), .A2(KEYINPUT107), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n980), .A2(new_n982), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n988), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n983), .B2(new_n984), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n980), .B2(new_n982), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n970), .A2(new_n978), .ZN(new_n994));
  OR3_X1    g0794(.A1(new_n990), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n990), .B2(new_n993), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n944), .B1(new_n977), .B2(new_n997), .ZN(G387));
  INV_X1    g0798(.A(new_n949), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n698), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n696), .A2(new_n697), .A3(new_n949), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1000), .A2(new_n655), .A3(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n649), .A2(new_n775), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n704), .A2(new_n656), .B1(new_n486), .B2(new_n654), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n230), .A2(new_n267), .ZN(new_n1005));
  AOI211_X1 g0805(.A(G45), .B(new_n656), .C1(G68), .C2(G77), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT50), .B1(new_n369), .B2(new_n201), .ZN(new_n1007));
  AND3_X1   g0807(.A1(new_n369), .A2(KEYINPUT50), .A3(new_n201), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n707), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1004), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n716), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n703), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n734), .A2(new_n201), .B1(new_n730), .B2(new_n203), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n280), .B(new_n1014), .C1(G150), .C2(new_n739), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n726), .A2(new_n575), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n931), .B1(G159), .B2(new_n747), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n748), .A2(new_n369), .B1(new_n742), .B2(G77), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n357), .B1(new_n739), .B2(G326), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n748), .A2(G311), .B1(G317), .B2(new_n733), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n735), .B2(new_n754), .C1(new_n761), .C2(new_n431), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT48), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n726), .A2(G283), .B1(G294), .B2(new_n742), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT113), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT49), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1020), .B1(new_n438), .B2(new_n743), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1019), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1003), .B(new_n1013), .C1(new_n1032), .C2(new_n715), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n999), .B2(new_n946), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1002), .A2(new_n1034), .ZN(G393));
  NAND2_X1  g0835(.A1(new_n1000), .A2(new_n973), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n949), .B1(new_n696), .B2(new_n697), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n973), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n779), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n946), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n238), .A2(new_n708), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n716), .B1(new_n436), .B2(new_n211), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n703), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n761), .A2(new_n243), .B1(new_n201), .B2(new_n765), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n725), .A2(new_n299), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT114), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n747), .A2(G150), .B1(G159), .B2(new_n733), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT51), .Z(new_n1050));
  AOI211_X1 g0850(.A(new_n280), .B(new_n799), .C1(G143), .C2(new_n739), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n203), .C2(new_n741), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n725), .A2(new_n438), .B1(new_n431), .B2(new_n765), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT115), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n747), .A2(G317), .B1(G311), .B2(new_n733), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT52), .Z(new_n1057));
  NAND2_X1  g0857(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n280), .B1(new_n738), .B2(new_n735), .C1(new_n504), .C2(new_n730), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n753), .B(new_n1059), .C1(G283), .C2(new_n742), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1057), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n1048), .A2(new_n1052), .B1(new_n1055), .B2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT116), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1044), .B1(new_n1063), .B2(new_n715), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n978), .B2(new_n775), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1041), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1040), .A2(new_n1067), .ZN(G390));
  NAND3_X1  g0868(.A1(new_n684), .A2(G330), .A3(new_n787), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(new_n851), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT117), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n619), .A2(new_n788), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n790), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n619), .A2(KEYINPUT100), .A3(new_n788), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n905), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n903), .B1(new_n1076), .B2(new_n851), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n902), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n903), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n787), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n906), .B1(new_n692), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1079), .B1(new_n1081), .B2(new_n871), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1082), .A2(new_n889), .A3(new_n886), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1072), .B1(new_n1078), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1079), .B1(new_n907), .B2(new_n871), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n900), .A2(new_n901), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1072), .B(new_n1083), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1071), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1081), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1069), .A2(new_n851), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1070), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1069), .B(new_n871), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(new_n1076), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n407), .A2(G330), .A3(new_n684), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1094), .A2(new_n632), .A3(new_n897), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1071), .B1(new_n1098), .B2(KEYINPUT117), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1089), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(KEYINPUT117), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1070), .B1(new_n1102), .B2(new_n1087), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1096), .B1(new_n1103), .B2(new_n1099), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1101), .A2(new_n1104), .A3(new_n655), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n807), .B1(G87), .B2(new_n742), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n800), .B2(new_n754), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n280), .B1(new_n738), .B2(new_n504), .C1(new_n734), .C2(new_n438), .ZN(new_n1108));
  OR3_X1    g0908(.A1(new_n1107), .A2(new_n1046), .A3(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n761), .A2(new_n436), .B1(new_n486), .B2(new_n765), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT119), .Z(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT54), .B(G143), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n761), .A2(new_n1112), .B1(new_n927), .B2(new_n765), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT118), .Z(new_n1114));
  INV_X1    g0914(.A(G125), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n357), .B1(new_n738), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(G128), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n754), .A2(new_n1117), .B1(new_n743), .B2(new_n201), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1116), .B(new_n1118), .C1(G132), .C2(new_n733), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n741), .A2(new_n812), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT53), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1119), .B(new_n1121), .C1(new_n767), .C2(new_n725), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1109), .A2(new_n1111), .B1(new_n1114), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT120), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n821), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n1124), .B2(new_n1123), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1126), .B(new_n703), .C1(new_n369), .C2(new_n797), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n902), .B2(new_n712), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1102), .A2(new_n1087), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1099), .B1(new_n1129), .B2(new_n1071), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1128), .B1(new_n1130), .B2(new_n946), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1105), .A2(new_n1131), .ZN(G378));
  NAND3_X1  g0932(.A1(new_n875), .A2(G330), .A3(new_n890), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n296), .A2(new_n261), .A3(new_n638), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n261), .A2(new_n638), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n292), .A2(new_n295), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1134), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1133), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1144), .A2(G330), .A3(new_n875), .A4(new_n890), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n909), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1143), .A2(new_n1145), .A3(new_n909), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1142), .A2(new_n712), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n702), .B(new_n655), .C1(new_n201), .C2(new_n796), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT122), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n734), .A2(new_n486), .B1(new_n339), .B2(new_n730), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n266), .B(new_n280), .C1(new_n738), .C2(new_n800), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n747), .A2(G116), .B1(new_n742), .B2(G77), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n743), .A2(new_n202), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G97), .B2(new_n748), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n925), .A2(new_n1155), .A3(new_n1156), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT58), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(G33), .A2(G41), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT121), .ZN(new_n1162));
  AOI21_X1  g0962(.A(G50), .B1(new_n280), .B2(new_n266), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1159), .A2(new_n1160), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n734), .A2(new_n1117), .B1(new_n730), .B2(new_n927), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G132), .B2(new_n748), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1112), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n747), .A2(G125), .B1(new_n742), .B2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1166), .B(new_n1168), .C1(new_n812), .C2(new_n725), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1162), .B1(G124), .B2(new_n739), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(new_n767), .C2(new_n743), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1164), .B1(new_n1160), .B2(new_n1159), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1152), .B1(new_n1174), .B2(new_n715), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1149), .A2(new_n946), .B1(new_n1150), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n898), .A2(new_n1095), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1101), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT57), .B1(new_n1179), .B2(new_n1149), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1177), .B1(new_n1130), .B2(new_n1097), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1148), .ZN(new_n1182));
  OAI21_X1  g0982(.A(KEYINPUT57), .B1(new_n1182), .B2(new_n1146), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n655), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1176), .B1(new_n1180), .B2(new_n1184), .ZN(G375));
  INV_X1    g0985(.A(new_n1094), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1177), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1187), .A2(new_n976), .A3(new_n1096), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n754), .A2(new_n504), .B1(new_n741), .B2(new_n436), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n921), .B(new_n1189), .C1(G116), .C2(new_n748), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n762), .A2(G107), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n280), .B1(new_n734), .B2(new_n800), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G303), .B2(new_n739), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1190), .A2(new_n1016), .A3(new_n1191), .A4(new_n1193), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n357), .B1(new_n738), .B2(new_n1117), .C1(new_n812), .C2(new_n730), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1157), .B(new_n1195), .C1(G159), .C2(new_n742), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n201), .B2(new_n725), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT123), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n748), .A2(new_n1167), .B1(G137), .B2(new_n733), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n808), .B2(new_n754), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1194), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n715), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1202), .B(new_n703), .C1(G68), .C2(new_n797), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n851), .B2(new_n712), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1094), .B2(new_n946), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1188), .A2(new_n1205), .ZN(G381));
  INV_X1    g1006(.A(G375), .ZN(new_n1207));
  INV_X1    g1007(.A(G378), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(G381), .A2(G387), .A3(G390), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1002), .A2(new_n781), .A3(new_n1034), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(G384), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT124), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .A4(new_n1212), .ZN(G407));
  INV_X1    g1013(.A(G343), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(G213), .ZN(new_n1215));
  OR3_X1    g1015(.A1(G375), .A2(G378), .A3(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(G407), .A2(new_n1216), .A3(G213), .ZN(G409));
  INV_X1    g1017(.A(new_n1210), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n781), .B1(new_n1002), .B2(new_n1034), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1038), .A2(new_n999), .B1(new_n696), .B2(new_n697), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n945), .B1(new_n1221), .B2(new_n975), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n995), .A2(new_n996), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(G390), .A2(new_n1224), .A3(new_n944), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1066), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(G387), .A2(new_n1226), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1220), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1219), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1225), .A2(new_n1227), .B1(new_n1210), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT126), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1228), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1229), .A2(new_n1210), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1220), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT126), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1232), .A2(new_n1237), .ZN(new_n1238));
  OAI211_X1 g1038(.A(G378), .B(new_n1176), .C1(new_n1180), .C2(new_n1184), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1103), .A2(new_n1099), .A3(new_n1096), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1149), .B(new_n976), .C1(new_n1240), .C2(new_n1177), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1176), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1208), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1239), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT62), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1096), .A2(KEYINPUT60), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1187), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n655), .B1(new_n1187), .B2(new_n1246), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1205), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(G384), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(G384), .B(new_n1205), .C1(new_n1247), .C2(new_n1248), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1244), .A2(new_n1245), .A3(new_n1215), .A4(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT61), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1239), .A2(new_n1243), .B1(G213), .B2(new_n1214), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1257));
  INV_X1    g1057(.A(G2897), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1215), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1251), .B(new_n1252), .C1(new_n1258), .C2(new_n1215), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1254), .B(new_n1255), .C1(new_n1256), .C2(new_n1262), .ZN(new_n1263));
  XOR2_X1   g1063(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1256), .B2(new_n1253), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1238), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1244), .A2(new_n1215), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT61), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT63), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n1268), .B2(new_n1257), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1256), .A2(KEYINPUT63), .A3(new_n1253), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1269), .A2(new_n1271), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1266), .A2(new_n1274), .ZN(G405));
  INV_X1    g1075(.A(new_n1239), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1149), .B(KEYINPUT57), .C1(new_n1240), .C2(new_n1177), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1101), .A2(new_n1178), .B1(new_n1148), .B2(new_n1147), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1277), .B(new_n655), .C1(new_n1278), .C2(KEYINPUT57), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G378), .B1(new_n1279), .B2(new_n1176), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1253), .B1(new_n1276), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G375), .A2(new_n1208), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n1257), .A3(new_n1239), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1238), .A3(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT127), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1238), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1281), .A2(new_n1238), .A3(KEYINPUT127), .A4(new_n1283), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1286), .A2(new_n1289), .A3(new_n1290), .ZN(G402));
endmodule


