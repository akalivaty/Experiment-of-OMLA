//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1139, new_n1140, new_n1141;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n457), .A2(G567), .ZN(new_n460));
  INV_X1    g035(.A(G2106), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n470), .A3(G125), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n466), .B1(new_n471), .B2(KEYINPUT68), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(new_n474), .A3(G125), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n464), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n469), .B1(new_n467), .B2(KEYINPUT69), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G137), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n482), .B(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n476), .A2(new_n485), .ZN(G160));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G112), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n464), .B1(new_n477), .B2(new_n479), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(G124), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n480), .A2(G136), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  NOR2_X1   g069(.A1(new_n464), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n490), .B2(G126), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(new_n480), .B2(G138), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n473), .A2(new_n464), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n498), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT71), .B1(new_n506), .B2(G651), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT6), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT72), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(new_n506), .A3(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n511), .A2(new_n515), .A3(G543), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n511), .A2(new_n515), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G88), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(new_n509), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n518), .A2(new_n526), .A3(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  XOR2_X1   g105(.A(KEYINPUT73), .B(KEYINPUT7), .Z(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n517), .A2(G51), .ZN(new_n536));
  XOR2_X1   g111(.A(KEYINPUT74), .B(G89), .Z(new_n537));
  NAND2_X1  g112(.A1(new_n525), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(new_n517), .A2(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n525), .A2(G90), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n509), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  XNOR2_X1  g121(.A(KEYINPUT75), .B(G43), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n517), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n525), .A2(G81), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n509), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  NAND4_X1  g133(.A1(new_n511), .A2(new_n515), .A3(G53), .A4(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n507), .A2(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n561), .A2(new_n562), .A3(G53), .A4(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AND4_X1   g139(.A1(G91), .A2(new_n511), .A3(new_n515), .A4(new_n523), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n568));
  AND2_X1   g143(.A1(KEYINPUT5), .A2(G543), .ZN(new_n569));
  NOR2_X1   g144(.A1(KEYINPUT5), .A2(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n521), .A2(KEYINPUT77), .A3(new_n522), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n567), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n574), .B(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n564), .A2(new_n566), .A3(new_n577), .ZN(G299));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n524), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n580), .B(new_n581), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n523), .A2(G74), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n517), .A2(G49), .B1(G651), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(G288));
  NAND2_X1  g160(.A1(new_n523), .A2(G61), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(KEYINPUT79), .B1(G73), .B2(G543), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n523), .A2(new_n588), .A3(G61), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n509), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(G48), .ZN(new_n591));
  INV_X1    g166(.A(G86), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n591), .A2(new_n516), .B1(new_n524), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G305));
  INV_X1    g170(.A(G47), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n596), .A2(new_n516), .B1(new_n524), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n600), .A2(new_n601), .B1(new_n509), .B2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n525), .A2(G92), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT10), .Z(new_n606));
  NAND2_X1  g181(.A1(new_n571), .A2(new_n572), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n509), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(G54), .B2(new_n517), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n604), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n604), .B1(new_n612), .B2(G868), .ZN(G321));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(G299), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G168), .B2(new_n615), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(G168), .B2(new_n615), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n552), .A2(new_n615), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n611), .A2(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n615), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT81), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND3_X1   g200(.A1(new_n468), .A2(new_n470), .A3(new_n464), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G2104), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n630), .A2(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n480), .A2(G135), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n490), .A2(G123), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n464), .A2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND3_X1  g213(.A1(new_n631), .A2(new_n632), .A3(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT84), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2430), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(G14), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n650), .ZN(G401));
  XOR2_X1   g230(.A(G2067), .B(G2678), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT85), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(G2072), .A2(G2078), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n442), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n657), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(KEYINPUT17), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n657), .A2(new_n664), .A3(new_n658), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n658), .B1(new_n657), .B2(new_n661), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT86), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(new_n657), .B2(new_n664), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n663), .B(new_n665), .C1(new_n668), .C2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n678), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT20), .Z(new_n682));
  AOI211_X1 g257(.A(new_n680), .B(new_n682), .C1(new_n675), .C2(new_n679), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1981), .B(G1986), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT87), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n685), .B(new_n689), .ZN(G229));
  MUX2_X1   g265(.A(G24), .B(G290), .S(G16), .Z(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(G1986), .Z(new_n692));
  OR2_X1    g267(.A1(G95), .A2(G2105), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n693), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT88), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n480), .A2(G131), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n490), .A2(G119), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G25), .B(new_n698), .S(G29), .Z(new_n699));
  XOR2_X1   g274(.A(KEYINPUT35), .B(G1991), .Z(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT89), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G6), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n594), .B2(new_n703), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT90), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT32), .B(G1981), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n703), .A2(G23), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G288), .B2(G16), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT33), .B(G1976), .Z(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n710), .A2(new_n712), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n703), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n703), .ZN(new_n716));
  INV_X1    g291(.A(G1971), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n708), .A2(new_n713), .A3(new_n714), .A4(new_n718), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n692), .B(new_n702), .C1(new_n719), .C2(KEYINPUT34), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(KEYINPUT34), .B2(new_n719), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n637), .A2(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(KEYINPUT95), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(KEYINPUT95), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT31), .B(G11), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT30), .B(G28), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(new_n724), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n726), .A2(new_n727), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n703), .A2(G21), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G168), .B2(new_n703), .ZN(new_n733));
  NOR2_X1   g308(.A1(G5), .A2(G16), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT96), .Z(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G301), .B2(new_n703), .ZN(new_n736));
  INV_X1    g311(.A(G1961), .ZN(new_n737));
  OAI22_X1  g312(.A1(new_n733), .A2(G1966), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n731), .B(new_n738), .C1(G1966), .C2(new_n733), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT97), .ZN(new_n740));
  AND2_X1   g315(.A1(KEYINPUT24), .A2(G34), .ZN(new_n741));
  NOR2_X1   g316(.A1(KEYINPUT24), .A2(G34), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n724), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT93), .Z(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G160), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT94), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2084), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n612), .A2(G16), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G4), .B2(G16), .ZN(new_n749));
  INV_X1    g324(.A(G1348), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n724), .A2(G35), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G162), .B2(new_n724), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT29), .Z(new_n754));
  INV_X1    g329(.A(G2090), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n749), .B2(new_n750), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n740), .A2(new_n747), .A3(new_n751), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n724), .A2(G32), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT26), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n467), .A2(G2105), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n762), .A2(new_n763), .B1(G105), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n490), .A2(G129), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n480), .A2(G141), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n759), .B1(new_n770), .B2(new_n724), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT27), .B(G1996), .Z(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT25), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G139), .B2(new_n480), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n464), .B2(new_n778), .ZN(new_n779));
  MUX2_X1   g354(.A(G33), .B(new_n779), .S(G29), .Z(new_n780));
  OAI21_X1  g355(.A(new_n774), .B1(G2072), .B2(new_n780), .ZN(new_n781));
  AOI211_X1 g356(.A(new_n773), .B(new_n781), .C1(G2072), .C2(new_n780), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n553), .A2(new_n703), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n703), .B2(G19), .ZN(new_n784));
  INV_X1    g359(.A(G1341), .ZN(new_n785));
  NAND2_X1  g360(.A1(G164), .A2(G29), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G27), .B2(G29), .ZN(new_n787));
  INV_X1    g362(.A(G2078), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n784), .A2(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n754), .A2(new_n755), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n724), .A2(G26), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n490), .A2(G128), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT91), .Z(new_n795));
  OAI21_X1  g370(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n796));
  INV_X1    g371(.A(G116), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G2105), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n480), .B2(G140), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n793), .B1(new_n800), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2067), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n782), .A2(new_n789), .A3(new_n790), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n784), .A2(new_n785), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n737), .B2(new_n736), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n703), .A2(G20), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT23), .ZN(new_n807));
  INV_X1    g382(.A(G299), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(new_n703), .ZN(new_n809));
  INV_X1    g384(.A(G1956), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n805), .B(new_n811), .C1(new_n788), .C2(new_n787), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n758), .A2(new_n803), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n723), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT98), .ZN(G311));
  INV_X1    g390(.A(KEYINPUT99), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n814), .B(new_n816), .ZN(G150));
  NAND2_X1  g392(.A1(new_n612), .A2(G559), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT38), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n517), .A2(G55), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n525), .A2(G93), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n820), .B(new_n821), .C1(new_n509), .C2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n553), .B(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n819), .B(new_n824), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n826), .A2(new_n827), .A3(G860), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n823), .A2(G860), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT37), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n828), .A2(new_n830), .ZN(G145));
  XNOR2_X1  g406(.A(new_n800), .B(new_n504), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n698), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n490), .A2(G130), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT101), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n835), .A2(new_n464), .A3(G118), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n464), .B2(G118), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n837), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n834), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G142), .B2(new_n480), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n629), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n779), .B(new_n769), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n833), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(G162), .B(new_n637), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT100), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(G160), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n844), .B(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(KEYINPUT102), .B(G37), .Z(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g426(.A1(new_n823), .A2(new_n615), .ZN(new_n852));
  XNOR2_X1  g427(.A(G288), .B(KEYINPUT103), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n594), .ZN(new_n854));
  XNOR2_X1  g429(.A(G290), .B(G166), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT42), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n611), .B(new_n808), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT41), .Z(new_n859));
  XOR2_X1   g434(.A(new_n622), .B(new_n824), .Z(new_n860));
  MUX2_X1   g435(.A(new_n858), .B(new_n859), .S(new_n860), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n857), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n852), .B1(new_n862), .B2(new_n615), .ZN(G295));
  OAI21_X1  g438(.A(new_n852), .B1(new_n862), .B2(new_n615), .ZN(G331));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n824), .B(G301), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G168), .ZN(new_n867));
  INV_X1    g442(.A(new_n858), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n859), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n856), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n869), .A2(new_n856), .A3(new_n870), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(new_n849), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT43), .ZN(new_n876));
  AOI21_X1  g451(.A(G37), .B1(new_n871), .B2(new_n872), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT43), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(new_n878), .A3(new_n874), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n865), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  AND4_X1   g455(.A1(new_n878), .A2(new_n873), .A3(new_n849), .A4(new_n874), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n878), .B1(new_n877), .B2(new_n874), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n880), .B1(new_n865), .B2(new_n883), .ZN(G397));
  INV_X1    g459(.A(KEYINPUT113), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT57), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n560), .A2(new_n563), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n576), .B1(new_n607), .B2(G65), .ZN(new_n890));
  INV_X1    g465(.A(G91), .ZN(new_n891));
  OAI22_X1  g466(.A1(new_n890), .A2(new_n509), .B1(new_n891), .B2(new_n524), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n888), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(KEYINPUT113), .A2(KEYINPUT57), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT114), .Z(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  NAND3_X1  g472(.A1(G299), .A2(new_n888), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G1384), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n478), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT3), .B1(new_n478), .B2(G2104), .ZN(new_n902));
  OAI211_X1 g477(.A(G138), .B(new_n464), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  AOI22_X1  g478(.A1(new_n903), .A2(KEYINPUT4), .B1(new_n626), .B2(new_n502), .ZN(new_n904));
  OAI21_X1  g479(.A(G2105), .B1(new_n901), .B2(new_n902), .ZN(new_n905));
  INV_X1    g480(.A(G126), .ZN(new_n906));
  OAI22_X1  g481(.A1(new_n905), .A2(new_n906), .B1(new_n495), .B2(new_n496), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n900), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT50), .ZN(new_n909));
  XOR2_X1   g484(.A(KEYINPUT104), .B(G40), .Z(new_n910));
  NOR3_X1   g485(.A1(new_n476), .A2(new_n485), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT50), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n504), .A2(new_n913), .A3(new_n900), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n810), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n908), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n900), .ZN(new_n919));
  XNOR2_X1  g494(.A(KEYINPUT56), .B(G2072), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n918), .A2(new_n919), .A3(new_n911), .A4(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n899), .A2(new_n916), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT115), .B1(new_n912), .B2(new_n915), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT115), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n909), .A2(new_n924), .A3(new_n911), .A4(new_n914), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n750), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT116), .ZN(new_n927));
  INV_X1    g502(.A(G2067), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n626), .A2(new_n502), .ZN(new_n929));
  AOI211_X1 g504(.A(new_n501), .B(G2105), .C1(new_n477), .C2(new_n479), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n929), .B1(new_n930), .B2(new_n499), .ZN(new_n931));
  AOI21_X1  g506(.A(G1384), .B1(new_n931), .B2(new_n498), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n911), .A2(new_n928), .A3(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n926), .A2(new_n927), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n927), .B1(new_n926), .B2(new_n933), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n934), .A2(new_n935), .A3(new_n611), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n569), .A2(new_n570), .A3(new_n568), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT77), .B1(new_n521), .B2(new_n522), .ZN(new_n938));
  OAI21_X1  g513(.A(G65), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n576), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n565), .B1(new_n941), .B2(G651), .ZN(new_n942));
  AOI211_X1 g517(.A(new_n887), .B(new_n895), .C1(new_n942), .C2(new_n564), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n897), .B1(G299), .B2(new_n888), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n471), .A2(KEYINPUT68), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(new_n475), .A3(new_n465), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(G2105), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n481), .A2(new_n484), .ZN(new_n949));
  INV_X1    g524(.A(new_n910), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(KEYINPUT50), .B2(new_n908), .ZN(new_n952));
  AOI21_X1  g527(.A(G1956), .B1(new_n952), .B2(new_n914), .ZN(new_n953));
  INV_X1    g528(.A(new_n921), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n945), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n922), .B1(new_n936), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT119), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n958), .A2(KEYINPUT61), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n955), .A2(new_n922), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(KEYINPUT61), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n955), .A2(new_n922), .A3(new_n958), .A4(KEYINPUT61), .ZN(new_n963));
  XNOR2_X1  g538(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n964));
  INV_X1    g539(.A(G1996), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n918), .A2(new_n965), .A3(new_n919), .A4(new_n911), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n911), .A2(new_n932), .ZN(new_n967));
  XOR2_X1   g542(.A(KEYINPUT58), .B(G1341), .Z(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT117), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n553), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n966), .A2(new_n969), .A3(KEYINPUT117), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n964), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT117), .B1(new_n966), .B2(new_n969), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n976), .A2(new_n552), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT59), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(KEYINPUT118), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n977), .B(new_n979), .C1(new_n971), .C2(new_n970), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n962), .A2(new_n963), .A3(new_n975), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT120), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n974), .A2(new_n976), .A3(new_n552), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n960), .A2(new_n961), .B1(new_n983), .B2(new_n979), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT120), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n984), .A2(new_n985), .A3(new_n963), .A4(new_n975), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT60), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT60), .B1(new_n934), .B2(new_n935), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n612), .ZN(new_n990));
  OAI211_X1 g565(.A(KEYINPUT60), .B(new_n611), .C1(new_n934), .C2(new_n935), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n957), .B1(new_n987), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G2084), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n952), .A2(new_n994), .A3(new_n914), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT111), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n918), .A2(new_n919), .A3(new_n911), .ZN(new_n997));
  INV_X1    g572(.A(G1966), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n952), .A2(new_n1000), .A3(new_n994), .A4(new_n914), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n996), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G8), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT121), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n996), .A2(G168), .A3(new_n999), .A4(new_n1001), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(G8), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1002), .A2(G286), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1004), .B(KEYINPUT51), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT121), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n1002), .B2(G8), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n1011));
  OAI211_X1 g586(.A(G8), .B(new_n1005), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT107), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n911), .B1(new_n932), .B2(KEYINPUT45), .ZN(new_n1015));
  INV_X1    g590(.A(new_n919), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n918), .A2(KEYINPUT107), .A3(new_n919), .A4(new_n911), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(new_n717), .A3(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n952), .A2(new_n755), .A3(new_n914), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT108), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G303), .A2(G8), .ZN(new_n1024));
  XOR2_X1   g599(.A(KEYINPUT109), .B(KEYINPUT55), .Z(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(KEYINPUT109), .A2(KEYINPUT55), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1026), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1019), .A2(KEYINPUT108), .A3(new_n1020), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1023), .A2(G8), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1021), .A2(G8), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n1028), .ZN(new_n1033));
  INV_X1    g608(.A(G1976), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT52), .B1(G288), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n582), .A2(G1976), .A3(new_n584), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n967), .A2(new_n1037), .A3(G8), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1037), .B1(new_n967), .B2(G8), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1035), .B(new_n1036), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n587), .A2(new_n589), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G651), .ZN(new_n1043));
  INV_X1    g618(.A(new_n593), .ZN(new_n1044));
  INV_X1    g619(.A(G1981), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n1047));
  OAI21_X1  g622(.A(G1981), .B1(new_n590), .B2(new_n593), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1047), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1050));
  OAI22_X1  g625(.A1(new_n1039), .A2(new_n1040), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1041), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1040), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1038), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1053), .B1(new_n1055), .B2(new_n1036), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1031), .A2(new_n1033), .A3(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(G301), .B(KEYINPUT54), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(G2078), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT122), .B(G1961), .Z(new_n1063));
  NAND3_X1  g638(.A1(new_n923), .A2(new_n925), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n788), .A2(KEYINPUT53), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1062), .B(new_n1064), .C1(new_n997), .C2(new_n1065), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n918), .A2(G40), .A3(G160), .ZN(new_n1068));
  XOR2_X1   g643(.A(new_n1068), .B(KEYINPUT124), .Z(new_n1069));
  NOR2_X1   g644(.A1(new_n1016), .A2(new_n1065), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1059), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1059), .A2(new_n1066), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1013), .A2(new_n1058), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n993), .A2(new_n1073), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1031), .A2(new_n1057), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1002), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1023), .A2(G8), .A3(new_n1030), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1076), .B1(new_n1077), .B2(new_n1028), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1002), .A2(G8), .A3(G168), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1031), .A2(new_n1033), .A3(new_n1057), .A4(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT63), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT112), .ZN(new_n1085));
  OR3_X1    g660(.A1(new_n1031), .A2(new_n1056), .A3(new_n1052), .ZN(new_n1086));
  AND4_X1   g661(.A1(new_n1034), .A2(new_n1051), .A3(new_n582), .A4(new_n584), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1046), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1055), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .A4(new_n1089), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1075), .A2(new_n1078), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT112), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1013), .A2(KEYINPUT62), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT62), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1008), .A2(new_n1095), .A3(new_n1012), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1066), .A2(G171), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1094), .A2(new_n1058), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1074), .A2(new_n1090), .A3(new_n1093), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n918), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n911), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(G1996), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n770), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1103), .B(KEYINPUT105), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1101), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n800), .A2(G2067), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n795), .A2(new_n928), .A3(new_n799), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n965), .B2(new_n770), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1104), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n698), .B(new_n700), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT106), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1110), .B1(new_n1101), .B2(new_n1112), .ZN(new_n1113));
  OR2_X1    g688(.A1(G290), .A2(G1986), .ZN(new_n1114));
  NAND2_X1  g689(.A1(G290), .A2(G1986), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1101), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1099), .A2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1102), .A2(KEYINPUT46), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1101), .B1(new_n1108), .B2(new_n770), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1102), .A2(KEYINPUT46), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  XOR2_X1   g697(.A(new_n1122), .B(KEYINPUT47), .Z(new_n1123));
  NOR2_X1   g698(.A1(new_n1114), .A2(new_n1101), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT125), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT48), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1123), .B1(new_n1113), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n700), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n698), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1110), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1101), .B1(new_n1130), .B2(new_n1107), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1118), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1118), .A2(KEYINPUT126), .A3(new_n1132), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g712(.A1(G229), .A2(G227), .A3(G401), .A4(new_n462), .ZN(new_n1139));
  XOR2_X1   g713(.A(new_n1139), .B(KEYINPUT127), .Z(new_n1140));
  NAND2_X1  g714(.A1(new_n1140), .A2(new_n850), .ZN(new_n1141));
  NOR2_X1   g715(.A1(new_n1141), .A2(new_n883), .ZN(G308));
  OR2_X1    g716(.A1(new_n1141), .A2(new_n883), .ZN(G225));
endmodule


