//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G353));
  NOR2_X1   g0006(.A1(G97), .A2(G107), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  AND2_X1   g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G20), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n202), .A2(new_n203), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n213), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n216), .B1(new_n218), .B2(new_n220), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n233), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n201), .A2(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n203), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n242), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(KEYINPUT67), .ZN(new_n249));
  AND2_X1   g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G1), .A2(G13), .ZN(new_n251));
  OAI21_X1  g0051(.A(G274), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G274), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n255), .B1(new_n217), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(KEYINPUT67), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n250), .A2(new_n251), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n260), .ZN(new_n264));
  INV_X1    g0064(.A(G226), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT68), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n265), .A2(KEYINPUT68), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  OR2_X1    g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n273), .A2(G223), .B1(new_n276), .B2(G77), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n271), .A2(new_n272), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G222), .A3(new_n270), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n263), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n269), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G179), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n211), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G150), .ZN(new_n288));
  OR2_X1    g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(G20), .B2(new_n204), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n251), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n296), .A2(new_n251), .A3(new_n292), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(G50), .C1(G1), .C2(new_n211), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(G50), .B2(new_n296), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n282), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n285), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  XOR2_X1   g0103(.A(new_n303), .B(KEYINPUT69), .Z(new_n304));
  INV_X1    g0104(.A(KEYINPUT9), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n283), .A2(G190), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n282), .A2(G200), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n295), .A2(new_n299), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT9), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n306), .A2(new_n307), .A3(new_n308), .A4(new_n310), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n311), .A2(KEYINPUT10), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(KEYINPUT10), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n289), .A2(KEYINPUT70), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n289), .A2(KEYINPUT70), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n316), .A2(new_n286), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT15), .B(G87), .ZN(new_n319));
  INV_X1    g0119(.A(G77), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n319), .A2(new_n287), .B1(new_n211), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n293), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n296), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n320), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n297), .B(G77), .C1(G1), .C2(new_n211), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n273), .A2(G238), .B1(new_n276), .B2(G107), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n235), .B1(new_n271), .B2(new_n272), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n270), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n263), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n254), .A2(new_n261), .B1(new_n264), .B2(G244), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n327), .B1(new_n301), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n334), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n284), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n326), .B1(new_n334), .B2(G200), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(KEYINPUT71), .B1(G190), .B2(new_n336), .ZN(new_n340));
  INV_X1    g0140(.A(G200), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n327), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT71), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  AND4_X1   g0145(.A1(new_n304), .A2(new_n314), .A3(new_n338), .A4(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT13), .ZN(new_n347));
  OAI211_X1 g0147(.A(G226), .B(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT72), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n278), .A2(KEYINPUT72), .A3(G226), .A4(new_n270), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n329), .A2(G1698), .B1(G33), .B2(G97), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n263), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n264), .A2(G238), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n262), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n347), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n217), .A2(new_n256), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n352), .B2(new_n353), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n361), .A2(new_n357), .A3(KEYINPUT13), .ZN(new_n362));
  OAI21_X1  g0162(.A(G169), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT14), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n355), .A2(new_n358), .A3(new_n347), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT13), .B1(new_n361), .B2(new_n357), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(G179), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n366), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT14), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n369), .A3(G169), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n364), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n287), .A2(new_n320), .B1(new_n211), .B2(G68), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT73), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n372), .A2(new_n373), .B1(new_n201), .B2(new_n289), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n372), .A2(new_n373), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n293), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT11), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OR3_X1    g0178(.A1(new_n296), .A2(KEYINPUT12), .A3(G68), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT12), .B1(new_n296), .B2(G68), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n203), .B1(new_n210), .B2(G20), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n379), .A2(new_n380), .B1(new_n297), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n376), .B2(new_n377), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n371), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(G200), .B1(new_n359), .B2(new_n362), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n365), .A2(G190), .A3(new_n366), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G223), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n270), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n265), .A2(G1698), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n392), .B(new_n393), .C1(new_n274), .C2(new_n275), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G33), .A2(G87), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(new_n263), .B1(new_n264), .B2(G232), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT76), .ZN(new_n398));
  INV_X1    g0198(.A(G190), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .A4(new_n262), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n396), .A2(new_n263), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n264), .A2(G232), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n262), .A2(new_n402), .A3(new_n399), .A4(new_n403), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n404), .A2(KEYINPUT76), .ZN(new_n405));
  NOR2_X1   g0205(.A1(G223), .A2(G1698), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n265), .B2(G1698), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(new_n278), .B1(G33), .B2(G87), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n403), .B1(new_n408), .B2(new_n360), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n254), .A2(new_n261), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n341), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n401), .B1(new_n405), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT77), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n286), .B1(new_n210), .B2(G20), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n297), .B1(new_n323), .B2(new_n286), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G58), .A2(G68), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT75), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(KEYINPUT75), .A2(G58), .A3(G68), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n219), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n289), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n421), .A2(G20), .B1(G159), .B2(new_n422), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n274), .A2(new_n275), .A3(G20), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT7), .ZN(new_n425));
  OAI21_X1  g0225(.A(G68), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n271), .A2(new_n211), .A3(new_n272), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n423), .B(KEYINPUT16), .C1(new_n426), .C2(new_n430), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n431), .A2(new_n293), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT16), .ZN(new_n433));
  INV_X1    g0233(.A(new_n423), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n429), .A2(new_n427), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n272), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n203), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n433), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n416), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT17), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n431), .A2(new_n293), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n435), .A2(new_n436), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G68), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT16), .B1(new_n443), .B2(new_n423), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n415), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(G169), .B1(new_n409), .B2(new_n410), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n397), .A2(G179), .A3(new_n262), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT18), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n413), .A2(KEYINPUT17), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n413), .A2(KEYINPUT17), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n404), .A2(KEYINPUT76), .ZN(new_n453));
  AOI21_X1  g0253(.A(G200), .B1(new_n397), .B2(new_n262), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n400), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n451), .B(new_n452), .C1(new_n455), .C2(new_n445), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT18), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n445), .A2(new_n448), .A3(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n440), .A2(new_n450), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n346), .A2(new_n390), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n210), .A2(G45), .ZN(new_n463));
  OR2_X1    g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  NAND2_X1  g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(new_n263), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n467), .A2(G270), .B1(new_n257), .B2(new_n466), .ZN(new_n468));
  OAI211_X1 g0268(.A(G257), .B(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n271), .A2(G303), .A3(new_n272), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT82), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n273), .A2(new_n472), .A3(G264), .ZN(new_n473));
  OAI211_X1 g0273(.A(G264), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT82), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n471), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n468), .B1(new_n476), .B2(new_n360), .ZN(new_n477));
  INV_X1    g0277(.A(G13), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(G1), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G116), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G20), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G283), .ZN(new_n484));
  INV_X1    g0284(.A(G97), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n484), .B(new_n211), .C1(G33), .C2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(new_n293), .A3(new_n482), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT20), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n486), .A2(KEYINPUT20), .A3(new_n293), .A4(new_n482), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n483), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n210), .A2(G33), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n297), .A2(KEYINPUT83), .A3(G116), .A4(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT83), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n296), .A2(new_n492), .A3(new_n251), .A4(new_n292), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(new_n481), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n477), .A2(new_n498), .A3(G169), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT21), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n469), .A2(new_n470), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n472), .B1(new_n273), .B2(G264), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n474), .A2(KEYINPUT82), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n263), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n498), .A2(new_n506), .A3(G179), .A4(new_n468), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n477), .A2(new_n498), .A3(KEYINPUT21), .A4(G169), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n501), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n477), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G190), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n498), .B1(new_n477), .B2(G200), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n211), .B(G87), .C1(new_n274), .C2(new_n275), .ZN(new_n514));
  OR2_X1    g0314(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n517), .B(KEYINPUT85), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT85), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n517), .B(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(new_n514), .A3(new_n515), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  OR3_X1    g0323(.A1(new_n211), .A2(KEYINPUT23), .A3(G107), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n211), .A2(G33), .A3(G116), .ZN(new_n525));
  NAND2_X1  g0325(.A1(KEYINPUT86), .A2(KEYINPUT24), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n524), .A2(new_n525), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT86), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n523), .A2(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n531), .ZN(new_n533));
  AOI211_X1 g0333(.A(new_n533), .B(new_n528), .C1(new_n519), .C2(new_n522), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n293), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT87), .ZN(new_n536));
  OR2_X1    g0336(.A1(new_n536), .A2(KEYINPUT25), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n211), .A2(G107), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(KEYINPUT25), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n537), .A2(new_n479), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n479), .A2(new_n538), .ZN(new_n541));
  INV_X1    g0341(.A(G107), .ZN(new_n542));
  OAI221_X1 g0342(.A(new_n540), .B1(new_n541), .B2(new_n539), .C1(new_n542), .C2(new_n495), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n535), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(G257), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n546));
  OAI211_X1 g0346(.A(G250), .B(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G294), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n263), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n467), .A2(G264), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n466), .A2(new_n257), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT88), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT88), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n550), .A2(new_n551), .A3(new_n555), .A4(new_n552), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(G169), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n553), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G179), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n545), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(G190), .B1(new_n554), .B2(new_n556), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n558), .A2(G200), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n535), .B(new_n544), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(G244), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n566));
  OAI211_X1 g0366(.A(G238), .B(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G116), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n263), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n463), .A2(G250), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n259), .A2(G1), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n360), .A2(new_n571), .B1(new_n257), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT80), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n570), .A2(KEYINPUT80), .A3(new_n573), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n284), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n278), .A2(new_n211), .A3(G68), .ZN(new_n579));
  NAND3_X1  g0379(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n211), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n208), .B2(G87), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT19), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n287), .B2(new_n485), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n579), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n585), .A2(new_n293), .B1(new_n323), .B2(new_n319), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n319), .B2(new_n495), .ZN(new_n587));
  INV_X1    g0387(.A(new_n577), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT80), .B1(new_n570), .B2(new_n573), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n578), .B(new_n587), .C1(new_n590), .C2(G169), .ZN(new_n591));
  OAI211_X1 g0391(.A(G244), .B(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT4), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .A4(new_n270), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n484), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n263), .ZN(new_n598));
  INV_X1    g0398(.A(new_n465), .ZN(new_n599));
  NOR2_X1   g0399(.A1(KEYINPUT5), .A2(G41), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n572), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n601), .A2(G257), .A3(new_n360), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n552), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT79), .B1(new_n605), .B2(G179), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n603), .B1(new_n597), .B2(new_n263), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT79), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(new_n608), .A3(new_n284), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n605), .A2(new_n301), .ZN(new_n610));
  AND2_X1   g0410(.A1(G97), .A2(G107), .ZN(new_n611));
  OAI22_X1  g0411(.A1(new_n611), .A2(new_n207), .B1(KEYINPUT78), .B2(KEYINPUT6), .ZN(new_n612));
  NOR2_X1   g0412(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(KEYINPUT6), .B2(new_n485), .ZN(new_n614));
  XNOR2_X1  g0414(.A(G97), .B(G107), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n612), .B(G20), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n422), .A2(G77), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n542), .B1(new_n435), .B2(new_n436), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n293), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  MUX2_X1   g0420(.A(new_n296), .B(new_n495), .S(G97), .Z(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n606), .A2(new_n609), .A3(new_n610), .A4(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(G200), .B1(new_n588), .B2(new_n589), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n576), .A2(G190), .A3(new_n577), .ZN(new_n625));
  INV_X1    g0425(.A(G87), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n495), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT81), .ZN(new_n628));
  XNOR2_X1  g0428(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n586), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n624), .A2(new_n625), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n605), .A2(G200), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n607), .A2(G190), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n633), .A2(new_n620), .A3(new_n621), .A4(new_n634), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n591), .A2(new_n623), .A3(new_n632), .A4(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n462), .A2(new_n513), .A3(new_n565), .A4(new_n636), .ZN(new_n637));
  XOR2_X1   g0437(.A(new_n637), .B(KEYINPUT89), .Z(G372));
  NAND2_X1  g0438(.A1(new_n450), .A2(new_n458), .ZN(new_n639));
  INV_X1    g0439(.A(new_n338), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n389), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n386), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n440), .A2(new_n456), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n314), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n304), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT91), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(KEYINPUT91), .B(new_n304), .C1(new_n644), .C2(new_n645), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n622), .B1(G169), .B2(new_n607), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n607), .A2(new_n608), .A3(new_n284), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n608), .B1(new_n607), .B2(new_n284), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n574), .A2(new_n301), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n578), .A2(new_n587), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n574), .A2(G200), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n625), .A2(new_n631), .A3(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n654), .A2(new_n655), .A3(new_n657), .A4(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n660), .A2(new_n657), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n591), .A2(new_n632), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT26), .B1(new_n662), .B2(new_n623), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n535), .A2(new_n544), .B1(new_n557), .B2(new_n559), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT90), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n301), .B1(new_n506), .B2(new_n468), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT21), .B1(new_n666), .B2(new_n498), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n508), .A2(new_n507), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n501), .A2(KEYINPUT90), .A3(new_n507), .A4(new_n508), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n664), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n659), .A2(new_n657), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n672), .A2(new_n564), .A3(new_n623), .A4(new_n635), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n661), .B(new_n663), .C1(new_n671), .C2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n650), .B1(new_n461), .B2(new_n675), .ZN(G369));
  NOR2_X1   g0476(.A1(new_n667), .A2(new_n668), .ZN(new_n677));
  OR3_X1    g0477(.A1(new_n480), .A2(KEYINPUT27), .A3(G20), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT27), .B1(new_n480), .B2(G20), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n565), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n682), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n664), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT92), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT92), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n684), .A2(new_n689), .A3(new_n686), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G330), .ZN(new_n692));
  INV_X1    g0492(.A(new_n498), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n513), .B1(new_n693), .B2(new_n685), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n669), .A2(new_n498), .A3(new_n670), .A4(new_n682), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n692), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n545), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n565), .B1(new_n697), .B2(new_n685), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n561), .B2(new_n685), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n691), .A2(new_n700), .ZN(G399));
  INV_X1    g0501(.A(new_n214), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G41), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G1), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n220), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n659), .A2(new_n657), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT26), .B1(new_n709), .B2(new_n623), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n654), .A2(new_n655), .A3(new_n591), .A4(new_n632), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n710), .A2(new_n711), .A3(new_n657), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n564), .A2(new_n623), .A3(new_n635), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT93), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n677), .A2(new_n561), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT93), .B1(new_n664), .B2(new_n509), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n713), .A2(new_n715), .A3(new_n716), .A4(new_n672), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n682), .B1(new_n712), .B2(new_n717), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n718), .A2(KEYINPUT94), .A3(KEYINPUT29), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT29), .B1(new_n674), .B2(new_n685), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT94), .B1(new_n718), .B2(KEYINPUT29), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n510), .A2(G179), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n550), .A2(new_n551), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n576), .A2(new_n607), .A3(new_n726), .A4(new_n577), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n607), .A2(new_n726), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n477), .A2(new_n284), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n729), .A2(new_n590), .A3(new_n730), .A4(KEYINPUT30), .ZN(new_n731));
  AOI21_X1  g0531(.A(G179), .B1(new_n570), .B2(new_n573), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n605), .A2(new_n477), .A3(new_n553), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n728), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT31), .B1(new_n734), .B2(new_n682), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n636), .A2(new_n565), .A3(new_n513), .A4(new_n685), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n692), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n723), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n708), .B1(new_n743), .B2(G1), .ZN(G364));
  OR2_X1    g0544(.A1(new_n696), .A2(KEYINPUT95), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n478), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n210), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n703), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n696), .A2(KEYINPUT95), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n694), .A2(new_n692), .A3(new_n695), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n745), .A2(new_n750), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n251), .B1(G20), .B2(new_n301), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n211), .A2(new_n284), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n399), .A2(new_n341), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G326), .ZN(new_n760));
  INV_X1    g0560(.A(new_n756), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n761), .A2(new_n399), .A3(G200), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G322), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n760), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G190), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n756), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n278), .B(new_n765), .C1(G311), .C2(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n399), .A2(G179), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n211), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G294), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n341), .A2(G190), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n756), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(KEYINPUT33), .B(G317), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n775), .B1(new_n776), .B2(KEYINPUT99), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(KEYINPUT99), .B2(new_n776), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n211), .A2(G179), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n757), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G303), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n779), .A2(new_n766), .ZN(new_n782));
  INV_X1    g0582(.A(G329), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n780), .A2(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n774), .A2(new_n779), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n784), .B1(G283), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n769), .A2(new_n773), .A3(new_n778), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n771), .A2(new_n485), .ZN(new_n789));
  INV_X1    g0589(.A(new_n775), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(G68), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT98), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n780), .A2(new_n626), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n758), .A2(new_n201), .B1(new_n767), .B2(new_n320), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n793), .B(new_n794), .C1(G58), .C2(new_n762), .ZN(new_n795));
  XOR2_X1   g0595(.A(KEYINPUT97), .B(G159), .Z(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n782), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT32), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n278), .B1(new_n542), .B2(new_n785), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(new_n798), .B2(new_n797), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n792), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n755), .B1(new_n788), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n754), .ZN(new_n806));
  INV_X1    g0606(.A(new_n220), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n278), .B(new_n702), .C1(new_n259), .C2(new_n807), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n247), .A2(new_n259), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n214), .A2(new_n278), .ZN(new_n810));
  INV_X1    g0610(.A(G355), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n810), .A2(new_n811), .B1(G116), .B2(new_n214), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n808), .A2(new_n809), .B1(KEYINPUT96), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(KEYINPUT96), .B2(new_n812), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n750), .B(new_n802), .C1(new_n806), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n694), .A2(new_n695), .ZN(new_n816));
  INV_X1    g0616(.A(new_n805), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n753), .A2(new_n818), .ZN(G396));
  NOR2_X1   g0619(.A1(new_n338), .A2(new_n682), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n326), .A2(new_n682), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n345), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n820), .B1(new_n822), .B2(new_n338), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n675), .B2(new_n682), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n673), .A2(new_n671), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n663), .A2(new_n660), .A3(new_n657), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n823), .B(new_n685), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n749), .B1(new_n829), .B2(new_n741), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n741), .B2(new_n829), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n754), .A2(new_n803), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT100), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n750), .B1(new_n834), .B2(new_n320), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G137), .A2(new_n759), .B1(new_n790), .B2(G150), .ZN(new_n836));
  XNOR2_X1  g0636(.A(KEYINPUT102), .B(G143), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n836), .B1(new_n767), .B2(new_n796), .C1(new_n763), .C2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT34), .ZN(new_n839));
  INV_X1    g0639(.A(new_n780), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G50), .A2(new_n840), .B1(new_n786), .B2(G68), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n202), .B2(new_n771), .ZN(new_n842));
  INV_X1    g0642(.A(new_n782), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n276), .B1(new_n843), .B2(G132), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n844), .A2(KEYINPUT103), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(KEYINPUT103), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n842), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G303), .A2(new_n759), .B1(new_n790), .B2(G283), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n481), .B2(new_n767), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT101), .Z(new_n850));
  AOI22_X1  g0650(.A1(new_n762), .A2(G294), .B1(G311), .B2(new_n843), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n542), .B2(new_n780), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n276), .B1(new_n785), .B2(new_n626), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n852), .A2(new_n789), .A3(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n839), .A2(new_n847), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n835), .B1(new_n755), .B2(new_n855), .C1(new_n823), .C2(new_n804), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n831), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  NOR2_X1   g0658(.A1(new_n746), .A2(new_n210), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n203), .B1(new_n429), .B2(KEYINPUT7), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n429), .B2(new_n428), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT16), .B1(new_n861), .B2(new_n423), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n415), .B1(new_n441), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n680), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n411), .A2(KEYINPUT76), .A3(new_n404), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n438), .A2(new_n293), .A3(new_n431), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n867), .A2(new_n868), .A3(new_n415), .A4(new_n400), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n863), .A2(new_n448), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(new_n870), .A3(new_n865), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT37), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n445), .A2(new_n864), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n869), .A2(new_n449), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n459), .A2(new_n866), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT105), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n459), .A2(new_n866), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n872), .A2(new_n875), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT105), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n459), .A2(new_n445), .A3(new_n864), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n869), .A2(new_n449), .A3(new_n873), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n875), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n878), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n389), .A2(new_n364), .A3(new_n367), .A4(new_n370), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n384), .A2(new_n685), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT104), .ZN(new_n892));
  INV_X1    g0692(.A(new_n890), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n386), .A2(new_n389), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT104), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n889), .A2(new_n895), .A3(new_n890), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n892), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT106), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n735), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n737), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n734), .A2(KEYINPUT106), .A3(KEYINPUT31), .A4(new_n682), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n739), .A2(new_n899), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n897), .A2(new_n902), .A3(new_n823), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT40), .B1(new_n888), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n897), .A2(new_n902), .A3(new_n823), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n876), .A2(KEYINPUT38), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT40), .B1(new_n906), .B2(new_n881), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n462), .A2(new_n902), .ZN(new_n910));
  OAI21_X1  g0710(.A(G330), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n911), .A2(KEYINPUT107), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n909), .A2(new_n910), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(KEYINPUT107), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n820), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n828), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n906), .A2(new_n881), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n917), .A2(new_n918), .A3(new_n897), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n639), .A2(new_n680), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n922), .B(new_n878), .C1(new_n882), .C2(new_n887), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n371), .A2(new_n385), .A3(new_n685), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n906), .A2(KEYINPUT39), .A3(new_n881), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n921), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n718), .A2(KEYINPUT94), .A3(KEYINPUT29), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n718), .A2(KEYINPUT29), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT94), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n929), .B1(new_n932), .B2(new_n720), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n462), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n650), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n928), .B(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n859), .B1(new_n915), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n936), .B2(new_n915), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n218), .A2(new_n481), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT35), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n941), .B2(new_n940), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT36), .Z(new_n944));
  NAND4_X1  g0744(.A1(new_n807), .A2(G77), .A3(new_n419), .A4(new_n420), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n243), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(G1), .A3(new_n478), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n938), .A2(new_n944), .A3(new_n947), .ZN(G367));
  NAND2_X1  g0748(.A1(new_n630), .A2(new_n682), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT108), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n950), .A2(new_n578), .A3(new_n587), .A4(new_n656), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT109), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n951), .B(KEYINPUT109), .C1(new_n709), .C2(new_n950), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n805), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n702), .A2(new_n278), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n232), .ZN(new_n957));
  INV_X1    g0757(.A(new_n806), .ZN(new_n958));
  INV_X1    g0758(.A(new_n319), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n958), .B1(new_n702), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n750), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n786), .A2(G77), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n775), .B2(new_n796), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n276), .B(new_n963), .C1(G58), .C2(new_n840), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n767), .A2(new_n201), .ZN(new_n965));
  INV_X1    g0765(.A(G137), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n758), .A2(new_n837), .B1(new_n782), .B2(new_n966), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n965), .B(new_n967), .C1(G150), .C2(new_n762), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n964), .B(new_n968), .C1(new_n203), .C2(new_n771), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n278), .B1(new_n790), .B2(G294), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n772), .A2(G107), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n840), .A2(KEYINPUT46), .A3(G116), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT46), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n780), .B2(new_n481), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n970), .A2(new_n971), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n762), .A2(G303), .B1(new_n759), .B2(G311), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(KEYINPUT115), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(KEYINPUT115), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n786), .A2(G97), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G283), .A2(new_n768), .B1(new_n843), .B2(G317), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n977), .A2(new_n978), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n969), .B1(new_n975), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT47), .Z(new_n983));
  OAI211_X1 g0783(.A(new_n955), .B(new_n961), .C1(new_n755), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(KEYINPUT113), .A2(KEYINPUT44), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT110), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n654), .A2(new_n986), .A3(new_n682), .ZN(new_n987));
  OAI21_X1  g0787(.A(KEYINPUT110), .B1(new_n623), .B2(new_n685), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n623), .A2(new_n635), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n685), .B1(new_n620), .B2(new_n621), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n987), .A2(new_n988), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n688), .A2(new_n690), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(KEYINPUT113), .A2(KEYINPUT44), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n985), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n994), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n684), .A2(new_n689), .A3(new_n686), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n689), .B1(new_n684), .B2(new_n686), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n996), .B1(new_n999), .B2(new_n992), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n987), .A2(new_n988), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n989), .A2(new_n991), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT45), .B1(new_n691), .B2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(KEYINPUT45), .B(new_n1003), .C1(new_n997), .C2(new_n998), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n995), .A2(new_n1000), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n700), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n999), .A2(new_n992), .A3(new_n996), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n993), .A2(new_n994), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1010), .A2(new_n1011), .A3(new_n985), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT45), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n999), .B2(new_n992), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n1005), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(new_n1015), .A3(new_n700), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1009), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n684), .B1(new_n699), .B2(new_n683), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n745), .A2(new_n751), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT114), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n696), .B(new_n684), .C1(new_n699), .C2(new_n683), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n745), .A2(new_n1018), .A3(KEYINPUT114), .A4(new_n751), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n743), .B1(new_n1017), .B2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n703), .B(KEYINPUT41), .Z(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n748), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT42), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1003), .A2(new_n1029), .A3(new_n565), .A4(new_n683), .ZN(new_n1030));
  OAI21_X1  g0830(.A(KEYINPUT42), .B1(new_n992), .B2(new_n684), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1003), .A2(new_n664), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n682), .B1(new_n1033), .B2(new_n623), .ZN(new_n1034));
  OAI21_X1  g0834(.A(KEYINPUT111), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n992), .A2(new_n561), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n685), .B1(new_n1036), .B2(new_n654), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT111), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1037), .A2(new_n1038), .A3(new_n1031), .A4(new_n1030), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT43), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n954), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1035), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n952), .A2(new_n953), .A3(KEYINPUT43), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1035), .A2(new_n1039), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT112), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(KEYINPUT112), .B1(new_n1050), .B2(new_n1042), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1047), .A2(new_n1051), .B1(new_n700), .B2(new_n992), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1046), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1050), .A2(KEYINPUT112), .A3(new_n1042), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n700), .A2(new_n992), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n984), .B1(new_n1028), .B2(new_n1057), .ZN(G387));
  INV_X1    g0858(.A(new_n1024), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n704), .B1(new_n1059), .B2(new_n743), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n743), .B2(new_n1059), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n699), .A2(new_n817), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n810), .A2(new_n705), .B1(G107), .B2(new_n214), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n705), .ZN(new_n1064));
  AOI211_X1 g0864(.A(G45), .B(new_n1064), .C1(G68), .C2(G77), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n286), .A2(G50), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT50), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n702), .B(new_n278), .C1(new_n1065), .C2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n238), .A2(G45), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1063), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n749), .B1(new_n1070), .B2(new_n958), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT116), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n780), .A2(new_n320), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n979), .A2(new_n278), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(G68), .C2(new_n768), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n759), .A2(G159), .B1(new_n843), .B2(G150), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n775), .A2(new_n286), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n762), .B2(G50), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n772), .A2(new_n959), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n278), .B1(new_n843), .B2(G326), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n762), .A2(G317), .B1(G303), .B2(new_n768), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G322), .A2(new_n759), .B1(new_n790), .B2(G311), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT117), .Z(new_n1085));
  INV_X1    g0885(.A(KEYINPUT48), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n772), .A2(G283), .B1(new_n840), .B2(G294), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT49), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1081), .B1(new_n481), .B2(new_n785), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1080), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1072), .B1(new_n1094), .B2(new_n754), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1059), .A2(new_n748), .B1(new_n1062), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1061), .A2(new_n1096), .ZN(G393));
  INV_X1    g0897(.A(new_n1016), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n700), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n1098), .A2(new_n1099), .B1(new_n742), .B2(new_n1024), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1059), .A2(new_n743), .A3(new_n1009), .A4(new_n1016), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1100), .A2(new_n1101), .A3(new_n703), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n992), .A2(new_n805), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n806), .B1(new_n485), .B2(new_n214), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n956), .B2(new_n242), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n762), .A2(G311), .B1(new_n759), .B2(G317), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT52), .Z(new_n1108));
  INV_X1    g0908(.A(G294), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n276), .B1(new_n785), .B2(new_n542), .C1(new_n1109), .C2(new_n767), .ZN(new_n1110));
  INV_X1    g0910(.A(G283), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n780), .A2(new_n1111), .B1(new_n782), .B2(new_n764), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1110), .B1(KEYINPUT118), .B2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1108), .B(new_n1113), .C1(KEYINPUT118), .C2(new_n1112), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n771), .A2(new_n481), .B1(new_n775), .B2(new_n781), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT119), .Z(new_n1116));
  AOI22_X1  g0916(.A1(new_n762), .A2(G159), .B1(new_n759), .B2(G150), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT51), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n771), .A2(new_n320), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1120), .B(new_n278), .C1(new_n626), .C2(new_n785), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n203), .A2(new_n780), .B1(new_n767), .B2(new_n286), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n775), .A2(new_n201), .B1(new_n782), .B2(new_n837), .ZN(new_n1123));
  OR3_X1    g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1114), .A2(new_n1116), .B1(new_n1118), .B2(new_n1124), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n750), .B(new_n1106), .C1(new_n1125), .C2(new_n754), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1103), .A2(new_n748), .B1(new_n1104), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1102), .A2(new_n1127), .ZN(G390));
  AOI22_X1  g0928(.A1(new_n340), .A2(new_n344), .B1(new_n326), .B2(new_n682), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n916), .B(G330), .C1(new_n640), .C2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n897), .A2(new_n902), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n917), .A2(new_n897), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1133), .A2(new_n924), .B1(new_n923), .B2(new_n926), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n924), .B(new_n878), .C1(new_n882), .C2(new_n887), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n822), .A2(new_n338), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n718), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n916), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1135), .B1(new_n1138), .B2(new_n897), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1132), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  AND4_X1   g0940(.A1(new_n877), .A2(new_n879), .A3(KEYINPUT38), .A4(new_n880), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n887), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n877), .B1(new_n876), .B2(KEYINPUT38), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n820), .B1(new_n718), .B2(new_n1136), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n897), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1144), .B(new_n924), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1130), .B1(new_n738), .B2(new_n739), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n897), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n923), .A2(new_n926), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n925), .B1(new_n917), .B2(new_n897), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1147), .B(new_n1149), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1140), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n748), .ZN(new_n1154));
  INV_X1    g0954(.A(G128), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n780), .A2(new_n288), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT53), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n278), .B1(new_n1155), .B2(new_n758), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G50), .A2(new_n786), .B1(new_n843), .B2(G125), .ZN(new_n1159));
  INV_X1    g0959(.A(G132), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1159), .B1(new_n1160), .B2(new_n763), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1158), .B(new_n1161), .C1(new_n1157), .C2(new_n1156), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT54), .B(G143), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n966), .A2(new_n775), .B1(new_n767), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G159), .B2(new_n772), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT121), .Z(new_n1166));
  NAND2_X1  g0966(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n758), .A2(new_n1111), .B1(new_n785), .B2(new_n203), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1168), .A2(new_n278), .A3(new_n793), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n762), .A2(G116), .B1(G294), .B2(new_n843), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G97), .A2(new_n768), .B1(new_n790), .B2(G107), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1169), .A2(new_n1120), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n755), .B1(new_n1167), .B2(new_n1172), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n750), .B(new_n1173), .C1(new_n286), .C2(new_n834), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n1150), .B2(new_n804), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1154), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n462), .A2(G330), .A3(new_n902), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n650), .B(new_n1177), .C1(new_n723), .C2(new_n461), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1148), .A2(new_n897), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n917), .B1(new_n1132), .B2(new_n1179), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n902), .A2(new_n1131), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1149), .B(new_n1145), .C1(new_n1181), .C2(new_n897), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1178), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1184), .A2(KEYINPUT120), .A3(new_n1152), .A4(new_n1140), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT120), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1140), .A2(new_n1152), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1188), .A2(new_n934), .A3(new_n650), .A4(new_n1177), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1186), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1185), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n704), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1176), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(G378));
  AOI21_X1  g0994(.A(new_n750), .B1(new_n834), .B2(new_n201), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n763), .A2(new_n1155), .B1(new_n775), .B2(new_n1160), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G125), .A2(new_n759), .B1(new_n768), .B2(G137), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n780), .B2(new_n1163), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1196), .B(new_n1198), .C1(G150), .C2(new_n772), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT59), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n843), .A2(G124), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n796), .A2(new_n785), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1204), .A2(G33), .A3(G41), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n762), .A2(G107), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT122), .Z(new_n1208));
  OAI22_X1  g1008(.A1(new_n775), .A2(new_n485), .B1(new_n782), .B2(new_n1111), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n771), .A2(new_n203), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n276), .A2(new_n258), .ZN(new_n1211));
  NOR4_X1   g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1073), .A4(new_n1211), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n767), .A2(new_n319), .B1(new_n785), .B2(new_n202), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G116), .B2(new_n759), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1208), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT58), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1211), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1219));
  AND4_X1   g1019(.A1(new_n1206), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n314), .A2(new_n303), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n309), .A2(new_n680), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1222), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n314), .A2(new_n303), .A3(new_n1224), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1223), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1226), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1224), .B1(new_n314), .B2(new_n303), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n303), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1230), .B(new_n1222), .C1(new_n312), .C2(new_n313), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1228), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1227), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1195), .B1(new_n755), .B2(new_n1220), .C1(new_n1234), .C2(new_n804), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT123), .Z(new_n1236));
  AOI211_X1 g1036(.A(new_n692), .B(new_n1233), .C1(new_n904), .C2(new_n908), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1234), .B1(new_n909), .B2(G330), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1237), .A2(new_n1238), .A3(new_n928), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n921), .A2(new_n927), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n909), .A2(G330), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1233), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n909), .A2(new_n1234), .A3(G330), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1240), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1239), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1236), .B1(new_n1245), .B2(new_n748), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1178), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT120), .B1(new_n1153), .B2(new_n1184), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1187), .A2(new_n1189), .A3(new_n1186), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1247), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT57), .B1(new_n1250), .B2(new_n1245), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1178), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1252));
  OAI21_X1  g1052(.A(KEYINPUT57), .B1(new_n1239), .B2(new_n1244), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n703), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1246), .B1(new_n1251), .B2(new_n1254), .ZN(G375));
  NAND2_X1  g1055(.A1(new_n1146), .A2(new_n803), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n749), .B1(new_n833), .B2(G68), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n762), .A2(G137), .B1(G150), .B2(new_n768), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1258), .B1(new_n1160), .B2(new_n758), .C1(new_n775), .C2(new_n1163), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(G159), .A2(new_n840), .B1(new_n843), .B2(G128), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n276), .B1(new_n786), .B2(G58), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1260), .B(new_n1261), .C1(new_n201), .C2(new_n771), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G116), .A2(new_n790), .B1(new_n843), .B2(G303), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1263), .B1(new_n542), .B2(new_n767), .C1(new_n1111), .C2(new_n763), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(G294), .A2(new_n759), .B1(new_n840), .B2(G97), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1265), .A2(new_n276), .A3(new_n962), .A4(new_n1079), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n1259), .A2(new_n1262), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1257), .B1(new_n1267), .B2(new_n754), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1188), .A2(new_n748), .B1(new_n1256), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1189), .A2(new_n1027), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1178), .A2(new_n1183), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(G381));
  INV_X1    g1072(.A(G396), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1061), .A2(new_n1273), .A3(new_n1096), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(G390), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n1276), .A3(new_n857), .ZN(new_n1277));
  NOR4_X1   g1077(.A1(new_n1277), .A2(G378), .A3(G387), .A4(G381), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1278), .B(new_n1246), .C1(new_n1251), .C2(new_n1254), .ZN(G407));
  NAND2_X1  g1079(.A1(new_n681), .A2(G213), .ZN(new_n1280));
  OR3_X1    g1080(.A1(G375), .A2(G378), .A3(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(G407), .A2(G213), .A3(new_n1281), .ZN(G409));
  NAND2_X1  g1082(.A1(G387), .A2(new_n1276), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1273), .B1(new_n1061), .B2(new_n1096), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1275), .A2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G390), .B(new_n984), .C1(new_n1028), .C2(new_n1057), .ZN(new_n1286));
  AND4_X1   g1086(.A1(KEYINPUT124), .A2(new_n1283), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT124), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1289), .A2(new_n1285), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G378), .B(new_n1246), .C1(new_n1251), .C2(new_n1254), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1239), .A2(new_n1244), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1252), .A2(new_n1294), .A3(new_n1026), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1236), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1294), .B2(new_n747), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1193), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1293), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1271), .B1(KEYINPUT60), .B2(new_n1189), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1178), .A2(new_n1183), .A3(KEYINPUT60), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n703), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1269), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1303));
  OR2_X1    g1103(.A1(new_n1303), .A2(new_n857), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n857), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1299), .A2(new_n1280), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(KEYINPUT62), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n681), .A2(G213), .A3(G2897), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1306), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1304), .A2(new_n1305), .A3(new_n1310), .ZN(new_n1313));
  AND2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1299), .A2(new_n1280), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT61), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1309), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1308), .A2(KEYINPUT62), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1292), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  AOI22_X1  g1120(.A1(new_n1293), .A2(new_n1298), .B1(G213), .B2(new_n681), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1321), .A2(KEYINPUT63), .A3(new_n1307), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT63), .B1(new_n1321), .B2(new_n1307), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n1291), .B(new_n1317), .C1(new_n1325), .C2(new_n1321), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT125), .B1(new_n1324), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT63), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1308), .A2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1321), .A2(KEYINPUT63), .A3(new_n1307), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT125), .ZN(new_n1333));
  NOR3_X1   g1133(.A1(new_n1332), .A2(new_n1333), .A3(new_n1326), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1320), .B1(new_n1328), .B2(new_n1334), .ZN(G405));
  INV_X1    g1135(.A(KEYINPUT127), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1336), .B1(new_n1306), .B2(KEYINPUT126), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1337), .B1(new_n1336), .B2(new_n1306), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(G375), .A2(new_n1193), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1293), .ZN(new_n1340));
  MUX2_X1   g1140(.A(new_n1338), .B(new_n1337), .S(new_n1340), .Z(new_n1341));
  XNOR2_X1  g1141(.A(new_n1341), .B(new_n1292), .ZN(G402));
endmodule


