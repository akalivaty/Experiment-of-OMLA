

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589;

  XNOR2_X2 U324 ( .A(n378), .B(n377), .ZN(n471) );
  XNOR2_X1 U325 ( .A(n317), .B(n316), .ZN(n319) );
  XOR2_X1 U326 ( .A(n350), .B(n349), .Z(n292) );
  NOR2_X1 U327 ( .A1(n573), .A2(n552), .ZN(n399) );
  XOR2_X1 U328 ( .A(G99GAT), .B(G85GAT), .Z(n363) );
  XNOR2_X1 U329 ( .A(n315), .B(KEYINPUT19), .ZN(n316) );
  XNOR2_X1 U330 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n405) );
  NOR2_X1 U331 ( .A1(n470), .A2(n469), .ZN(n487) );
  NOR2_X1 U332 ( .A1(n461), .A2(n572), .ZN(n444) );
  XNOR2_X1 U333 ( .A(n406), .B(n405), .ZN(n529) );
  XNOR2_X1 U334 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U335 ( .A(n360), .B(n388), .Z(n579) );
  NOR2_X1 U336 ( .A1(n571), .A2(n458), .ZN(n548) );
  XNOR2_X1 U337 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U338 ( .A(n329), .B(n328), .Z(n533) );
  XNOR2_X1 U339 ( .A(KEYINPUT38), .B(n492), .ZN(n500) );
  XNOR2_X1 U340 ( .A(n446), .B(KEYINPUT120), .ZN(n447) );
  XNOR2_X1 U341 ( .A(n448), .B(n447), .ZN(G1348GAT) );
  XOR2_X1 U342 ( .A(G29GAT), .B(G43GAT), .Z(n294) );
  XNOR2_X1 U343 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n294), .B(n293), .ZN(n367) );
  XOR2_X1 U345 ( .A(G15GAT), .B(G1GAT), .Z(n389) );
  XOR2_X1 U346 ( .A(n367), .B(n389), .Z(n296) );
  NAND2_X1 U347 ( .A1(G229GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U349 ( .A(G8GAT), .B(KEYINPUT67), .Z(n298) );
  XNOR2_X1 U350 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U352 ( .A(n300), .B(n299), .Z(n308) );
  XOR2_X1 U353 ( .A(G113GAT), .B(G36GAT), .Z(n302) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(G50GAT), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U356 ( .A(KEYINPUT30), .B(G141GAT), .Z(n304) );
  XNOR2_X1 U357 ( .A(G22GAT), .B(G197GAT), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U360 ( .A(n308), .B(n307), .Z(n534) );
  INV_X1 U361 ( .A(n534), .ZN(n573) );
  NAND2_X1 U362 ( .A1(G227GAT), .A2(G233GAT), .ZN(n314) );
  XOR2_X1 U363 ( .A(KEYINPUT78), .B(G99GAT), .Z(n310) );
  XNOR2_X1 U364 ( .A(G43GAT), .B(G15GAT), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n312) );
  XOR2_X1 U366 ( .A(G190GAT), .B(G134GAT), .Z(n311) );
  XNOR2_X1 U367 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n329) );
  XNOR2_X1 U369 ( .A(KEYINPUT80), .B(KEYINPUT17), .ZN(n317) );
  INV_X1 U370 ( .A(KEYINPUT79), .ZN(n315) );
  XNOR2_X1 U371 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n408) );
  XNOR2_X1 U373 ( .A(n408), .B(G71GAT), .ZN(n327) );
  XOR2_X1 U374 ( .A(G120GAT), .B(G127GAT), .Z(n321) );
  XNOR2_X1 U375 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n428) );
  XOR2_X1 U377 ( .A(G183GAT), .B(n428), .Z(n325) );
  XOR2_X1 U378 ( .A(G176GAT), .B(KEYINPUT81), .Z(n323) );
  XNOR2_X1 U379 ( .A(KEYINPUT20), .B(KEYINPUT82), .ZN(n322) );
  XOR2_X1 U380 ( .A(n323), .B(n322), .Z(n324) );
  INV_X1 U381 ( .A(n533), .ZN(n455) );
  XOR2_X1 U382 ( .A(G78GAT), .B(G204GAT), .Z(n335) );
  XOR2_X1 U383 ( .A(KEYINPUT84), .B(KEYINPUT24), .Z(n331) );
  XNOR2_X1 U384 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n333) );
  XNOR2_X1 U386 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n332), .B(KEYINPUT2), .ZN(n432) );
  XNOR2_X1 U388 ( .A(n333), .B(n432), .ZN(n334) );
  XNOR2_X1 U389 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U390 ( .A(G106GAT), .B(G148GAT), .Z(n355) );
  XOR2_X1 U391 ( .A(G22GAT), .B(G155GAT), .Z(n381) );
  XOR2_X1 U392 ( .A(n355), .B(n381), .Z(n337) );
  NAND2_X1 U393 ( .A1(G228GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U395 ( .A(n339), .B(n338), .Z(n344) );
  XOR2_X1 U396 ( .A(KEYINPUT83), .B(G218GAT), .Z(n341) );
  XNOR2_X1 U397 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U399 ( .A(G197GAT), .B(n342), .Z(n407) );
  XOR2_X1 U400 ( .A(G50GAT), .B(G162GAT), .Z(n366) );
  XNOR2_X1 U401 ( .A(n407), .B(n366), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n461) );
  XNOR2_X1 U403 ( .A(KEYINPUT32), .B(n363), .ZN(n346) );
  AND2_X1 U404 ( .A1(G230GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U406 ( .A(KEYINPUT70), .B(KEYINPUT33), .Z(n348) );
  XNOR2_X1 U407 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n348), .B(n347), .ZN(n349) );
  INV_X1 U409 ( .A(G204GAT), .ZN(n354) );
  XOR2_X1 U410 ( .A(KEYINPUT71), .B(G64GAT), .Z(n352) );
  XNOR2_X1 U411 ( .A(G176GAT), .B(G92GAT), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n414) );
  XNOR2_X1 U414 ( .A(n355), .B(n414), .ZN(n356) );
  XNOR2_X1 U415 ( .A(n292), .B(n356), .ZN(n360) );
  XOR2_X1 U416 ( .A(KEYINPUT13), .B(KEYINPUT69), .Z(n358) );
  XNOR2_X1 U417 ( .A(G71GAT), .B(G78GAT), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U419 ( .A(G57GAT), .B(n359), .Z(n388) );
  XOR2_X1 U420 ( .A(KEYINPUT11), .B(KEYINPUT73), .Z(n362) );
  XNOR2_X1 U421 ( .A(KEYINPUT10), .B(KEYINPUT9), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n378) );
  XOR2_X1 U423 ( .A(KEYINPUT65), .B(n363), .Z(n365) );
  XOR2_X1 U424 ( .A(G36GAT), .B(G190GAT), .Z(n410) );
  XNOR2_X1 U425 ( .A(G218GAT), .B(n410), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n367), .B(n366), .ZN(n369) );
  AND2_X1 U428 ( .A1(G232GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U430 ( .A(n371), .B(n370), .Z(n376) );
  XOR2_X1 U431 ( .A(G134GAT), .B(KEYINPUT74), .Z(n431) );
  XOR2_X1 U432 ( .A(G92GAT), .B(KEYINPUT66), .Z(n373) );
  XNOR2_X1 U433 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n431), .B(n374), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U437 ( .A(KEYINPUT36), .B(n471), .ZN(n486) );
  XOR2_X1 U438 ( .A(KEYINPUT76), .B(G64GAT), .Z(n380) );
  XNOR2_X1 U439 ( .A(G127GAT), .B(G211GAT), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n393) );
  XOR2_X1 U441 ( .A(G8GAT), .B(G183GAT), .Z(n409) );
  XOR2_X1 U442 ( .A(n381), .B(n409), .Z(n383) );
  NAND2_X1 U443 ( .A1(G231GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U444 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U445 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n385) );
  XNOR2_X1 U446 ( .A(KEYINPUT77), .B(KEYINPUT12), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U448 ( .A(n387), .B(n386), .Z(n391) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n472) );
  INV_X1 U452 ( .A(n472), .ZN(n585) );
  NOR2_X1 U453 ( .A1(n486), .A2(n585), .ZN(n395) );
  XOR2_X1 U454 ( .A(KEYINPUT45), .B(KEYINPUT112), .Z(n394) );
  XOR2_X1 U455 ( .A(n395), .B(n394), .Z(n396) );
  NAND2_X1 U456 ( .A1(n573), .A2(n396), .ZN(n397) );
  NOR2_X1 U457 ( .A1(n579), .A2(n397), .ZN(n398) );
  XOR2_X1 U458 ( .A(KEYINPUT113), .B(n398), .Z(n404) );
  XOR2_X1 U459 ( .A(KEYINPUT111), .B(n585), .Z(n563) );
  NAND2_X1 U460 ( .A1(n563), .A2(n471), .ZN(n401) );
  XNOR2_X1 U461 ( .A(KEYINPUT41), .B(n579), .ZN(n552) );
  XNOR2_X1 U462 ( .A(n399), .B(KEYINPUT46), .ZN(n400) );
  NOR2_X1 U463 ( .A1(n401), .A2(n400), .ZN(n402) );
  XOR2_X1 U464 ( .A(KEYINPUT47), .B(n402), .Z(n403) );
  NOR2_X1 U465 ( .A1(n404), .A2(n403), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n418) );
  XOR2_X1 U467 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n412) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U470 ( .A(n414), .B(n413), .Z(n416) );
  NAND2_X1 U471 ( .A1(G226GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n518) );
  NOR2_X1 U474 ( .A1(n529), .A2(n518), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n419), .B(KEYINPUT54), .ZN(n441) );
  XOR2_X1 U476 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n421) );
  XNOR2_X1 U477 ( .A(KEYINPUT85), .B(KEYINPUT6), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n440) );
  XOR2_X1 U479 ( .A(G85GAT), .B(G148GAT), .Z(n423) );
  XNOR2_X1 U480 ( .A(G1GAT), .B(G155GAT), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U482 ( .A(KEYINPUT4), .B(KEYINPUT88), .Z(n425) );
  XNOR2_X1 U483 ( .A(G57GAT), .B(KEYINPUT86), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U485 ( .A(n427), .B(n426), .Z(n438) );
  XOR2_X1 U486 ( .A(n428), .B(KEYINPUT87), .Z(n430) );
  NAND2_X1 U487 ( .A1(G225GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n436) );
  XOR2_X1 U489 ( .A(n431), .B(G162GAT), .Z(n434) );
  XNOR2_X1 U490 ( .A(G29GAT), .B(n432), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n468) );
  INV_X1 U495 ( .A(n468), .ZN(n530) );
  NAND2_X1 U496 ( .A1(n441), .A2(n530), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n442), .B(KEYINPUT64), .ZN(n572) );
  XNOR2_X1 U498 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n445) );
  NAND2_X1 U500 ( .A1(n455), .A2(n445), .ZN(n567) );
  NOR2_X1 U501 ( .A1(n573), .A2(n567), .ZN(n448) );
  INV_X1 U502 ( .A(G169GAT), .ZN(n446) );
  XOR2_X1 U503 ( .A(n518), .B(KEYINPUT91), .Z(n449) );
  XNOR2_X1 U504 ( .A(KEYINPUT27), .B(n449), .ZN(n458) );
  XOR2_X1 U505 ( .A(n461), .B(KEYINPUT28), .Z(n525) );
  INV_X1 U506 ( .A(n525), .ZN(n450) );
  NOR2_X1 U507 ( .A1(n458), .A2(n450), .ZN(n531) );
  NAND2_X1 U508 ( .A1(n531), .A2(KEYINPUT92), .ZN(n451) );
  NOR2_X1 U509 ( .A1(n530), .A2(n451), .ZN(n453) );
  NOR2_X1 U510 ( .A1(n531), .A2(KEYINPUT92), .ZN(n452) );
  NOR2_X1 U511 ( .A1(n453), .A2(n452), .ZN(n454) );
  NOR2_X1 U512 ( .A1(n455), .A2(n454), .ZN(n470) );
  NOR2_X1 U513 ( .A1(n455), .A2(KEYINPUT92), .ZN(n466) );
  XOR2_X1 U514 ( .A(KEYINPUT93), .B(KEYINPUT26), .Z(n457) );
  NAND2_X1 U515 ( .A1(n461), .A2(n533), .ZN(n456) );
  XNOR2_X1 U516 ( .A(n457), .B(n456), .ZN(n571) );
  INV_X1 U517 ( .A(KEYINPUT94), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n548), .B(n459), .ZN(n464) );
  NOR2_X1 U519 ( .A1(n518), .A2(n533), .ZN(n460) );
  NOR2_X1 U520 ( .A1(n461), .A2(n460), .ZN(n462) );
  XNOR2_X1 U521 ( .A(KEYINPUT25), .B(n462), .ZN(n463) );
  NAND2_X1 U522 ( .A1(n464), .A2(n463), .ZN(n465) );
  NOR2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  NOR2_X1 U524 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n471), .A2(n472), .ZN(n473) );
  XNOR2_X1 U526 ( .A(KEYINPUT16), .B(n473), .ZN(n474) );
  NOR2_X1 U527 ( .A1(n487), .A2(n474), .ZN(n475) );
  XOR2_X1 U528 ( .A(KEYINPUT95), .B(n475), .Z(n503) );
  NOR2_X1 U529 ( .A1(n579), .A2(n573), .ZN(n476) );
  XNOR2_X1 U530 ( .A(n476), .B(KEYINPUT72), .ZN(n491) );
  NAND2_X1 U531 ( .A1(n503), .A2(n491), .ZN(n483) );
  NOR2_X1 U532 ( .A1(n530), .A2(n483), .ZN(n477) );
  XOR2_X1 U533 ( .A(G1GAT), .B(n477), .Z(n478) );
  XNOR2_X1 U534 ( .A(KEYINPUT34), .B(n478), .ZN(G1324GAT) );
  NOR2_X1 U535 ( .A1(n518), .A2(n483), .ZN(n479) );
  XOR2_X1 U536 ( .A(G8GAT), .B(n479), .Z(G1325GAT) );
  NOR2_X1 U537 ( .A1(n533), .A2(n483), .ZN(n481) );
  XNOR2_X1 U538 ( .A(KEYINPUT35), .B(KEYINPUT96), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U541 ( .A1(n525), .A2(n483), .ZN(n485) );
  XNOR2_X1 U542 ( .A(G22GAT), .B(KEYINPUT97), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1327GAT) );
  XNOR2_X1 U544 ( .A(KEYINPUT39), .B(KEYINPUT99), .ZN(n494) );
  NOR2_X1 U545 ( .A1(n486), .A2(n487), .ZN(n488) );
  NAND2_X1 U546 ( .A1(n585), .A2(n488), .ZN(n489) );
  XNOR2_X1 U547 ( .A(KEYINPUT37), .B(n489), .ZN(n490) );
  XNOR2_X1 U548 ( .A(KEYINPUT98), .B(n490), .ZN(n515) );
  NAND2_X1 U549 ( .A1(n515), .A2(n491), .ZN(n492) );
  NOR2_X1 U550 ( .A1(n530), .A2(n500), .ZN(n493) );
  XNOR2_X1 U551 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U552 ( .A(n495), .B(G29GAT), .Z(G1328GAT) );
  NOR2_X1 U553 ( .A1(n518), .A2(n500), .ZN(n496) );
  XOR2_X1 U554 ( .A(G36GAT), .B(n496), .Z(G1329GAT) );
  NOR2_X1 U555 ( .A1(n500), .A2(n533), .ZN(n498) );
  XNOR2_X1 U556 ( .A(KEYINPUT40), .B(KEYINPUT100), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U558 ( .A(G43GAT), .B(n499), .Z(G1330GAT) );
  XNOR2_X1 U559 ( .A(G50GAT), .B(KEYINPUT101), .ZN(n502) );
  NOR2_X1 U560 ( .A1(n525), .A2(n500), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n502), .B(n501), .ZN(G1331GAT) );
  XNOR2_X1 U562 ( .A(KEYINPUT102), .B(n552), .ZN(n558) );
  NOR2_X1 U563 ( .A1(n558), .A2(n534), .ZN(n516) );
  NAND2_X1 U564 ( .A1(n503), .A2(n516), .ZN(n511) );
  NOR2_X1 U565 ( .A1(n530), .A2(n511), .ZN(n505) );
  XNOR2_X1 U566 ( .A(KEYINPUT103), .B(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U569 ( .A1(n518), .A2(n511), .ZN(n507) );
  XOR2_X1 U570 ( .A(KEYINPUT104), .B(n507), .Z(n508) );
  XNOR2_X1 U571 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U572 ( .A1(n533), .A2(n511), .ZN(n510) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(G1334GAT) );
  NOR2_X1 U575 ( .A1(n525), .A2(n511), .ZN(n513) );
  XNOR2_X1 U576 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(n514), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n516), .A2(n515), .ZN(n524) );
  NOR2_X1 U580 ( .A1(n530), .A2(n524), .ZN(n517) );
  XOR2_X1 U581 ( .A(G85GAT), .B(n517), .Z(G1336GAT) );
  NOR2_X1 U582 ( .A1(n518), .A2(n524), .ZN(n520) );
  XNOR2_X1 U583 ( .A(G92GAT), .B(KEYINPUT107), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(G1337GAT) );
  NOR2_X1 U585 ( .A1(n533), .A2(n524), .ZN(n522) );
  XNOR2_X1 U586 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(n523), .ZN(G1338GAT) );
  NOR2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n527) );
  XNOR2_X1 U590 ( .A(KEYINPUT110), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U592 ( .A(G106GAT), .B(n528), .Z(G1339GAT) );
  NOR2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n547) );
  NAND2_X1 U594 ( .A1(n531), .A2(n547), .ZN(n532) );
  NOR2_X1 U595 ( .A1(n533), .A2(n532), .ZN(n536) );
  NAND2_X1 U596 ( .A1(n536), .A2(n534), .ZN(n535) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  INV_X1 U598 ( .A(n536), .ZN(n543) );
  NOR2_X1 U599 ( .A1(n558), .A2(n543), .ZN(n538) );
  XNOR2_X1 U600 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U602 ( .A(G120GAT), .B(n539), .Z(G1341GAT) );
  NOR2_X1 U603 ( .A1(n563), .A2(n543), .ZN(n541) );
  XNOR2_X1 U604 ( .A(KEYINPUT116), .B(KEYINPUT50), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U606 ( .A(G127GAT), .B(n542), .Z(G1342GAT) );
  NOR2_X1 U607 ( .A1(n471), .A2(n543), .ZN(n545) );
  XNOR2_X1 U608 ( .A(KEYINPUT117), .B(KEYINPUT51), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U610 ( .A(G134GAT), .B(n546), .Z(G1343GAT) );
  NAND2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n556) );
  NOR2_X1 U612 ( .A1(n573), .A2(n556), .ZN(n549) );
  XOR2_X1 U613 ( .A(G141GAT), .B(n549), .Z(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n551) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n554) );
  NOR2_X1 U617 ( .A1(n552), .A2(n556), .ZN(n553) );
  XOR2_X1 U618 ( .A(n554), .B(n553), .Z(G1345GAT) );
  NOR2_X1 U619 ( .A1(n585), .A2(n556), .ZN(n555) );
  XOR2_X1 U620 ( .A(G155GAT), .B(n555), .Z(G1346GAT) );
  NOR2_X1 U621 ( .A1(n471), .A2(n556), .ZN(n557) );
  XOR2_X1 U622 ( .A(G162GAT), .B(n557), .Z(G1347GAT) );
  NOR2_X1 U623 ( .A1(n558), .A2(n567), .ZN(n560) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(n562) );
  XOR2_X1 U626 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  NOR2_X1 U628 ( .A1(n563), .A2(n567), .ZN(n565) );
  INV_X1 U629 ( .A(KEYINPUT122), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U632 ( .A1(n567), .A2(n471), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G190GAT), .B(n570), .ZN(G1351GAT) );
  OR2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n587) );
  NOR2_X1 U637 ( .A1(n573), .A2(n587), .ZN(n578) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n575) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(KEYINPUT124), .B(n576), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  INV_X1 U643 ( .A(n579), .ZN(n580) );
  NOR2_X1 U644 ( .A1(n587), .A2(n580), .ZN(n584) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n582) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n587), .ZN(n586) );
  XOR2_X1 U650 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
  NOR2_X1 U651 ( .A1(n486), .A2(n587), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

