//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n454), .A2(new_n458), .B1(new_n449), .B2(new_n455), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT66), .Z(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT70), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n464), .B1(new_n465), .B2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  OR2_X1    g046(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(G137), .A3(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n471), .A2(KEYINPUT69), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n477), .B1(new_n470), .B2(new_n474), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n463), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n467), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n482), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n483));
  INV_X1    g058(.A(new_n473), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OR2_X1    g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n479), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G160));
  NOR2_X1   g064(.A1(new_n470), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n470), .A2(new_n486), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  OAI221_X1 g068(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n486), .C2(G112), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  XOR2_X1   g070(.A(new_n495), .B(KEYINPUT71), .Z(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  NAND3_X1  g072(.A1(new_n472), .A2(G138), .A3(new_n473), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n498), .A2(new_n481), .A3(KEYINPUT4), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT4), .B1(new_n470), .B2(new_n498), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(KEYINPUT73), .B(KEYINPUT4), .C1(new_n470), .C2(new_n498), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(G126), .A2(G2105), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n466), .A2(new_n469), .A3(new_n467), .A4(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n507), .A2(new_n508), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n461), .A2(G114), .ZN(new_n511));
  OAI21_X1  g086(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(KEYINPUT74), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT5), .A3(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n522), .A2(G62), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  XOR2_X1   g099(.A(new_n524), .B(KEYINPUT75), .Z(new_n525));
  OAI21_X1  g100(.A(G651), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT76), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT76), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n528), .B(G651), .C1(new_n523), .C2(new_n525), .ZN(new_n529));
  OR2_X1    g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n522), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n517), .B1(new_n530), .B2(new_n531), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n534), .A2(G88), .B1(G50), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n527), .A2(new_n529), .A3(new_n536), .ZN(G303));
  INV_X1    g112(.A(G303), .ZN(G166));
  AND2_X1   g113(.A1(new_n534), .A2(G89), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n535), .A2(G51), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n539), .A2(new_n544), .ZN(G168));
  AOI22_X1  g120(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G651), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n535), .A2(G52), .ZN(new_n549));
  INV_X1    g124(.A(G90), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n533), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(G171));
  AND2_X1   g127(.A1(G68), .A2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n522), .B2(G56), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(new_n547), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT77), .ZN(new_n556));
  OR3_X1    g131(.A1(new_n554), .A2(KEYINPUT77), .A3(new_n547), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n535), .A2(G43), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n533), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n556), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT78), .ZN(G188));
  NAND2_X1  g144(.A1(new_n535), .A2(G53), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT79), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g148(.A(KEYINPUT79), .B(KEYINPUT9), .Z(new_n574));
  NAND3_X1  g149(.A1(new_n535), .A2(new_n574), .A3(G53), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n573), .A2(KEYINPUT80), .A3(new_n575), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n519), .A2(new_n581), .A3(new_n521), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n581), .B1(new_n519), .B2(new_n521), .ZN(new_n583));
  OAI21_X1  g158(.A(G65), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(G78), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n517), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n547), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n534), .A2(G91), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n580), .A2(new_n591), .ZN(G299));
  INV_X1    g167(.A(G171), .ZN(G301));
  INV_X1    g168(.A(G168), .ZN(G286));
  AOI22_X1  g169(.A1(new_n534), .A2(G87), .B1(G49), .B2(new_n535), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G288));
  AOI22_X1  g172(.A1(new_n534), .A2(G86), .B1(G48), .B2(new_n535), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n522), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n547), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n598), .A2(new_n600), .ZN(G305));
  AOI22_X1  g176(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n547), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n535), .A2(G47), .ZN(new_n604));
  INV_X1    g179(.A(G85), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n533), .B2(new_n605), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n603), .A2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT82), .ZN(new_n609));
  AND3_X1   g184(.A1(new_n520), .A2(KEYINPUT5), .A3(G543), .ZN(new_n610));
  AOI21_X1  g185(.A(G543), .B1(new_n520), .B2(KEYINPUT5), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT81), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n519), .A2(new_n581), .A3(new_n521), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g189(.A1(new_n614), .A2(G66), .ZN(new_n615));
  AND2_X1   g190(.A1(G79), .A2(G543), .ZN(new_n616));
  OAI21_X1  g191(.A(G651), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n534), .A2(KEYINPUT10), .A3(G92), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT10), .ZN(new_n619));
  INV_X1    g194(.A(G92), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n533), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n618), .A2(new_n621), .B1(G54), .B2(new_n535), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n609), .B1(G868), .B2(new_n623), .ZN(G284));
  OAI21_X1  g199(.A(new_n609), .B1(G868), .B2(new_n623), .ZN(G321));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n586), .B1(new_n614), .B2(G65), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n589), .B1(new_n627), .B2(new_n547), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n578), .B2(new_n579), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n626), .B1(new_n629), .B2(G868), .ZN(G297));
  OAI21_X1  g205(.A(new_n626), .B1(new_n629), .B2(G868), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n623), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND2_X1  g208(.A1(new_n623), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g212(.A1(new_n468), .A2(G2105), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n482), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT13), .ZN(new_n641));
  AOI22_X1  g216(.A1(new_n640), .A2(new_n641), .B1(KEYINPUT83), .B2(G2100), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(new_n643));
  NOR2_X1   g218(.A1(KEYINPUT83), .A2(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n490), .A2(G135), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT84), .Z(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  INV_X1    g223(.A(new_n486), .ZN(new_n649));
  INV_X1    g224(.A(G111), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n492), .B2(G123), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n653), .A2(G2096), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(G2096), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n645), .A2(new_n654), .A3(new_n655), .ZN(G156));
  XOR2_X1   g231(.A(G2451), .B(G2454), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT14), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2427), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2430), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT15), .B(G2435), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n664), .B2(new_n663), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n660), .B(new_n666), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2443), .B(G2446), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g245(.A(G14), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n670), .B2(new_n668), .ZN(G401));
  XNOR2_X1  g247(.A(G2072), .B(G2078), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT17), .Z(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(new_n675), .B2(new_n673), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT85), .Z(new_n682));
  NAND3_X1  g257(.A1(new_n678), .A2(new_n675), .A3(new_n673), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT18), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n679), .A2(new_n675), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n674), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G2096), .B(G2100), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G227));
  XOR2_X1   g264(.A(G1971), .B(G1976), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1956), .B(G2474), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1961), .B(G1966), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(new_n694), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT20), .Z(new_n698));
  AOI211_X1 g273(.A(new_n696), .B(new_n698), .C1(new_n691), .C2(new_n695), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT86), .ZN(new_n700));
  XOR2_X1   g275(.A(G1981), .B(G1986), .Z(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n700), .B(new_n705), .ZN(G229));
  NOR2_X1   g281(.A1(G16), .A2(G24), .ZN(new_n707));
  XNOR2_X1  g282(.A(G290), .B(KEYINPUT87), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(G16), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT88), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G1986), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G25), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n490), .A2(G131), .ZN(new_n714));
  OAI221_X1 g289(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n486), .C2(G107), .ZN(new_n715));
  INV_X1    g290(.A(new_n492), .ZN(new_n716));
  INV_X1    g291(.A(G119), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n714), .B(new_n715), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n713), .B1(new_n719), .B2(new_n712), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT35), .B(G1991), .Z(new_n721));
  XOR2_X1   g296(.A(new_n720), .B(new_n721), .Z(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(KEYINPUT90), .B2(KEYINPUT36), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n711), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(G6), .A2(G16), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n598), .A2(new_n600), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(G16), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT32), .ZN(new_n729));
  INV_X1    g304(.A(G1981), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(G303), .A2(G16), .ZN(new_n732));
  INV_X1    g307(.A(G1971), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G22), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT89), .Z(new_n736));
  NAND3_X1  g311(.A1(new_n732), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n734), .A2(G23), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n595), .A2(new_n596), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(new_n734), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT33), .B(G1976), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n733), .B1(new_n732), .B2(new_n736), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n731), .A2(new_n737), .A3(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(KEYINPUT34), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(KEYINPUT34), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n725), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(KEYINPUT90), .B2(KEYINPUT36), .ZN(new_n749));
  NOR2_X1   g324(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n725), .A2(new_n750), .A3(new_n746), .A4(new_n747), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(G115), .A2(G2104), .ZN(new_n753));
  INV_X1    g328(.A(G127), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n481), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(new_n649), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n486), .A2(G103), .A3(G2104), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT94), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(KEYINPUT25), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n758), .A2(KEYINPUT94), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n758), .A2(KEYINPUT94), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n490), .A2(G139), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n765), .A2(KEYINPUT95), .A3(new_n766), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n757), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT96), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI211_X1 g348(.A(KEYINPUT96), .B(new_n757), .C1(new_n769), .C2(new_n770), .ZN(new_n774));
  OAI21_X1  g349(.A(G29), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G33), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(G29), .B2(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(G2072), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(G2072), .ZN(new_n779));
  OAI21_X1  g354(.A(KEYINPUT97), .B1(G29), .B2(G32), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n490), .A2(G141), .ZN(new_n781));
  NAND3_X1  g356(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT26), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n784), .A2(new_n785), .B1(G105), .B2(new_n638), .ZN(new_n786));
  INV_X1    g361(.A(G129), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n781), .B(new_n786), .C1(new_n716), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(new_n712), .ZN(new_n789));
  MUX2_X1   g364(.A(new_n780), .B(KEYINPUT97), .S(new_n789), .Z(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT27), .B(G1996), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT24), .ZN(new_n792));
  INV_X1    g367(.A(G34), .ZN(new_n793));
  AOI21_X1  g368(.A(G29), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n792), .B2(new_n793), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G160), .B2(new_n712), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n790), .A2(new_n791), .B1(G2084), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n778), .A2(new_n779), .A3(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(KEYINPUT98), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n712), .A2(G35), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G162), .B2(new_n712), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2090), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n802), .B(new_n803), .Z(new_n804));
  NOR2_X1   g379(.A1(G4), .A2(G16), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n623), .B2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT91), .B(G1348), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(G1341), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n563), .A2(G16), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G16), .B2(G19), .ZN(new_n811));
  OAI221_X1 g386(.A(new_n808), .B1(new_n809), .B2(new_n811), .C1(G2084), .C2(new_n796), .ZN(new_n812));
  NOR2_X1   g387(.A1(G168), .A2(new_n734), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n734), .B2(G21), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT99), .B(G1966), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT30), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n817), .A2(G28), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n712), .B1(new_n817), .B2(G28), .ZN(new_n819));
  AND2_X1   g394(.A1(KEYINPUT31), .A2(G11), .ZN(new_n820));
  NOR2_X1   g395(.A1(KEYINPUT31), .A2(G11), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n818), .A2(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n653), .ZN(new_n823));
  NOR2_X1   g398(.A1(G171), .A2(new_n734), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G5), .B2(new_n734), .ZN(new_n825));
  INV_X1    g400(.A(G1961), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n823), .A2(G29), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n814), .A2(new_n815), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n827), .B(new_n828), .C1(new_n826), .C2(new_n825), .ZN(new_n829));
  NOR4_X1   g404(.A1(new_n812), .A2(new_n816), .A3(new_n822), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n734), .A2(G20), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT23), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n629), .B2(new_n734), .ZN(new_n833));
  INV_X1    g408(.A(G1956), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n811), .A2(new_n809), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n791), .B2(new_n790), .ZN(new_n837));
  NOR2_X1   g412(.A1(G27), .A2(G29), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G164), .B2(G29), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G2078), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n712), .A2(G26), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT28), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n843));
  INV_X1    g418(.A(G116), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n649), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n490), .B2(G140), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n492), .A2(G128), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n847), .A2(KEYINPUT92), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(KEYINPUT92), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n842), .B1(new_n851), .B2(new_n712), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT93), .B(G2067), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NOR3_X1   g429(.A1(new_n837), .A2(new_n840), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n804), .A2(new_n830), .A3(new_n835), .A4(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n798), .B2(KEYINPUT98), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n752), .A2(new_n799), .A3(new_n857), .ZN(G150));
  INV_X1    g433(.A(G150), .ZN(G311));
  AOI22_X1  g434(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(new_n547), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n535), .A2(G55), .ZN(new_n862));
  INV_X1    g437(.A(G93), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n862), .B1(new_n533), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(G860), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT37), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n623), .A2(G559), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n562), .A2(new_n866), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n560), .B1(new_n555), .B2(KEYINPUT77), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(new_n557), .A3(new_n865), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n870), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT39), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT101), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n879));
  INV_X1    g454(.A(new_n875), .ZN(new_n880));
  AOI21_X1  g455(.A(G860), .B1(new_n880), .B2(KEYINPUT39), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n879), .B1(new_n878), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n868), .B1(new_n882), .B2(new_n883), .ZN(G145));
  NAND2_X1  g459(.A1(new_n769), .A2(new_n770), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n756), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT96), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n771), .A2(new_n772), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT104), .B1(new_n773), .B2(new_n774), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n515), .B(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n788), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n515), .B(KEYINPUT103), .ZN(new_n895));
  INV_X1    g470(.A(new_n788), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(new_n897), .A3(new_n850), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n850), .B1(new_n894), .B2(new_n897), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n890), .B(new_n891), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n888), .B1(new_n887), .B2(new_n889), .ZN(new_n902));
  INV_X1    g477(.A(new_n900), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(new_n903), .A3(new_n898), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n490), .A2(G142), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n492), .A2(G130), .ZN(new_n906));
  OAI221_X1 g481(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n486), .C2(G118), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n640), .B(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(new_n718), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n901), .A2(new_n904), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n823), .A2(new_n488), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n653), .A2(G160), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(G162), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT106), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n901), .A2(new_n904), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n910), .B(KEYINPUT105), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n911), .B(new_n916), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n901), .A2(new_n918), .A3(new_n904), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n918), .B1(new_n901), .B2(new_n904), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n915), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n919), .A2(new_n922), .A3(new_n923), .A4(new_n925), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(G395));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n930));
  INV_X1    g505(.A(G290), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(G303), .ZN(new_n932));
  NAND4_X1  g507(.A1(G290), .A2(new_n529), .A3(new_n527), .A4(new_n536), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n739), .A2(G305), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n727), .A2(G288), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n932), .A2(new_n933), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  AOI22_X1  g512(.A1(new_n932), .A2(new_n933), .B1(new_n935), .B2(new_n934), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n930), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n932), .A2(new_n933), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n935), .A2(new_n934), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(KEYINPUT108), .A3(new_n936), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT42), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n936), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(KEYINPUT42), .B2(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n874), .B(new_n634), .Z(new_n948));
  NAND2_X1  g523(.A1(new_n629), .A2(new_n623), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n617), .A2(new_n622), .ZN(new_n950));
  NAND2_X1  g525(.A1(G299), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT41), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n949), .A2(KEYINPUT41), .A3(new_n951), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n948), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n952), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n957), .B1(new_n958), .B2(new_n948), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n947), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n947), .A2(new_n959), .ZN(new_n961));
  OAI21_X1  g536(.A(G868), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(G868), .B2(new_n865), .ZN(G295));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n964));
  XNOR2_X1  g539(.A(G295), .B(new_n964), .ZN(G331));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n871), .A2(G301), .A3(new_n873), .ZN(new_n967));
  AOI21_X1  g542(.A(G301), .B1(new_n871), .B2(new_n873), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n967), .A2(new_n968), .A3(G286), .ZN(new_n969));
  INV_X1    g544(.A(new_n873), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n865), .B1(new_n872), .B2(new_n557), .ZN(new_n971));
  OAI21_X1  g546(.A(G171), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n871), .A2(G301), .A3(new_n873), .ZN(new_n973));
  AOI21_X1  g548(.A(G168), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n958), .B1(new_n969), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(G286), .B1(new_n967), .B2(new_n968), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(G168), .A3(new_n973), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n976), .A2(new_n954), .A3(new_n977), .A4(new_n955), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n944), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n923), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n944), .B1(new_n975), .B2(new_n978), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n980), .A2(KEYINPUT43), .A3(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n969), .A2(new_n974), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n954), .A2(new_n955), .ZN(new_n984));
  AOI22_X1  g559(.A1(KEYINPUT110), .A2(new_n975), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n986), .B(new_n958), .C1(new_n969), .C2(new_n974), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n944), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT43), .B1(new_n988), .B2(new_n980), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n982), .B1(new_n989), .B2(KEYINPUT112), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n975), .A2(KEYINPUT110), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(new_n987), .A3(new_n978), .ZN(new_n992));
  INV_X1    g567(.A(new_n944), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n980), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n995));
  OR3_X1    g570(.A1(new_n994), .A2(KEYINPUT112), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n966), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n992), .A2(new_n993), .ZN(new_n999));
  INV_X1    g574(.A(new_n980), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n995), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT43), .B1(new_n980), .B2(new_n981), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT111), .B1(new_n994), .B2(new_n995), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n1003), .A2(new_n1004), .A3(KEYINPUT44), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n997), .A2(new_n1005), .ZN(G397));
  INV_X1    g581(.A(G1384), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n504), .B2(new_n513), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n479), .A2(new_n487), .A3(G40), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1996), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT46), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1012), .ZN(new_n1016));
  INV_X1    g591(.A(G2067), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n850), .B(new_n1017), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1018), .A2(new_n896), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1015), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT47), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1021), .A2(KEYINPUT127), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(KEYINPUT127), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n788), .B(new_n1013), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1018), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1025), .A2(new_n721), .A3(new_n719), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n851), .A2(new_n1017), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1016), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n718), .B(new_n721), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1016), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(G290), .A2(G1986), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT48), .B1(new_n1012), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1012), .A2(KEYINPUT48), .A3(new_n1031), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1028), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1022), .A2(new_n1023), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(G303), .A2(G8), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1037), .B(KEYINPUT55), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1008), .A2(KEYINPUT50), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1041), .B(new_n1007), .C1(new_n504), .C2(new_n513), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1011), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(G2090), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1011), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT45), .B(new_n1007), .C1(new_n504), .C2(new_n513), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1971), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1039), .B(G8), .C1(new_n1045), .C2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n739), .A2(G1976), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1050), .B(G8), .C1(new_n1008), .C2(new_n1011), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n739), .A2(G1976), .ZN(new_n1052));
  OR3_X1    g627(.A1(new_n1051), .A2(KEYINPUT52), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(KEYINPUT49), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n598), .A2(new_n600), .A3(new_n730), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1056), .B1(new_n1057), .B2(KEYINPUT114), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n727), .A2(new_n730), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1057), .A2(KEYINPUT114), .A3(new_n1056), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1057), .A2(KEYINPUT114), .A3(new_n1056), .ZN(new_n1063));
  OAI22_X1  g638(.A1(new_n1063), .A2(new_n1058), .B1(new_n730), .B2(new_n727), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1065));
  INV_X1    g640(.A(G8), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1062), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1051), .A2(KEYINPUT52), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1053), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(G288), .A2(G1976), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1068), .A2(new_n1071), .B1(new_n730), .B2(new_n727), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1067), .ZN(new_n1073));
  OAI22_X1  g648(.A1(new_n1049), .A2(new_n1070), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT63), .ZN(new_n1075));
  OAI21_X1  g650(.A(G8), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1038), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1053), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(new_n1049), .ZN(new_n1079));
  INV_X1    g654(.A(G2084), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1040), .A2(new_n1080), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT116), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1010), .A2(new_n1043), .A3(new_n1047), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n815), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1011), .B1(new_n1008), .B2(KEYINPUT50), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1085), .A2(new_n1086), .A3(new_n1080), .A4(new_n1042), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1082), .A2(new_n1084), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(G8), .A3(G168), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1075), .B1(new_n1079), .B2(new_n1089), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1044), .A2(G2090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1048), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1066), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1070), .B1(new_n1093), .B2(new_n1039), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1089), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1094), .A2(KEYINPUT63), .A3(new_n1095), .A4(new_n1077), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1074), .B1(new_n1090), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G2078), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1046), .A2(new_n1098), .A3(new_n1047), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1044), .A2(new_n826), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1100), .A2(G2078), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1046), .A2(new_n1047), .A3(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(G171), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1079), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1082), .A2(new_n1084), .A3(G168), .A4(new_n1087), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1108), .A2(new_n1109), .A3(G8), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1088), .A2(G286), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(G8), .A3(new_n1108), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1110), .B1(new_n1112), .B2(KEYINPUT51), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1107), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1088), .A2(G286), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1108), .A2(G8), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT51), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1110), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n1114), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1097), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n1123));
  OAI211_X1 g698(.A(G40), .B(new_n487), .C1(new_n479), .C2(new_n1123), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n479), .A2(new_n1123), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n1010), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1010), .A3(KEYINPUT124), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1047), .A2(new_n1103), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1099), .A2(new_n1100), .B1(new_n1044), .B2(new_n826), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(new_n1133), .A3(G301), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT54), .B1(new_n1106), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1135), .A2(new_n1079), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT125), .B1(new_n1105), .B2(G171), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(G171), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1133), .A2(new_n1140), .A3(G301), .A4(new_n1104), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1137), .A2(new_n1139), .A3(KEYINPUT54), .A4(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1122), .A2(new_n1136), .A3(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1010), .A2(new_n1013), .A3(new_n1043), .A4(new_n1047), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(G1341), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(new_n563), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT57), .ZN(new_n1151));
  NOR2_X1   g726(.A1(G299), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n576), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(new_n628), .B2(KEYINPUT117), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1155), .B(new_n589), .C1(new_n627), .C2(new_n547), .ZN(new_n1156));
  AOI21_X1  g731(.A(KEYINPUT57), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT118), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1152), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT117), .B1(new_n588), .B2(new_n590), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1160), .A2(new_n576), .A3(new_n1156), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1158), .B1(new_n1161), .B2(new_n1151), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT56), .B(G2072), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1046), .A2(new_n1047), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(G1956), .B1(new_n1085), .B2(new_n1042), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1159), .B(new_n1163), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1044), .A2(new_n834), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1046), .A2(new_n1047), .A3(new_n1164), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1161), .A2(new_n1158), .A3(new_n1151), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n629), .A2(KEYINPUT57), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1168), .B(new_n1169), .C1(new_n1172), .C2(new_n1162), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1167), .A2(KEYINPUT61), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1044), .A2(new_n807), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1008), .A2(G2067), .A3(new_n1011), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n950), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  AOI211_X1 g753(.A(new_n623), .B(new_n1176), .C1(new_n1044), .C2(new_n807), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT60), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1148), .A2(new_n563), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT120), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1176), .B1(new_n1044), .B2(new_n807), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n950), .A2(KEYINPUT60), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1181), .A2(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AND4_X1   g761(.A1(new_n1150), .A2(new_n1174), .A3(new_n1180), .A4(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT121), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1167), .A2(new_n1188), .A3(new_n1173), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1190), .A2(KEYINPUT121), .A3(new_n1163), .A4(new_n1159), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(KEYINPUT122), .B1(new_n1189), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1167), .A2(new_n1188), .A3(new_n1173), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT122), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1195), .A2(new_n1196), .A3(new_n1192), .A4(new_n1191), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1187), .A2(new_n1194), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1167), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1173), .B1(new_n1199), .B2(new_n1178), .ZN(new_n1200));
  AOI22_X1  g775(.A1(KEYINPUT126), .A2(new_n1143), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1122), .A2(new_n1136), .A3(new_n1202), .A4(new_n1142), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1121), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1030), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1031), .A2(KEYINPUT113), .ZN(new_n1206));
  NAND2_X1  g781(.A1(G290), .A2(G1986), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1206), .B(new_n1207), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1205), .B1(new_n1016), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1036), .B1(new_n1204), .B2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g785(.A1(G229), .A2(G227), .A3(G401), .A4(new_n459), .ZN(new_n1212));
  NAND2_X1  g786(.A1(new_n924), .A2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g787(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1214));
  NOR2_X1   g788(.A1(new_n1213), .A2(new_n1214), .ZN(G308));
  OAI211_X1 g789(.A(new_n924), .B(new_n1212), .C1(new_n1003), .C2(new_n1004), .ZN(G225));
endmodule


