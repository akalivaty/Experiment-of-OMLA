//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1289, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G107), .ZN(new_n220));
  INV_X1    g0020(.A(G264), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n211), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT66), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n211), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n214), .B(new_n227), .C1(new_n216), .C2(new_n221), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n228), .A2(KEYINPUT0), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(KEYINPUT0), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n202), .A2(new_n203), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n233), .A2(G20), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n229), .A2(new_n230), .A3(new_n236), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n225), .B(new_n237), .C1(KEYINPUT1), .C2(new_n223), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n219), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n208), .A2(G20), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NOR3_X1   g0056(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT72), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n234), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT72), .B1(new_n254), .B2(new_n256), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n262), .A2(new_n263), .B1(new_n254), .B2(new_n259), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n268), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n269));
  AOI21_X1  g0069(.A(KEYINPUT70), .B1(new_n268), .B2(KEYINPUT3), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n267), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT7), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(new_n272), .A3(new_n209), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT70), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(new_n266), .B2(G33), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n268), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT7), .B1(new_n278), .B2(G20), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n273), .A2(new_n279), .A3(G68), .ZN(new_n280));
  XNOR2_X1  g0080(.A(G58), .B(G68), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n281), .A2(G20), .B1(G159), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(KEYINPUT16), .A3(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n284), .A2(new_n261), .ZN(new_n285));
  OAI21_X1  g0085(.A(KEYINPUT71), .B1(new_n266), .B2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT71), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(new_n268), .A3(KEYINPUT3), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n274), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT7), .B1(new_n289), .B2(G20), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n267), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(new_n272), .A3(new_n209), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(G68), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n283), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT16), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n265), .B1(new_n285), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G87), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT73), .ZN(new_n301));
  MUX2_X1   g0101(.A(G223), .B(G226), .S(G1698), .Z(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(new_n278), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G41), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(G1), .A3(G13), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n299), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n208), .B(G274), .C1(G41), .C2(G45), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n307), .B1(new_n309), .B2(new_n219), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT74), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(KEYINPUT74), .B(new_n307), .C1(new_n309), .C2(new_n219), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n306), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n276), .A2(new_n277), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(new_n302), .A3(new_n267), .ZN(new_n317));
  INV_X1    g0117(.A(new_n301), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n305), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n310), .ZN(new_n322));
  AOI21_X1  g0122(.A(G200), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT76), .B1(new_n315), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n305), .B1(new_n317), .B2(new_n318), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n310), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT76), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n327), .B(new_n328), .C1(new_n314), .C2(new_n306), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n298), .A2(KEYINPUT17), .A3(new_n324), .A4(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT17), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n324), .A2(new_n329), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n284), .A2(new_n261), .ZN(new_n333));
  AOI21_X1  g0133(.A(KEYINPUT16), .B1(new_n294), .B2(new_n283), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n264), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n331), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n321), .A2(new_n338), .A3(new_n312), .A4(new_n313), .ZN(new_n339));
  INV_X1    g0139(.A(G169), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n326), .B2(new_n310), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n297), .A2(new_n261), .A3(new_n284), .ZN(new_n343));
  AOI211_X1 g0143(.A(KEYINPUT18), .B(new_n342), .C1(new_n343), .C2(new_n264), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT18), .ZN(new_n345));
  INV_X1    g0145(.A(new_n342), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n335), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT75), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n335), .A2(new_n346), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT18), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT75), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n335), .A2(new_n346), .A3(new_n345), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n337), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n204), .A2(G20), .ZN(new_n355));
  XOR2_X1   g0155(.A(KEYINPUT8), .B(G58), .Z(new_n356));
  NOR2_X1   g0156(.A1(new_n268), .A2(G20), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n356), .A2(new_n357), .B1(G150), .B2(new_n282), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n261), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n259), .A2(new_n261), .ZN(new_n361));
  INV_X1    g0161(.A(G50), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n256), .A2(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n361), .A2(new_n363), .B1(new_n362), .B2(new_n259), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT9), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT3), .B(G33), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(G223), .A3(G1698), .ZN(new_n369));
  INV_X1    g0169(.A(G1698), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(G222), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G77), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n369), .B(new_n371), .C1(new_n372), .C2(new_n368), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n320), .ZN(new_n374));
  INV_X1    g0174(.A(new_n307), .ZN(new_n375));
  INV_X1    g0175(.A(new_n309), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(G226), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G200), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n360), .A2(KEYINPUT9), .A3(new_n364), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n367), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT68), .B1(new_n378), .B2(new_n299), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT10), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT68), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n374), .A2(new_n384), .A3(G190), .A4(new_n377), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n381), .A2(new_n382), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n367), .A2(new_n385), .A3(new_n379), .A4(new_n380), .ZN(new_n387));
  INV_X1    g0187(.A(new_n382), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT10), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n378), .A2(G169), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n338), .B2(new_n378), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n365), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G13), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n396), .A2(G1), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(G20), .A3(new_n203), .ZN(new_n398));
  XOR2_X1   g0198(.A(new_n398), .B(KEYINPUT12), .Z(new_n399));
  NAND2_X1  g0199(.A1(new_n357), .A2(G77), .ZN(new_n400));
  INV_X1    g0200(.A(new_n282), .ZN(new_n401));
  OAI221_X1 g0201(.A(new_n400), .B1(new_n209), .B2(G68), .C1(new_n362), .C2(new_n401), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n402), .A2(new_n261), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n399), .B1(KEYINPUT11), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT67), .B1(new_n259), .B2(new_n261), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT67), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n258), .A2(new_n406), .A3(new_n234), .A4(new_n260), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n405), .A2(G68), .A3(new_n255), .A4(new_n407), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n404), .B(new_n408), .C1(KEYINPUT11), .C2(new_n403), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n368), .A2(G226), .A3(new_n370), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n368), .A2(G232), .A3(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G97), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n320), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n375), .B1(new_n376), .B2(G238), .ZN(new_n415));
  XNOR2_X1  g0215(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n415), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT13), .ZN(new_n420));
  OAI211_X1 g0220(.A(G179), .B(new_n417), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n416), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n340), .B1(new_n423), .B2(new_n417), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT14), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n417), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n416), .B1(new_n414), .B2(new_n415), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n425), .B(G169), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n409), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT15), .B(G87), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n433), .A2(new_n357), .B1(G20), .B2(G77), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n254), .B2(new_n401), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n261), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n405), .A2(G77), .A3(new_n255), .A4(new_n407), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n259), .A2(new_n372), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n368), .A2(G232), .A3(new_n370), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n220), .B2(new_n368), .ZN(new_n441));
  INV_X1    g0241(.A(G238), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n292), .A2(new_n442), .A3(new_n370), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n320), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n375), .B1(new_n376), .B2(G244), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n444), .A2(G179), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n340), .B1(new_n444), .B2(new_n445), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n439), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n444), .A2(new_n299), .A3(new_n445), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(G200), .B1(new_n444), .B2(new_n445), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n448), .B1(new_n452), .B2(new_n439), .ZN(new_n453));
  OAI211_X1 g0253(.A(G190), .B(new_n417), .C1(new_n419), .C2(new_n420), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n325), .B1(new_n423), .B2(new_n417), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(new_n409), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n453), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AND4_X1   g0257(.A1(new_n354), .A2(new_n395), .A3(new_n431), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G116), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n208), .B2(G33), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n405), .A2(new_n407), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n397), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(G20), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT81), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT81), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n397), .A2(new_n465), .A3(G20), .A4(new_n459), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n260), .A2(new_n234), .B1(G20), .B2(new_n459), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G283), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n470), .B(new_n209), .C1(G33), .C2(new_n215), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(KEYINPUT20), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT20), .B1(new_n469), .B2(new_n471), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT82), .B1(new_n468), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n474), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n472), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT82), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n478), .A2(new_n479), .A3(new_n461), .A4(new_n467), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G264), .A2(G1698), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n216), .B2(G1698), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n267), .B(new_n483), .C1(new_n269), .C2(new_n270), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n292), .A2(G303), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n305), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G41), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n208), .B(G45), .C1(new_n487), .C2(KEYINPUT5), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT5), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G41), .ZN(new_n490));
  OAI211_X1 g0290(.A(G270), .B(new_n305), .C1(new_n488), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(G41), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(new_n208), .A3(G45), .A4(G274), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT78), .B1(new_n489), .B2(G41), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT78), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(new_n487), .A3(KEYINPUT5), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n491), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(KEYINPUT21), .B(G169), .C1(new_n486), .C2(new_n498), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n497), .A2(new_n493), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n278), .A2(new_n483), .B1(G303), .B2(new_n292), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n491), .B(new_n500), .C1(new_n501), .C2(new_n305), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n499), .B1(new_n338), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n481), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n486), .A2(new_n498), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(G200), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n486), .A2(new_n498), .A3(G190), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n480), .B(new_n476), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(G169), .B1(new_n486), .B2(new_n498), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n509), .B1(new_n476), .B2(new_n480), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n504), .B(new_n508), .C1(KEYINPUT21), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT83), .ZN(new_n512));
  INV_X1    g0312(.A(new_n509), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n481), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT21), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT83), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(new_n508), .A4(new_n504), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n433), .A2(new_n258), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n316), .A2(new_n209), .A3(G68), .A4(new_n267), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT19), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n522), .A2(new_n209), .A3(G33), .A4(G97), .ZN(new_n523));
  NOR2_X1   g0323(.A1(G87), .A2(G97), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n524), .A2(new_n220), .B1(new_n412), .B2(new_n209), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n523), .B1(new_n525), .B2(new_n522), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n520), .B1(new_n527), .B2(new_n261), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n208), .A2(G33), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n258), .A2(new_n529), .A3(new_n234), .A4(new_n260), .ZN(new_n530));
  OR3_X1    g0330(.A1(new_n530), .A2(KEYINPUT79), .A3(new_n432), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT79), .B1(new_n530), .B2(new_n432), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT80), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n528), .A2(new_n533), .A3(KEYINPUT80), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G244), .A2(G1698), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n442), .B2(G1698), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n267), .B(new_n539), .C1(new_n269), .C2(new_n270), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n268), .A2(new_n459), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n305), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(G45), .ZN(new_n544));
  OAI21_X1  g0344(.A(G250), .B1(new_n544), .B2(G1), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n208), .A2(G45), .A3(G274), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n305), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n340), .B1(new_n543), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n541), .B1(new_n278), .B2(new_n539), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n338), .B(new_n548), .C1(new_n551), .C2(new_n305), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n536), .A2(new_n537), .A3(new_n554), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n290), .A2(G107), .A3(new_n293), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT6), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n557), .A2(G97), .A3(G107), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n215), .A2(KEYINPUT6), .ZN(new_n559));
  NOR2_X1   g0359(.A1(KEYINPUT77), .A2(G107), .ZN(new_n560));
  NAND2_X1  g0360(.A1(KEYINPUT77), .A2(G107), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n558), .A2(new_n559), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n215), .A2(new_n220), .A3(KEYINPUT6), .ZN(new_n564));
  OR2_X1    g0364(.A1(KEYINPUT77), .A2(G107), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n557), .A2(G97), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .A4(new_n561), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n563), .A2(G20), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n282), .A2(G77), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n261), .B1(new_n556), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n259), .A2(G97), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(G97), .B2(new_n530), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n370), .A2(G244), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT4), .B1(new_n278), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n291), .A2(new_n267), .A3(G250), .A4(G1698), .ZN(new_n577));
  AND2_X1   g0377(.A1(KEYINPUT4), .A2(G244), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n291), .A2(new_n267), .A3(new_n578), .A4(new_n370), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(new_n579), .A3(new_n470), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n320), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G257), .B(new_n305), .C1(new_n488), .C2(new_n490), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n497), .A2(new_n493), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n581), .A2(new_n299), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(G200), .B1(new_n581), .B2(new_n585), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n571), .B(new_n574), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n581), .A2(G179), .A3(new_n585), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n340), .B1(new_n581), .B2(new_n585), .ZN(new_n590));
  INV_X1    g0390(.A(new_n261), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n568), .A2(new_n569), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n290), .A2(G107), .A3(new_n293), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI22_X1  g0394(.A1(new_n589), .A2(new_n590), .B1(new_n594), .B2(new_n573), .ZN(new_n595));
  OAI21_X1  g0395(.A(G200), .B1(new_n543), .B2(new_n549), .ZN(new_n596));
  INV_X1    g0396(.A(new_n530), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G87), .ZN(new_n598));
  OAI211_X1 g0398(.A(G190), .B(new_n548), .C1(new_n551), .C2(new_n305), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n596), .A2(new_n528), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n555), .A2(new_n588), .A3(new_n595), .A4(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT22), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(new_n213), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n316), .A2(new_n209), .A3(new_n267), .A4(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n213), .A2(G20), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n602), .B1(new_n292), .B2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(KEYINPUT84), .B(KEYINPUT23), .C1(new_n209), .C2(G107), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT23), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT84), .B1(new_n209), .B2(G107), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n609), .A2(new_n610), .B1(new_n541), .B2(new_n209), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n604), .A2(new_n607), .A3(new_n608), .A4(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT24), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n610), .A2(new_n609), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n541), .A2(new_n209), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n615), .A2(new_n616), .A3(new_n608), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n617), .A2(KEYINPUT24), .A3(new_n604), .A4(new_n607), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n614), .A2(new_n261), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n397), .A2(G20), .A3(new_n220), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT25), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(G107), .B2(new_n597), .ZN(new_n622));
  OAI211_X1 g0422(.A(G264), .B(new_n305), .C1(new_n488), .C2(new_n490), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(G257), .A2(G1698), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n214), .B2(G1698), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n267), .B(new_n626), .C1(new_n269), .C2(new_n270), .ZN(new_n627));
  INV_X1    g0427(.A(G294), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n268), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n624), .B1(new_n631), .B2(new_n320), .ZN(new_n632));
  AOI21_X1  g0432(.A(G200), .B1(new_n632), .B2(new_n500), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n629), .B1(new_n278), .B2(new_n626), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n500), .B(new_n623), .C1(new_n634), .C2(new_n305), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(G190), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n619), .B(new_n622), .C1(new_n633), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n618), .A2(new_n261), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n615), .A2(new_n616), .A3(new_n608), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT22), .B1(new_n368), .B2(new_n605), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT24), .B1(new_n641), .B2(new_n604), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n622), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n635), .A2(G169), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n631), .A2(new_n320), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n645), .A2(G179), .A3(new_n500), .A4(new_n623), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT85), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n637), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n637), .A2(new_n648), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT85), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n601), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n458), .A2(new_n519), .A3(new_n653), .ZN(G372));
  NAND2_X1  g0454(.A1(new_n554), .A2(new_n534), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n637), .A2(new_n655), .A3(new_n600), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n588), .A2(new_n595), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n648), .B(new_n504), .C1(KEYINPUT21), .C2(new_n510), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n531), .A2(new_n532), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n591), .B1(new_n521), .B2(new_n526), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n660), .A2(new_n661), .A3(new_n520), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n553), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n596), .A2(new_n599), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n527), .A2(new_n261), .ZN(new_n665));
  INV_X1    g0465(.A(new_n520), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n666), .A3(new_n598), .ZN(new_n667));
  OAI22_X1  g0467(.A1(new_n662), .A2(new_n553), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n595), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n663), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n590), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n581), .A2(G179), .A3(new_n585), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n672), .A2(new_n673), .B1(new_n571), .B2(new_n574), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(new_n555), .A3(new_n600), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT26), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n659), .A2(new_n671), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n458), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n330), .A2(new_n336), .ZN(new_n679));
  INV_X1    g0479(.A(new_n431), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n448), .B1(new_n456), .B2(new_n454), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n344), .A2(new_n347), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI22_X1  g0484(.A1(new_n684), .A2(new_n390), .B1(new_n365), .B2(new_n392), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n678), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT86), .ZN(G369));
  OR3_X1    g0487(.A1(new_n462), .A2(KEYINPUT27), .A3(G20), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT27), .B1(new_n462), .B2(G20), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G213), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G343), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n512), .A2(new_n518), .B1(new_n481), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n516), .A2(new_n504), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n481), .A2(new_n692), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OR3_X1    g0496(.A1(new_n693), .A2(new_n696), .A3(KEYINPUT87), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT87), .B1(new_n693), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n652), .A2(new_n650), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n643), .A2(new_n692), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n692), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n648), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT88), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n701), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n648), .A2(new_n692), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n694), .A2(new_n692), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n710), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n709), .A2(new_n712), .ZN(G399));
  NOR2_X1   g0513(.A1(new_n227), .A2(G41), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR4_X1   g0515(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(G1), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n232), .B2(new_n715), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n677), .A2(new_n705), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n672), .A2(new_n673), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n571), .A2(new_n574), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n655), .A2(new_n723), .A3(new_n724), .A4(new_n600), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n655), .A2(KEYINPUT92), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT92), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n663), .A2(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n725), .A2(KEYINPUT26), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n674), .A2(new_n555), .A3(new_n670), .A4(new_n600), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n659), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(KEYINPUT29), .A3(new_n705), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n722), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n653), .A2(new_n519), .A3(new_n705), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n705), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT89), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(new_n505), .B2(G179), .ZN(new_n739));
  NOR4_X1   g0539(.A1(new_n486), .A2(new_n498), .A3(KEYINPUT89), .A4(new_n338), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n543), .A2(new_n549), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(new_n632), .A3(new_n581), .A4(new_n585), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n737), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n505), .A2(new_n742), .A3(G179), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT90), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n316), .A2(new_n267), .A3(new_n575), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT4), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n577), .A2(new_n579), .A3(new_n470), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n305), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n500), .A2(new_n582), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n746), .B(new_n635), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n581), .A2(new_n585), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n746), .B1(new_n755), .B2(new_n635), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n745), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n744), .A2(KEYINPUT91), .A3(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n741), .A2(new_n737), .A3(new_n743), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(KEYINPUT91), .B1(new_n744), .B2(new_n757), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n736), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n744), .A2(new_n757), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n692), .B1(new_n764), .B2(new_n759), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n735), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n734), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G330), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n733), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n719), .B1(new_n769), .B2(G1), .ZN(G364));
  NOR2_X1   g0570(.A1(new_n396), .A2(G20), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G45), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n715), .A2(G1), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n701), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G330), .B2(new_n699), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n774), .A2(KEYINPUT93), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n774), .A2(KEYINPUT93), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n234), .B1(G20), .B2(new_n340), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n209), .A2(G190), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G179), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G329), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n292), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n325), .A2(G179), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n787), .A2(G20), .A3(G190), .ZN(new_n791));
  INV_X1    g0591(.A(G303), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n789), .A2(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n783), .A2(G190), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G20), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n786), .B(new_n793), .C1(G294), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(G20), .A2(G179), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT96), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n299), .A2(new_n325), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(KEYINPUT98), .B(G326), .Z(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n299), .A2(G200), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n798), .A2(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n801), .A2(new_n803), .B1(new_n805), .B2(G322), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n796), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n798), .A2(new_n299), .A3(new_n325), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n798), .A2(new_n299), .A3(G200), .ZN(new_n810));
  XOR2_X1   g0610(.A(KEYINPUT33), .B(G317), .Z(new_n811));
  OAI221_X1 g0611(.A(new_n807), .B1(new_n808), .B2(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G159), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n784), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT32), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n788), .A2(G107), .ZN(new_n816));
  INV_X1    g0616(.A(new_n791), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G87), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n815), .A2(new_n368), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n805), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n820), .A2(new_n202), .B1(new_n362), .B2(new_n800), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n795), .A2(G97), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n810), .B2(new_n203), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT97), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n822), .B(new_n825), .C1(new_n372), .C2(new_n809), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n781), .B1(new_n812), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(G13), .A2(G33), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(G20), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n780), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT95), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n227), .A2(new_n459), .ZN(new_n834));
  XNOR2_X1  g0634(.A(G355), .B(KEYINPUT94), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n226), .A2(new_n368), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n233), .A2(G45), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n249), .B2(G45), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n227), .A2(new_n278), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n834), .B1(new_n835), .B2(new_n836), .C1(new_n838), .C2(new_n840), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n779), .B(new_n827), .C1(new_n833), .C2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n830), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n699), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n776), .A2(new_n844), .ZN(G396));
  NOR2_X1   g0645(.A1(new_n780), .A2(new_n828), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n779), .B1(new_n372), .B2(new_n846), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n820), .A2(new_n628), .B1(new_n792), .B2(new_n800), .ZN(new_n848));
  INV_X1    g0648(.A(new_n784), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n368), .B1(new_n849), .B2(G311), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n817), .A2(G107), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n788), .A2(G87), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n850), .A2(new_n851), .A3(new_n823), .A4(new_n852), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n459), .A2(new_n809), .B1(new_n810), .B2(new_n790), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n848), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(G137), .A2(new_n801), .B1(new_n805), .B2(G143), .ZN(new_n856));
  INV_X1    g0656(.A(G150), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n856), .B1(new_n857), .B2(new_n810), .C1(new_n813), .C2(new_n809), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT34), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n788), .A2(G68), .ZN(new_n860));
  INV_X1    g0660(.A(G132), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n860), .B1(new_n362), .B2(new_n791), .C1(new_n861), .C2(new_n784), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n271), .B(new_n862), .C1(G58), .C2(new_n795), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n855), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n451), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n439), .B1(new_n865), .B2(new_n449), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n439), .A2(new_n692), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n448), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n448), .A2(new_n692), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n847), .B1(new_n864), .B2(new_n781), .C1(new_n829), .C2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n677), .A2(new_n705), .A3(new_n870), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT99), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT99), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n677), .A2(new_n874), .A3(new_n705), .A4(new_n870), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n677), .A2(new_n705), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n877), .B2(new_n870), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n878), .A2(new_n768), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n773), .B1(new_n878), .B2(new_n768), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n871), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT100), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(G384));
  AOI211_X1 g0683(.A(new_n372), .B(new_n232), .C1(G58), .C2(G68), .ZN(new_n884));
  INV_X1    g0684(.A(new_n201), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n885), .A2(new_n203), .ZN(new_n886));
  OAI211_X1 g0686(.A(G1), .B(new_n396), .C1(new_n884), .C2(new_n886), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT101), .Z(new_n888));
  NAND3_X1  g0688(.A1(new_n235), .A2(G20), .A3(G116), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n563), .A2(new_n567), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT35), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n891), .B2(new_n890), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT36), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n888), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n894), .B2(new_n893), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT16), .B1(new_n280), .B2(new_n283), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n333), .A2(new_n897), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n898), .A2(new_n264), .B1(new_n342), .B2(new_n690), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n324), .A2(new_n343), .A3(new_n264), .A4(new_n329), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT37), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT104), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n335), .A2(new_n346), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n903), .B1(new_n335), .B2(new_n346), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n690), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n335), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT37), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n900), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n902), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n690), .B1(new_n898), .B2(new_n264), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n912), .B1(new_n354), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(KEYINPUT38), .B(new_n912), .C1(new_n354), .C2(new_n914), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT103), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n876), .A2(new_n869), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n431), .A2(KEYINPUT102), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT102), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n923), .B(new_n409), .C1(new_n426), .C2(new_n430), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n456), .A2(new_n454), .B1(new_n409), .B2(new_n692), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n680), .A2(new_n692), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n920), .B1(new_n921), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n869), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n873), .B2(new_n875), .ZN(new_n931));
  INV_X1    g0731(.A(new_n928), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n931), .A2(KEYINPUT103), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n919), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n344), .A2(new_n347), .A3(KEYINPUT75), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n351), .B1(new_n350), .B2(new_n352), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n679), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n913), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT38), .B1(new_n938), .B2(new_n912), .ZN(new_n939));
  INV_X1    g0739(.A(new_n918), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT39), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n909), .B1(new_n679), .B2(new_n683), .ZN(new_n942));
  INV_X1    g0742(.A(new_n906), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n904), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n900), .A2(new_n909), .A3(new_n910), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n900), .A2(new_n349), .A3(new_n909), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n944), .A2(new_n945), .B1(KEYINPUT37), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n916), .B1(new_n942), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n918), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n941), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n692), .B1(new_n922), .B2(new_n924), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n683), .A2(new_n908), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n934), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n458), .A2(new_n732), .A3(new_n722), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n957), .A2(new_n685), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n956), .B(new_n958), .Z(new_n959));
  OAI211_X1 g0759(.A(KEYINPUT31), .B(new_n692), .C1(new_n764), .C2(new_n759), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n734), .A2(new_n766), .A3(new_n960), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n961), .A2(new_n870), .A3(new_n928), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n939), .B2(new_n940), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT40), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n918), .A2(new_n948), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n962), .A2(new_n966), .A3(KEYINPUT40), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n458), .A2(new_n961), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT105), .Z(new_n970));
  OR2_X1    g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n968), .A2(new_n970), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(G330), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n959), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n208), .B2(new_n771), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n959), .A2(new_n973), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n896), .B1(new_n975), .B2(new_n976), .ZN(G367));
  AOI21_X1  g0777(.A(new_n832), .B1(new_n227), .B2(new_n433), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n839), .A2(new_n245), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n779), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n667), .A2(new_n692), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n663), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n668), .B2(new_n981), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n791), .A2(new_n459), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(KEYINPUT46), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT110), .Z(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(KEYINPUT46), .B2(new_n984), .C1(new_n628), .C2(new_n810), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n987), .A2(KEYINPUT111), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(KEYINPUT111), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n849), .A2(G317), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n788), .A2(G97), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n795), .A2(G107), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n990), .A2(new_n991), .A3(new_n271), .A4(new_n992), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n820), .A2(new_n792), .B1(new_n808), .B2(new_n800), .ZN(new_n994));
  INV_X1    g0794(.A(new_n809), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n993), .B(new_n994), .C1(G283), .C2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n988), .A2(new_n989), .A3(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT112), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n817), .A2(G58), .B1(new_n849), .B2(G137), .ZN(new_n999));
  INV_X1    g0799(.A(new_n795), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n999), .B1(new_n203), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n368), .B1(new_n789), .B2(new_n372), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1001), .B1(KEYINPUT113), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n813), .B2(new_n810), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n885), .B2(new_n995), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G143), .A2(new_n801), .B1(new_n805), .B2(G150), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(KEYINPUT113), .C2(new_n1002), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n998), .A2(KEYINPUT47), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n780), .ZN(new_n1009));
  AOI21_X1  g0809(.A(KEYINPUT47), .B1(new_n998), .B2(new_n1007), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n980), .B1(new_n843), .B2(new_n983), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n772), .A2(G1), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n724), .A2(new_n692), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n657), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n674), .A2(new_n692), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n712), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT44), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT45), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT107), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n712), .A2(new_n1020), .A3(new_n1016), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1020), .B1(new_n712), .B2(new_n1016), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1019), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1023), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1025), .A2(KEYINPUT45), .A3(new_n1021), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1018), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n708), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n700), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(KEYINPUT108), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT108), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1027), .A2(new_n1032), .A3(new_n1029), .ZN(new_n1033));
  AND4_X1   g0833(.A1(new_n709), .A2(new_n1018), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n708), .B1(new_n699), .B2(G330), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n709), .A2(new_n711), .A3(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1029), .A2(new_n1037), .B1(new_n694), .B2(new_n692), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n1040), .A3(new_n769), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT109), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1039), .A2(new_n1040), .A3(KEYINPUT109), .A4(new_n769), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n769), .B1(new_n1036), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n714), .B(KEYINPUT41), .Z(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1012), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1016), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n709), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n708), .A2(new_n711), .A3(new_n1016), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1052), .A2(KEYINPUT42), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(KEYINPUT42), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n595), .B1(new_n1014), .B2(new_n648), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n705), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .A4(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1053), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n983), .B(KEYINPUT43), .Z(new_n1060));
  AOI22_X1  g0860(.A1(new_n1058), .A2(KEYINPUT106), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1058), .A2(KEYINPUT106), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n1051), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1051), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1011), .B1(new_n1049), .B2(new_n1066), .ZN(G387));
  NAND2_X1  g0867(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n769), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n715), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1045), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1012), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n779), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n836), .A2(new_n716), .B1(G107), .B2(new_n226), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n356), .A2(new_n362), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT50), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n716), .B(new_n544), .C1(new_n203), .C2(new_n372), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n839), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT114), .Z(new_n1080));
  NAND2_X1  g0880(.A1(new_n242), .A2(G45), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1075), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1074), .B1(new_n1082), .B2(new_n832), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n991), .B1(new_n372), .B2(new_n791), .C1(new_n857), .C2(new_n784), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1000), .A2(new_n432), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n1084), .A2(new_n271), .A3(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G159), .A2(new_n801), .B1(new_n805), .B2(G50), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n810), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G68), .A2(new_n995), .B1(new_n1088), .B2(new_n356), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1086), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G322), .A2(new_n801), .B1(new_n805), .B2(G317), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1091), .B1(new_n792), .B2(new_n809), .C1(new_n808), .C2(new_n810), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT48), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n817), .A2(G294), .B1(new_n795), .B2(G283), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT49), .Z(new_n1098));
  AOI22_X1  g0898(.A1(new_n803), .A2(new_n849), .B1(new_n788), .B2(G116), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n271), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1090), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1083), .B1(new_n1101), .B2(new_n780), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n708), .B2(new_n843), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT115), .Z(new_n1104));
  NOR2_X1   g0904(.A1(new_n1073), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1071), .A2(new_n1105), .ZN(G393));
  NAND3_X1  g0906(.A1(new_n1035), .A2(new_n1030), .A3(new_n1012), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n833), .B1(new_n215), .B2(new_n226), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n840), .A2(new_n252), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1074), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n817), .A2(G283), .B1(new_n849), .B2(G322), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1111), .A2(new_n292), .A3(new_n816), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G116), .B2(new_n795), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n628), .B2(new_n809), .C1(new_n792), .C2(new_n810), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G317), .A2(new_n801), .B1(new_n805), .B2(G311), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT52), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n852), .B1(new_n203), .B2(new_n791), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1000), .A2(new_n372), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n849), .A2(G143), .ZN(new_n1119));
  NOR4_X1   g0919(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .A4(new_n271), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n201), .B2(new_n810), .C1(new_n254), .C2(new_n809), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(G150), .A2(new_n801), .B1(new_n805), .B2(G159), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT51), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n1114), .A2(new_n1116), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1110), .B1(new_n1124), .B2(new_n780), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n1016), .B2(new_n843), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1107), .A2(new_n1126), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n715), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1035), .A2(new_n1030), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1045), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1127), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(G390));
  NAND3_X1  g0934(.A1(new_n961), .A2(G330), .A3(new_n870), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n932), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n731), .A2(new_n705), .A3(new_n868), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n869), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n767), .A2(new_n928), .A3(G330), .A4(new_n870), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1136), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n767), .A2(G330), .A3(new_n870), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n932), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n961), .A2(new_n928), .A3(G330), .A4(new_n870), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1141), .B1(new_n1145), .B2(new_n931), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n458), .A2(G330), .A3(new_n961), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n957), .A2(new_n1147), .A3(new_n685), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT116), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n952), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n931), .B2(new_n932), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1151), .A2(new_n941), .A3(new_n950), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n952), .B1(new_n1138), .B2(new_n928), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n966), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1152), .A2(new_n1154), .A3(new_n1140), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1144), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1149), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1144), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1136), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n931), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1148), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT116), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1152), .A2(new_n1154), .A3(new_n1140), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1160), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1157), .A2(new_n1167), .A3(new_n714), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n779), .B1(new_n254), .B2(new_n846), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n820), .A2(new_n459), .B1(new_n790), .B2(new_n800), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n215), .A2(new_n809), .B1(new_n810), .B2(new_n220), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n849), .A2(G294), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n818), .A2(new_n1172), .A3(new_n292), .A4(new_n860), .ZN(new_n1173));
  NOR4_X1   g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1118), .A4(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n292), .B1(new_n788), .B2(new_n885), .ZN(new_n1175));
  INV_X1    g0975(.A(G125), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1175), .B1(new_n1176), .B2(new_n784), .C1(new_n813), .C2(new_n1000), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n791), .A2(new_n857), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT53), .ZN(new_n1179));
  INV_X1    g0979(.A(G128), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1179), .B1(new_n1180), .B2(new_n800), .C1(new_n861), .C2(new_n820), .ZN(new_n1181));
  XOR2_X1   g0981(.A(KEYINPUT54), .B(G143), .Z(new_n1182));
  AOI22_X1  g0982(.A1(G137), .A2(new_n1088), .B1(new_n995), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1177), .B(new_n1181), .C1(KEYINPUT117), .C2(new_n1184), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1184), .A2(KEYINPUT117), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1174), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1169), .B1(new_n1187), .B2(new_n781), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n949), .B1(new_n917), .B2(new_n918), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n950), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1188), .B1(new_n1191), .B2(new_n828), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(new_n1012), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1168), .A2(new_n1194), .ZN(G378));
  INV_X1    g0995(.A(new_n846), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n774), .B1(new_n885), .B2(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n805), .A2(G128), .B1(new_n817), .B2(new_n1182), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT119), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n995), .A2(G137), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n810), .A2(new_n861), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n800), .A2(new_n1176), .B1(new_n1000), .B2(new_n857), .ZN(new_n1202));
  NOR4_X1   g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT59), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n849), .A2(G124), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n268), .B(new_n487), .C1(new_n789), .C2(new_n813), .ZN(new_n1208));
  NOR4_X1   g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n271), .A2(new_n487), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n788), .A2(G58), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n372), .B2(new_n791), .C1(new_n790), .C2(new_n784), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1210), .B(new_n1212), .C1(G107), .C2(new_n805), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n800), .A2(new_n459), .B1(new_n1000), .B2(new_n203), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT118), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G97), .A2(new_n1088), .B1(new_n995), .B2(new_n433), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1213), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1217), .A2(KEYINPUT58), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(KEYINPUT58), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1210), .B(new_n362), .C1(G33), .C2(G41), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n780), .B1(new_n1209), .B2(new_n1221), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT120), .Z(new_n1223));
  AND3_X1   g1023(.A1(new_n394), .A2(new_n365), .A3(new_n908), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n394), .B1(new_n365), .B2(new_n908), .ZN(new_n1225));
  XOR2_X1   g1025(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1226));
  OR3_X1    g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1226), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1197), .B(new_n1223), .C1(new_n828), .C2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n961), .A2(new_n928), .A3(new_n870), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n917), .B2(new_n918), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n967), .B(G330), .C1(new_n1233), .C2(KEYINPUT40), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1230), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n965), .A2(G330), .A3(new_n967), .A4(new_n1229), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n956), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n954), .B1(new_n951), .B2(new_n952), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1235), .A2(new_n1239), .A3(new_n1236), .A4(new_n934), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1231), .B1(new_n1241), .B2(new_n1012), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1191), .A2(new_n1151), .B1(new_n966), .B2(new_n1153), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1166), .B(new_n1146), .C1(new_n1244), .C2(new_n1144), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1148), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1241), .A2(new_n1246), .A3(KEYINPUT121), .A4(KEYINPUT57), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n714), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1241), .A2(new_n1246), .A3(KEYINPUT57), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT57), .B1(new_n1241), .B2(new_n1246), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT121), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1250), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1243), .B1(new_n1249), .B2(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT122), .ZN(G375));
  NOR2_X1   g1055(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n928), .A2(new_n829), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n801), .A2(G132), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT123), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1088), .A2(new_n1182), .B1(new_n805), .B2(G137), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(KEYINPUT124), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n809), .A2(new_n857), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1211), .B1(new_n1180), .B2(new_n784), .C1(new_n813), .C2(new_n791), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n278), .B1(new_n1000), .B2(new_n362), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n820), .A2(new_n790), .B1(new_n628), .B2(new_n800), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n368), .B1(new_n788), .B2(G77), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1268), .B1(new_n215), .B2(new_n791), .C1(new_n792), .C2(new_n784), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n220), .A2(new_n809), .B1(new_n810), .B2(new_n459), .ZN(new_n1270));
  NOR4_X1   g1070(.A1(new_n1267), .A2(new_n1269), .A3(new_n1270), .A4(new_n1085), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n780), .B1(new_n1266), .B2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1272), .B(new_n1074), .C1(G68), .C2(new_n1196), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n1256), .A2(new_n1072), .B1(new_n1257), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1148), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1256), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(new_n1048), .A3(new_n1163), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(G381));
  INV_X1    g1079(.A(KEYINPUT125), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G378), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1168), .A2(new_n1194), .A3(KEYINPUT125), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(G375), .A2(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(G387), .A2(G390), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(G393), .A2(G396), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(G384), .A2(G381), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1284), .A2(new_n1285), .A3(new_n1286), .A4(new_n1287), .ZN(G407));
  NAND3_X1  g1088(.A1(new_n1284), .A2(G213), .A3(new_n691), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(G407), .A2(new_n1289), .A3(G213), .ZN(G409));
  NAND2_X1  g1090(.A1(new_n691), .A2(G213), .ZN(new_n1291));
  XOR2_X1   g1091(.A(new_n1277), .B(KEYINPUT60), .Z(new_n1292));
  INV_X1    g1092(.A(new_n1163), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1292), .A2(new_n715), .A3(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n882), .B1(new_n1294), .B2(new_n1274), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1163), .A2(new_n714), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G384), .B(new_n1275), .C1(new_n1292), .C2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1241), .A2(new_n1246), .A3(new_n1048), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1242), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1281), .A2(new_n1301), .A3(new_n1282), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(KEYINPUT126), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1281), .A2(new_n1301), .A3(new_n1304), .A4(new_n1282), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(G378), .ZN(new_n1307));
  AOI211_X1 g1107(.A(new_n1307), .B(new_n1243), .C1(new_n1249), .C2(new_n1253), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1291), .B(new_n1299), .C1(new_n1306), .C2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(KEYINPUT62), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1291), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n691), .A2(G213), .A3(G2897), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1295), .A2(new_n1297), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1312), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1311), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT61), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1253), .ZN(new_n1318));
  OAI211_X1 g1118(.A(G378), .B(new_n1242), .C1(new_n1318), .C2(new_n1248), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1319), .A2(new_n1303), .A3(new_n1305), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1320), .A2(new_n1321), .A3(new_n1291), .A4(new_n1299), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1310), .A2(new_n1316), .A3(new_n1317), .A4(new_n1322), .ZN(new_n1323));
  AOI22_X1  g1123(.A1(new_n1071), .A2(new_n1105), .B1(new_n776), .B2(new_n844), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1286), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT127), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1034), .B1(KEYINPUT108), .B2(new_n1030), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1327), .A2(new_n1043), .A3(new_n1044), .A4(new_n1033), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1047), .B1(new_n1328), .B2(new_n769), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1065), .B1(new_n1329), .B2(new_n1012), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1133), .B1(new_n1330), .B2(new_n1011), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1325), .B(new_n1326), .C1(new_n1285), .C2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(G387), .A2(G390), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1330), .A2(new_n1011), .A3(new_n1133), .ZN(new_n1335));
  OAI21_X1  g1135(.A(KEYINPUT127), .B1(new_n1286), .B2(new_n1324), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1333), .A2(new_n1334), .A3(new_n1335), .A4(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1332), .A2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1323), .A2(new_n1338), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1332), .A2(new_n1317), .A3(new_n1337), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1320), .A2(KEYINPUT63), .A3(new_n1291), .A4(new_n1299), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT63), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1342), .B1(new_n1311), .B2(new_n1315), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1309), .ZN(new_n1344));
  OAI211_X1 g1144(.A(new_n1340), .B(new_n1341), .C1(new_n1343), .C2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1339), .A2(new_n1345), .ZN(G405));
  NAND3_X1  g1146(.A1(G375), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(new_n1319), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1299), .B1(new_n1332), .B2(new_n1337), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1332), .A2(new_n1337), .A3(new_n1299), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1348), .A2(new_n1350), .A3(new_n1351), .ZN(new_n1352));
  AND3_X1   g1152(.A1(new_n1332), .A2(new_n1337), .A3(new_n1299), .ZN(new_n1353));
  OAI211_X1 g1153(.A(new_n1319), .B(new_n1347), .C1(new_n1353), .C2(new_n1349), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1352), .A2(new_n1354), .ZN(G402));
endmodule


