//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n567, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n451), .B(new_n452), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OR2_X1    g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n466), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  NOR2_X1   g049(.A1(new_n464), .A2(new_n465), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(new_n467), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n479));
  INV_X1    g054(.A(G136), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n477), .B(new_n479), .C1(new_n480), .C2(new_n468), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  NAND3_X1  g057(.A1(new_n466), .A2(G138), .A3(new_n467), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n484), .A2(KEYINPUT68), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(KEYINPUT68), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(G126), .B1(new_n464), .B2(new_n465), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n467), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n483), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n466), .A2(KEYINPUT4), .A3(G138), .ZN(new_n493));
  NAND2_X1  g068(.A1(G102), .A2(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(new_n467), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n492), .A2(new_n497), .ZN(G164));
  OR2_X1    g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OR2_X1    g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(G543), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n501), .A2(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT69), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n511), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  AOI22_X1  g093(.A1(new_n499), .A2(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n519), .A2(G89), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n510), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g101(.A(KEYINPUT70), .B(G543), .C1(new_n508), .C2(new_n509), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(new_n526), .B2(new_n527), .ZN(new_n534));
  INV_X1    g109(.A(new_n531), .ZN(new_n535));
  OAI21_X1  g110(.A(KEYINPUT71), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n524), .B1(new_n532), .B2(new_n536), .ZN(G168));
  NAND2_X1  g112(.A1(new_n528), .A2(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  AND2_X1   g114(.A1(KEYINPUT5), .A2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(KEYINPUT5), .A2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n544), .A2(G651), .B1(new_n519), .B2(G90), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n538), .A2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  NAND3_X1  g122(.A1(new_n501), .A2(new_n504), .A3(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n501), .B2(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n548), .B1(new_n551), .B2(new_n512), .ZN(new_n552));
  INV_X1    g127(.A(G43), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n526), .B2(new_n527), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT72), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n549), .B1(new_n542), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n557), .A2(G651), .B1(new_n519), .B2(G81), .ZN(new_n558));
  AOI21_X1  g133(.A(KEYINPUT70), .B1(new_n504), .B2(G543), .ZN(new_n559));
  INV_X1    g134(.A(new_n527), .ZN(new_n560));
  OAI21_X1  g135(.A(G43), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n558), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n555), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(new_n569));
  XOR2_X1   g144(.A(new_n569), .B(KEYINPUT73), .Z(G188));
  XNOR2_X1  g145(.A(new_n542), .B(KEYINPUT74), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g148(.A1(G78), .A2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n502), .B2(new_n503), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G53), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(KEYINPUT9), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(KEYINPUT9), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n579), .A2(new_n580), .B1(G91), .B2(new_n519), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n575), .A2(new_n581), .ZN(G299));
  NAND2_X1  g157(.A1(new_n532), .A2(new_n536), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(new_n523), .ZN(G286));
  OAI21_X1  g159(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n577), .A2(G49), .ZN(new_n586));
  INV_X1    g161(.A(G87), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n585), .B(new_n586), .C1(new_n587), .C2(new_n505), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT75), .ZN(G288));
  NAND2_X1  g164(.A1(new_n519), .A2(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n577), .A2(G48), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n501), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n512), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n592), .A2(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(new_n528), .A2(G47), .ZN(new_n596));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n542), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(new_n519), .B2(G85), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n571), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g179(.A1(G79), .A2(G543), .ZN(new_n605));
  OAI21_X1  g180(.A(G651), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n528), .A2(G54), .ZN(new_n607));
  AND3_X1   g182(.A1(new_n501), .A2(new_n504), .A3(G92), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT10), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n602), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n602), .B1(new_n611), .B2(G868), .ZN(G321));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(G299), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n614), .B2(G168), .ZN(G297));
  OAI21_X1  g191(.A(new_n615), .B1(new_n614), .B2(G168), .ZN(G280));
  INV_X1    g192(.A(G860), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n610), .B1(G559), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT76), .ZN(G148));
  NAND2_X1  g195(.A1(new_n555), .A2(new_n563), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(new_n614), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n610), .A2(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n614), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n466), .A2(new_n462), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT77), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  INV_X1    g207(.A(new_n468), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n633), .A2(G135), .B1(G123), .B2(new_n476), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  INV_X1    g210(.A(G111), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n635), .A2(KEYINPUT78), .B1(new_n636), .B2(G2105), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(KEYINPUT78), .B2(new_n635), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n631), .A2(new_n632), .A3(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT79), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT80), .ZN(new_n656));
  OAI21_X1  g231(.A(G14), .B1(new_n653), .B2(new_n654), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT17), .Z(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  INV_X1    g239(.A(new_n661), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(new_n659), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n663), .B(new_n664), .C1(new_n662), .C2(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n659), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT18), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT81), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n675), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n675), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(G229));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G33), .ZN(new_n692));
  NAND2_X1  g267(.A1(G115), .A2(G2104), .ZN(new_n693));
  INV_X1    g268(.A(G127), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n475), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n467), .B1(new_n695), .B2(KEYINPUT88), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(KEYINPUT88), .B2(new_n695), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT25), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n633), .B2(G139), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT89), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT90), .Z(new_n704));
  OAI21_X1  g279(.A(new_n692), .B1(new_n704), .B2(new_n691), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(G2072), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT91), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT82), .B(G29), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(G27), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G164), .B2(new_n709), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(G2078), .Z(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G20), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT23), .Z(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G299), .B2(G16), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT96), .B(G1956), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n712), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT24), .B(G34), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n708), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT92), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G160), .B2(G29), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(G2084), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT94), .Z(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT31), .B(G11), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT93), .B(G28), .Z(new_n727));
  AOI21_X1  g302(.A(G29), .B1(new_n727), .B2(KEYINPUT30), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(KEYINPUT30), .B2(new_n727), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n726), .B(new_n729), .C1(new_n639), .C2(new_n708), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n723), .B2(G2084), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n691), .A2(G32), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n633), .A2(G141), .B1(G105), .B2(new_n462), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n476), .A2(G129), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT26), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n732), .B1(new_n739), .B2(new_n691), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G1996), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n725), .A2(new_n731), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n713), .A2(G5), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G171), .B2(new_n713), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(G1961), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n709), .A2(G35), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G162), .B2(new_n709), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n749));
  INV_X1    g324(.A(G2090), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n748), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n745), .A2(G1961), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR4_X1   g329(.A1(new_n719), .A2(new_n743), .A3(new_n746), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n705), .A2(G2072), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n713), .A2(G21), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G168), .B2(new_n713), .ZN(new_n758));
  INV_X1    g333(.A(G1966), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  AND3_X1   g335(.A1(new_n755), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G4), .A2(G16), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n611), .B2(G16), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT85), .B(G1348), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n708), .A2(G26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n476), .A2(G128), .ZN(new_n768));
  INV_X1    g343(.A(G140), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(new_n468), .ZN(new_n770));
  OAI21_X1  g345(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n771));
  INV_X1    g346(.A(G116), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G2105), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT86), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n767), .B1(new_n775), .B2(new_n691), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2067), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n713), .A2(G19), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n564), .B2(new_n713), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n777), .B1(G1341), .B2(new_n779), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n765), .B(new_n780), .C1(G1341), .C2(new_n779), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT87), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n707), .A2(new_n761), .A3(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(KEYINPUT97), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(KEYINPUT97), .ZN(new_n785));
  MUX2_X1   g360(.A(G23), .B(new_n588), .S(G16), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT33), .ZN(new_n787));
  INV_X1    g362(.A(G1976), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n713), .A2(G22), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT83), .Z(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G166), .B2(new_n713), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1971), .ZN(new_n793));
  NOR2_X1   g368(.A1(G6), .A2(G16), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n592), .A2(new_n594), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT32), .B(G1981), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  OR3_X1    g373(.A1(new_n789), .A2(new_n793), .A3(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(KEYINPUT34), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(KEYINPUT34), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n709), .A2(G25), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n633), .A2(G131), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n476), .A2(G119), .ZN(new_n804));
  OR2_X1    g379(.A1(G95), .A2(G2105), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n805), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n802), .B1(new_n808), .B2(new_n709), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT35), .B(G1991), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G1986), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n713), .A2(G24), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G290), .B2(G16), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n811), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n812), .B2(new_n814), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n800), .A2(new_n801), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(KEYINPUT84), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n817), .B(new_n819), .Z(new_n820));
  OR2_X1    g395(.A1(new_n818), .A2(KEYINPUT84), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n784), .A2(new_n785), .B1(new_n820), .B2(new_n821), .ZN(G311));
  NAND2_X1  g397(.A1(new_n784), .A2(new_n785), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n820), .A2(new_n821), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(G150));
  NAND2_X1  g400(.A1(G80), .A2(G543), .ZN(new_n826));
  INV_X1    g401(.A(G67), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n542), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G651), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT99), .ZN(new_n830));
  OAI21_X1  g405(.A(G55), .B1(new_n559), .B2(new_n560), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT98), .B(G93), .Z(new_n832));
  AND3_X1   g407(.A1(new_n832), .A2(new_n501), .A3(new_n504), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n830), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(G55), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n526), .B2(new_n527), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n837), .A2(KEYINPUT99), .A3(new_n833), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n829), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G860), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT101), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n611), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n558), .A2(new_n561), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n845), .B(new_n829), .C1(new_n835), .C2(new_n838), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n831), .A2(new_n834), .A3(new_n830), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT99), .B1(new_n837), .B2(new_n833), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n848), .A2(new_n849), .B1(G651), .B2(new_n828), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n846), .B(new_n847), .C1(new_n621), .C2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n839), .A2(new_n564), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n847), .B1(new_n853), .B2(new_n846), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n844), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n618), .B1(new_n857), .B2(KEYINPUT39), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n842), .B1(new_n858), .B2(new_n859), .ZN(G145));
  XNOR2_X1  g435(.A(G164), .B(new_n775), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n739), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n704), .ZN(new_n863));
  INV_X1    g438(.A(new_n739), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n861), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n703), .ZN(new_n866));
  AOI22_X1  g441(.A1(new_n633), .A2(G142), .B1(G130), .B2(new_n476), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n467), .A2(G118), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n461), .B1(new_n868), .B2(KEYINPUT102), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT102), .B1(G106), .B2(G2105), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n869), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n627), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n807), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n863), .A2(new_n866), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n876), .B1(new_n863), .B2(new_n866), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(G162), .B(G160), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n639), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT104), .ZN(new_n883));
  AOI21_X1  g458(.A(G37), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n879), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n877), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT103), .B1(new_n886), .B2(new_n882), .ZN(new_n887));
  OAI211_X1 g462(.A(KEYINPUT103), .B(new_n882), .C1(new_n878), .C2(new_n879), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n884), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  AND2_X1   g466(.A1(new_n609), .A2(new_n607), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n892), .A2(new_n575), .A3(new_n581), .A4(new_n606), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n610), .A2(G299), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n855), .B1(G559), .B2(new_n610), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n623), .B1(new_n852), .B2(new_n854), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT105), .B1(new_n895), .B2(KEYINPUT41), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT41), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n893), .A2(new_n894), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n895), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n896), .A2(new_n907), .A3(new_n897), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n898), .B1(new_n899), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n908), .A2(new_n899), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n588), .B(KEYINPUT108), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(new_n795), .ZN(new_n912));
  XOR2_X1   g487(.A(G303), .B(G290), .Z(new_n913));
  XNOR2_X1  g488(.A(new_n912), .B(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT42), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n909), .A2(new_n910), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n909), .B2(new_n910), .ZN(new_n917));
  OAI21_X1  g492(.A(G868), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(G868), .B2(new_n850), .ZN(G295));
  OAI21_X1  g494(.A(new_n918), .B1(G868), .B2(new_n850), .ZN(G331));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n921));
  NAND2_X1  g496(.A1(G301), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n538), .A2(new_n545), .A3(KEYINPUT109), .ZN(new_n923));
  AND3_X1   g498(.A1(G168), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n922), .B1(G168), .B2(new_n923), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(new_n852), .B2(new_n854), .ZN(new_n927));
  INV_X1    g502(.A(new_n895), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n846), .B1(new_n850), .B2(new_n621), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT100), .ZN(new_n930));
  NAND3_X1  g505(.A1(G286), .A2(new_n921), .A3(G301), .ZN(new_n931));
  NAND3_X1  g506(.A1(G168), .A2(new_n922), .A3(new_n923), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n933), .A3(new_n851), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n927), .A2(new_n928), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT110), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n927), .A2(new_n934), .A3(new_n937), .A4(new_n928), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n927), .A2(new_n934), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT41), .B1(new_n893), .B2(new_n894), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n928), .B2(new_n905), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n936), .A2(new_n938), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n914), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n943), .A2(KEYINPUT111), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT111), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n939), .A2(new_n907), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n948), .A2(new_n914), .A3(new_n935), .ZN(new_n949));
  INV_X1    g524(.A(G37), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT43), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n914), .B1(new_n948), .B2(new_n935), .ZN(new_n953));
  OR3_X1    g528(.A1(new_n951), .A2(KEYINPUT43), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(KEYINPUT44), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n949), .A2(new_n956), .A3(new_n950), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(new_n945), .B2(new_n946), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT43), .B1(new_n951), .B2(new_n953), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT112), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n963));
  AOI211_X1 g538(.A(new_n963), .B(KEYINPUT44), .C1(new_n958), .C2(new_n959), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n955), .B1(new_n962), .B2(new_n964), .ZN(G397));
  INV_X1    g540(.A(G40), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n470), .A2(new_n473), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(G1384), .B1(new_n491), .B2(new_n496), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n968), .B1(new_n970), .B2(KEYINPUT50), .ZN(new_n971));
  INV_X1    g546(.A(G2084), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n969), .A2(KEYINPUT45), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n967), .B1(new_n969), .B2(KEYINPUT45), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n759), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G8), .ZN(new_n981));
  NOR2_X1   g556(.A1(G168), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT51), .B1(new_n982), .B2(KEYINPUT123), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n981), .B1(new_n975), .B2(new_n979), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n985), .B1(new_n986), .B2(new_n982), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n986), .A2(new_n982), .A3(new_n985), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n983), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n991));
  XOR2_X1   g566(.A(KEYINPUT113), .B(G1384), .Z(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(KEYINPUT45), .B(new_n993), .C1(new_n492), .C2(new_n497), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n994), .B(new_n967), .C1(KEYINPUT45), .C2(new_n969), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n991), .B1(new_n995), .B2(G2078), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n970), .A2(KEYINPUT50), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(new_n967), .A3(new_n974), .ZN(new_n998));
  INV_X1    g573(.A(G1961), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n978), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n991), .A2(G2078), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n976), .A3(new_n1002), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n1000), .A2(KEYINPUT125), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT125), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1005));
  OAI211_X1 g580(.A(G301), .B(new_n996), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(G164), .B2(new_n992), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1009), .A2(new_n967), .A3(new_n994), .A4(new_n1002), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n996), .A2(new_n1000), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1007), .B1(new_n1011), .B2(G171), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1971), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n995), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n971), .A2(new_n750), .A3(new_n974), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n981), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G303), .A2(G8), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  NAND4_X1  g597(.A1(G303), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1017), .B(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n969), .A2(new_n967), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n588), .A2(new_n788), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(G8), .A3(new_n1028), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1029), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT116), .B1(new_n1029), .B2(KEYINPUT52), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n1033));
  NOR2_X1   g608(.A1(G305), .A2(G1981), .ZN(new_n1034));
  INV_X1    g609(.A(G1981), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1033), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n981), .B1(new_n969), .B2(new_n967), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G305), .A2(G1981), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n795), .A2(new_n1035), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(KEYINPUT49), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n788), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(new_n1038), .A3(new_n1028), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1026), .B1(new_n1032), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1045), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1047), .B(KEYINPUT117), .C1(new_n1031), .C2(new_n1030), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n990), .A2(new_n1013), .A3(new_n1025), .A4(new_n1049), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n1051));
  OAI21_X1  g626(.A(new_n996), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(G171), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1011), .A2(G171), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1050), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1348), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n998), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1027), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n969), .A2(KEYINPUT121), .A3(new_n967), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G2067), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT60), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1058), .A2(new_n1064), .A3(new_n1065), .A4(new_n611), .ZN(new_n1066));
  INV_X1    g641(.A(G1996), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1001), .A2(new_n1067), .A3(new_n994), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT58), .B(G1341), .Z(new_n1069));
  NAND3_X1  g644(.A1(new_n1060), .A2(new_n1061), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n621), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1066), .B1(new_n1071), .B2(KEYINPUT59), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1058), .A2(new_n1064), .A3(new_n610), .ZN(new_n1073));
  AOI21_X1  g648(.A(G1348), .B1(new_n971), .B2(new_n974), .ZN(new_n1074));
  AOI21_X1  g649(.A(G2067), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n611), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1065), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1071), .A2(KEYINPUT59), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1072), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT56), .B(G2072), .Z(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n995), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1956), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n998), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1081), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1001), .A2(KEYINPUT120), .A3(new_n994), .A4(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1082), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT119), .B1(new_n579), .B2(new_n580), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1088), .A2(KEYINPUT57), .ZN(new_n1089));
  XNOR2_X1  g664(.A(G299), .B(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1082), .A2(new_n1084), .A3(new_n1090), .A4(new_n1086), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(KEYINPUT61), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT122), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1092), .A2(new_n1096), .A3(KEYINPUT61), .A4(new_n1093), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT61), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1079), .A2(new_n1095), .A3(new_n1097), .A4(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1093), .B(new_n611), .C1(new_n1075), .C2(new_n1074), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1102), .A2(new_n1092), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1056), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n986), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(G286), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1049), .A2(new_n1025), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT63), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT118), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1112), .A3(new_n1109), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1032), .A2(new_n1045), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1025), .A2(KEYINPUT63), .A3(new_n1114), .A4(new_n1107), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1024), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1017), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1042), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1119), .A2(G1976), .A3(G288), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1038), .B1(new_n1120), .B2(new_n1034), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1049), .A2(new_n1025), .A3(G171), .A4(new_n1052), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n1124));
  INV_X1    g699(.A(new_n982), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1106), .A2(new_n1125), .A3(new_n984), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n987), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1124), .B1(new_n1127), .B2(new_n983), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1123), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1127), .A2(new_n1124), .A3(new_n983), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1122), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1105), .A2(new_n1116), .A3(new_n1131), .ZN(new_n1132));
  OR3_X1    g707(.A1(new_n1009), .A2(KEYINPUT114), .A3(new_n968), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT114), .B1(new_n1009), .B2(new_n968), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n739), .B(new_n1067), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n775), .B(new_n1063), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n807), .B(new_n810), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(G290), .B(G1986), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1136), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1132), .A2(new_n1143), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1135), .A2(G1986), .A3(G290), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1147), .A2(KEYINPUT48), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1136), .A2(new_n1141), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(KEYINPUT48), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n810), .B(new_n808), .C1(new_n1135), .C2(new_n1139), .ZN(new_n1154));
  INV_X1    g729(.A(new_n775), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1154), .B1(G2067), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1135), .B1(new_n1156), .B2(KEYINPUT126), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(KEYINPUT126), .B2(new_n1156), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1136), .B1(new_n864), .B2(new_n1138), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1136), .A2(KEYINPUT46), .A3(new_n1067), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT46), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(new_n1135), .B2(G1996), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1159), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT47), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1153), .A2(new_n1158), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1144), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g741(.A1(G401), .A2(G229), .A3(new_n459), .A4(G227), .ZN(new_n1168));
  NAND3_X1  g742(.A1(new_n890), .A2(new_n960), .A3(new_n1168), .ZN(G225));
  INV_X1    g743(.A(G225), .ZN(G308));
endmodule


