//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996, new_n997, new_n998;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202));
  OAI21_X1  g001(.A(G127gat), .B1(new_n202), .B2(KEYINPUT1), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n204));
  INV_X1    g003(.A(G127gat), .ZN(new_n205));
  INV_X1    g004(.A(G113gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G120gat), .ZN(new_n207));
  INV_X1    g006(.A(G120gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G113gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n204), .B(new_n205), .C1(new_n207), .C2(new_n209), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n203), .A2(G134gat), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(G134gat), .B1(new_n203), .B2(new_n210), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT77), .ZN(new_n214));
  XNOR2_X1  g013(.A(G141gat), .B(G148gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n216), .B1(G155gat), .B2(G162gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n214), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G155gat), .B(G162gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G155gat), .ZN(new_n222));
  INV_X1    g021(.A(G162gat), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT2), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G141gat), .ZN(new_n225));
  INV_X1    g024(.A(G148gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G141gat), .A2(G148gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(new_n214), .A3(new_n219), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n221), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT4), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n213), .A2(KEYINPUT4), .A3(new_n231), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT4), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n241), .B1(new_n221), .B2(new_n230), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT78), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n218), .A2(new_n220), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n219), .B1(new_n229), .B2(new_n214), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n221), .A2(KEYINPUT78), .A3(new_n230), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n242), .B1(new_n248), .B2(KEYINPUT3), .ZN(new_n249));
  INV_X1    g048(.A(new_n213), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT80), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n252), .B1(new_n246), .B2(new_n247), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT80), .ZN(new_n254));
  NOR4_X1   g053(.A1(new_n253), .A2(new_n254), .A3(new_n213), .A4(new_n242), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n237), .B(new_n240), .C1(new_n251), .C2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT5), .ZN(new_n257));
  INV_X1    g056(.A(new_n248), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n232), .B1(new_n258), .B2(new_n213), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n257), .B1(new_n259), .B2(new_n239), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n239), .A2(KEYINPUT5), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n237), .B(new_n262), .C1(new_n251), .C2(new_n255), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G1gat), .B(G29gat), .Z(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G57gat), .B(G85gat), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n267), .B(new_n268), .Z(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT6), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n261), .A2(new_n269), .A3(new_n263), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n264), .A2(KEYINPUT6), .A3(new_n270), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT82), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n269), .B1(new_n261), .B2(new_n263), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(KEYINPUT82), .A3(KEYINPUT6), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n274), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  OR2_X1    g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(KEYINPUT24), .A3(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n282), .A2(KEYINPUT24), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT23), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(G169gat), .B2(G176gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT64), .B(G169gat), .ZN(new_n289));
  INV_X1    g088(.A(G176gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(KEYINPUT23), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n285), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT25), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n293), .B1(new_n295), .B2(KEYINPUT23), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n285), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT26), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT65), .B1(new_n295), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n295), .A2(new_n305), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT65), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n308), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n306), .A2(new_n286), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(new_n311), .A3(new_n282), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(new_n310), .B2(new_n282), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n304), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G226gat), .ZN(new_n316));
  INV_X1    g115(.A(G233gat), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n299), .B(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(new_n316), .B2(new_n317), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n302), .B(KEYINPUT28), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n310), .A2(new_n282), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT66), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n321), .B1(new_n312), .B2(new_n323), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n292), .A2(new_n293), .B1(new_n285), .B2(new_n297), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n320), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n318), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G211gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT73), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT73), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G211gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n331), .A3(G218gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT22), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G197gat), .B(G204gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G211gat), .B(G218gat), .Z(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n337), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n334), .A2(new_n339), .A3(new_n335), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT74), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n334), .B2(new_n335), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G8gat), .B(G36gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(G64gat), .ZN(new_n348));
  INV_X1    g147(.A(G92gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n340), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n343), .B1(new_n351), .B2(new_n342), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n338), .A2(KEYINPUT74), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n318), .A2(new_n326), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n346), .A2(new_n350), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT30), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT76), .ZN(new_n359));
  OR2_X1    g158(.A1(new_n356), .A2(new_n357), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n350), .B(KEYINPUT75), .ZN(new_n361));
  INV_X1    g160(.A(new_n346), .ZN(new_n362));
  INV_X1    g161(.A(new_n355), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n356), .A2(new_n365), .A3(new_n357), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n359), .A2(new_n360), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n280), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G78gat), .B(G106gat), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n370), .B(G22gat), .Z(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT31), .B(G50gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(KEYINPUT84), .B(new_n319), .C1(new_n341), .C2(new_n344), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n252), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT84), .B1(new_n354), .B2(new_n319), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n248), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n242), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n319), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n345), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G228gat), .A2(G233gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n378), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT85), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT85), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n378), .A2(new_n388), .A3(new_n385), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT29), .B1(new_n338), .B2(new_n340), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n230), .B(new_n221), .C1(new_n391), .C2(new_n241), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(KEYINPUT83), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n381), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n382), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n374), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n383), .B1(new_n393), .B2(new_n381), .ZN(new_n397));
  AOI211_X1 g196(.A(new_n373), .B(new_n397), .C1(new_n387), .C2(new_n389), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n372), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n378), .A2(new_n388), .A3(new_n385), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n388), .B1(new_n378), .B2(new_n385), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n395), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n373), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n390), .A2(new_n374), .A3(new_n395), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n404), .A3(new_n371), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n369), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT68), .B(G71gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(G99gat), .ZN(new_n409));
  XOR2_X1   g208(.A(G15gat), .B(G43gat), .Z(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G227gat), .A2(G233gat), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n250), .B1(new_n324), .B2(new_n325), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n299), .A2(new_n315), .A3(new_n213), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT67), .B(KEYINPUT33), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n411), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT32), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n413), .A2(new_n414), .ZN(new_n421));
  INV_X1    g220(.A(new_n412), .ZN(new_n422));
  AOI221_X4 g221(.A(new_n418), .B1(new_n416), .B2(new_n411), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT34), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n413), .A2(new_n412), .A3(new_n414), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n425), .B1(new_n426), .B2(KEYINPUT69), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(KEYINPUT69), .A3(new_n425), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OAI22_X1  g228(.A1(new_n424), .A2(KEYINPUT70), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n417), .B(new_n419), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT70), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n426), .A2(KEYINPUT69), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT34), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n431), .A2(new_n432), .A3(new_n434), .A4(new_n428), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT71), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n430), .A2(new_n435), .A3(new_n436), .A4(KEYINPUT36), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT72), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(new_n429), .B2(new_n427), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n434), .A2(KEYINPUT72), .A3(new_n428), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n424), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n431), .A2(new_n439), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT36), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT71), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n430), .A2(new_n435), .A3(KEYINPUT36), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n437), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT40), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT39), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n259), .A2(new_n239), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n237), .B1(new_n251), .B2(new_n255), .ZN(new_n452));
  AOI211_X1 g251(.A(new_n450), .B(new_n451), .C1(new_n452), .C2(new_n239), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n450), .A3(new_n239), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n269), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n449), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT86), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n458), .B(new_n449), .C1(new_n453), .C2(new_n455), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n452), .A2(new_n239), .ZN(new_n461));
  INV_X1    g260(.A(new_n451), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(KEYINPUT39), .A3(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n463), .A2(KEYINPUT40), .A3(new_n269), .A4(new_n454), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n367), .A2(new_n271), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n405), .B(new_n399), .C1(new_n460), .C2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT38), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n356), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n469));
  OAI22_X1  g268(.A1(new_n362), .A2(new_n363), .B1(new_n469), .B2(KEYINPUT37), .ZN(new_n470));
  XOR2_X1   g269(.A(KEYINPUT87), .B(KEYINPUT37), .Z(new_n471));
  NAND3_X1  g270(.A1(new_n346), .A2(new_n355), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n468), .B1(new_n473), .B2(new_n350), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n274), .A2(new_n277), .A3(new_n279), .A4(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n470), .A2(new_n467), .A3(new_n361), .A4(new_n472), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n407), .B(new_n448), .C1(new_n466), .C2(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n403), .A2(new_n404), .A3(new_n371), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n371), .B1(new_n403), .B2(new_n404), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n444), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n482), .A2(new_n280), .A3(new_n368), .A4(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT35), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND4_X1   g285(.A1(new_n405), .A2(new_n399), .A3(new_n435), .A4(new_n430), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n280), .A2(KEYINPUT35), .A3(new_n368), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n479), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G57gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(KEYINPUT93), .ZN(new_n492));
  OR2_X1    g291(.A1(KEYINPUT94), .A2(G64gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(KEYINPUT94), .A2(G64gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT93), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(G57gat), .ZN(new_n497));
  AND2_X1   g296(.A1(KEYINPUT94), .A2(G64gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(KEYINPUT94), .A2(G64gat), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G71gat), .ZN(new_n501));
  INV_X1    g300(.A(G78gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT9), .ZN(new_n503));
  NAND2_X1  g302(.A1(G71gat), .A2(G78gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n495), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n507));
  AND2_X1   g306(.A1(G57gat), .A2(G64gat), .ZN(new_n508));
  NOR2_X1   g307(.A1(G57gat), .A2(G64gat), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT92), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(KEYINPUT92), .A2(G71gat), .A3(G78gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n501), .A2(new_n502), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT95), .B1(new_n506), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT92), .B1(G71gat), .B2(G78gat), .ZN(new_n518));
  NOR2_X1   g317(.A1(G71gat), .A2(G78gat), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G57gat), .B(G64gat), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n520), .B(new_n513), .C1(new_n521), .C2(new_n507), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n495), .A2(new_n500), .A3(new_n505), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT95), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n526), .A2(KEYINPUT21), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n527), .B(new_n528), .Z(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT16), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n532), .A2(G1gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(G1gat), .B2(new_n531), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(G8gat), .ZN(new_n536));
  INV_X1    g335(.A(G8gat), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n534), .B(new_n537), .C1(G1gat), .C2(new_n531), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n539), .B1(new_n526), .B2(KEYINPUT21), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(G183gat), .ZN(new_n541));
  AND2_X1   g340(.A1(G231gat), .A2(G233gat), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n542), .ZN(new_n544));
  XNOR2_X1  g343(.A(G127gat), .B(G155gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(new_n328), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n543), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n547), .B1(new_n543), .B2(new_n544), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n530), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n550), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(new_n529), .A3(new_n548), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G99gat), .A2(G106gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT97), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(G99gat), .A3(G106gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n558), .A3(KEYINPUT8), .ZN(new_n559));
  INV_X1    g358(.A(G85gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n349), .ZN(new_n561));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT7), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT7), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(G85gat), .A3(G92gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n559), .A2(new_n561), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G99gat), .B(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n559), .A2(new_n566), .A3(new_n568), .A4(new_n561), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G29gat), .ZN(new_n573));
  INV_X1    g372(.A(G36gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(new_n574), .A3(KEYINPUT14), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT14), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n576), .B1(G29gat), .B2(G36gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(G29gat), .A2(G36gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT15), .ZN(new_n580));
  INV_X1    g379(.A(G50gat), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n580), .B1(G43gat), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G43gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(G50gat), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT90), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(new_n581), .B2(G43gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n581), .A2(G43gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n583), .A2(KEYINPUT90), .A3(G50gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT89), .B(KEYINPUT15), .Z(new_n591));
  AOI22_X1  g390(.A1(new_n590), .A2(new_n591), .B1(new_n584), .B2(new_n582), .ZN(new_n592));
  AND3_X1   g391(.A1(KEYINPUT91), .A2(G29gat), .A3(G36gat), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT91), .B1(G29gat), .B2(G36gat), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n575), .B(new_n577), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AOI221_X4 g395(.A(KEYINPUT17), .B1(new_n579), .B2(new_n585), .C1(new_n592), .C2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT17), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n590), .A2(new_n591), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n596), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n579), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n572), .B1(new_n597), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n605));
  INV_X1    g404(.A(new_n572), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n601), .A2(new_n602), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G190gat), .B(G218gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT96), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n611), .A2(KEYINPUT98), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n610), .ZN(new_n617));
  OR3_X1    g416(.A1(new_n609), .A2(KEYINPUT98), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n611), .B1(new_n618), .B2(new_n615), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n554), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n536), .A2(new_n538), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n623), .B1(new_n597), .B2(new_n603), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n539), .A2(new_n607), .ZN(new_n625));
  NAND2_X1  g424(.A1(G229gat), .A2(G233gat), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT18), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n539), .B(new_n607), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n626), .B(KEYINPUT13), .Z(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n624), .A2(KEYINPUT18), .A3(new_n625), .A4(new_n626), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n629), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G113gat), .B(G141gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G169gat), .B(G197gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n629), .A2(new_n632), .A3(new_n633), .A4(new_n640), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(new_n290), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G204gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n524), .B1(new_n522), .B2(new_n523), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n572), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n522), .A2(new_n523), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n653), .A2(new_n570), .A3(new_n571), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT10), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT10), .B1(new_n650), .B2(new_n651), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(new_n572), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n649), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n649), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n652), .A2(new_n659), .A3(new_n654), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n648), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n658), .A2(new_n660), .A3(new_n648), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n645), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n622), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n490), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n280), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT99), .B(G1gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1324gat));
  NOR2_X1   g470(.A1(new_n668), .A2(new_n368), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n532), .A2(new_n537), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n675), .A2(KEYINPUT42), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(KEYINPUT42), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n676), .B(new_n677), .C1(new_n537), .C2(new_n672), .ZN(G1325gat));
  INV_X1    g477(.A(G15gat), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n668), .A2(new_n679), .A3(new_n448), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n490), .A2(new_n483), .A3(new_n667), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(new_n679), .B2(new_n681), .ZN(G1326gat));
  NOR2_X1   g481(.A1(new_n668), .A2(new_n482), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT43), .B(G22gat), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT100), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n683), .B(new_n685), .ZN(G1327gat));
  NAND2_X1  g485(.A1(new_n490), .A2(new_n620), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n687), .A2(new_n554), .A3(new_n666), .ZN(new_n688));
  INV_X1    g487(.A(new_n280), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(new_n573), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT101), .B(KEYINPUT45), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n687), .A2(KEYINPUT44), .ZN(new_n693));
  AND4_X1   g492(.A1(KEYINPUT82), .A2(new_n264), .A3(KEYINPUT6), .A4(new_n270), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT82), .B1(new_n278), .B2(KEYINPUT6), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n367), .B1(new_n696), .B2(new_n274), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT102), .B1(new_n697), .B2(new_n482), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n464), .A2(new_n271), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n699), .A2(new_n457), .A3(new_n367), .A4(new_n459), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n482), .B(new_n700), .C1(new_n477), .C2(new_n475), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT102), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n369), .A2(new_n702), .A3(new_n406), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n698), .A2(new_n701), .A3(new_n448), .A4(new_n703), .ZN(new_n704));
  AOI22_X1  g503(.A1(new_n484), .A2(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n706), .A2(new_n707), .A3(new_n620), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n554), .A2(new_n666), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n709), .A2(new_n689), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n692), .B1(new_n573), .B2(new_n712), .ZN(G1328gat));
  NAND3_X1  g512(.A1(new_n688), .A2(new_n574), .A3(new_n367), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n714), .B(KEYINPUT46), .Z(new_n715));
  NAND3_X1  g514(.A1(new_n709), .A2(new_n367), .A3(new_n710), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT103), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n717), .B2(new_n574), .ZN(G1329gat));
  INV_X1    g517(.A(new_n448), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n709), .A2(new_n719), .A3(new_n710), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G43gat), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n688), .A2(new_n583), .A3(new_n483), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n723), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n721), .B(new_n724), .C1(new_n722), .C2(KEYINPUT47), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1330gat));
  AOI211_X1 g528(.A(KEYINPUT44), .B(new_n621), .C1(new_n704), .C2(new_n705), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n707), .B1(new_n490), .B2(new_n620), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n406), .B(new_n710), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n482), .A2(G50gat), .ZN(new_n733));
  AOI22_X1  g532(.A1(new_n732), .A2(G50gat), .B1(new_n688), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT48), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n735), .A2(KEYINPUT105), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(KEYINPUT105), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n736), .B1(new_n734), .B2(new_n737), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(G1331gat));
  NOR2_X1   g539(.A1(new_n622), .A2(new_n644), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n706), .A2(new_n664), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT106), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n689), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT107), .B(G57gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1332gat));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n742), .B(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n368), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  AND2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n749), .B2(new_n750), .ZN(G1333gat));
  OAI21_X1  g552(.A(new_n501), .B1(new_n748), .B2(new_n444), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n719), .A2(G71gat), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n754), .B(new_n755), .C1(new_n748), .C2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(G71gat), .B1(new_n743), .B2(new_n483), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n748), .A2(new_n756), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT50), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n743), .A2(new_n406), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  INV_X1    g562(.A(new_n664), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n554), .A2(new_n644), .A3(new_n764), .ZN(new_n765));
  AND4_X1   g564(.A1(G85gat), .A2(new_n709), .A3(new_n689), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n554), .A2(new_n644), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n706), .A2(new_n620), .A3(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n706), .A2(KEYINPUT51), .A3(new_n620), .A4(new_n767), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n772), .A2(new_n771), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n773), .A2(new_n774), .A3(new_n689), .A4(new_n664), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n766), .B1(new_n775), .B2(new_n560), .ZN(G1336gat));
  NOR2_X1   g575(.A1(new_n368), .A2(G92gat), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n773), .A2(new_n774), .A3(new_n664), .A4(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n367), .B(new_n765), .C1(new_n730), .C2(new_n731), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G92gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n780), .A2(new_n783), .A3(G92gat), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n780), .B2(G92gat), .ZN(new_n785));
  INV_X1    g584(.A(new_n777), .ZN(new_n786));
  AOI211_X1 g585(.A(new_n764), .B(new_n786), .C1(new_n770), .C2(new_n772), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n782), .B1(new_n788), .B2(new_n779), .ZN(G1337gat));
  NOR2_X1   g588(.A1(new_n444), .A2(G99gat), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n773), .A2(new_n774), .A3(new_n664), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n709), .A2(new_n719), .A3(new_n765), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G99gat), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(G1338gat));
  NOR3_X1   g593(.A1(new_n482), .A2(G106gat), .A3(new_n764), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n773), .A2(new_n774), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n709), .A2(new_n406), .A3(new_n765), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G106gat), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n773), .A2(new_n774), .A3(KEYINPUT111), .A4(new_n795), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n798), .A2(new_n799), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n770), .A2(new_n772), .B1(KEYINPUT110), .B2(new_n795), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n795), .A2(KEYINPUT110), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT53), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n803), .A2(new_n808), .ZN(G1339gat));
  NOR2_X1   g608(.A1(new_n630), .A2(new_n631), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n626), .B1(new_n624), .B2(new_n625), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n639), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n658), .A2(new_n660), .A3(new_n648), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n643), .B(new_n812), .C1(new_n813), .C2(new_n661), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT113), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT10), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n517), .A2(new_n525), .B1(new_n571), .B2(new_n570), .ZN(new_n818));
  INV_X1    g617(.A(new_n654), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n526), .A2(new_n606), .A3(KEYINPUT10), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n821), .A3(new_n659), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n658), .A2(new_n822), .A3(KEYINPUT54), .ZN(new_n823));
  INV_X1    g622(.A(new_n648), .ZN(new_n824));
  XOR2_X1   g623(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n658), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n816), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n659), .B1(new_n820), .B2(new_n821), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n648), .B1(new_n829), .B2(new_n825), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n658), .A2(new_n822), .A3(KEYINPUT54), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n644), .A2(new_n828), .A3(new_n663), .A4(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n620), .B1(new_n815), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n828), .A2(new_n663), .A3(new_n832), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n643), .A2(new_n812), .ZN(new_n836));
  NOR4_X1   g635(.A1(new_n835), .A2(new_n619), .A3(new_n616), .A4(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT114), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n554), .ZN(new_n839));
  INV_X1    g638(.A(new_n833), .ZN(new_n840));
  INV_X1    g639(.A(new_n836), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(KEYINPUT113), .A3(new_n664), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n814), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n621), .B1(new_n840), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n831), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT55), .B1(new_n830), .B2(new_n831), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n620), .A2(new_n663), .A3(new_n850), .A4(new_n841), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n846), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n838), .A2(new_n839), .A3(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n554), .A2(new_n621), .A3(new_n645), .A4(new_n764), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n280), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n855), .A2(new_n368), .A3(new_n482), .A4(new_n483), .ZN(new_n856));
  OAI21_X1  g655(.A(G113gat), .B1(new_n856), .B2(new_n645), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT115), .Z(new_n858));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n855), .A2(new_n859), .A3(new_n487), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n855), .B2(new_n487), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n368), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n644), .A2(new_n206), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n858), .B1(new_n863), .B2(new_n864), .ZN(G1340gat));
  INV_X1    g664(.A(new_n863), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n208), .A3(new_n664), .ZN(new_n867));
  OAI21_X1  g666(.A(G120gat), .B1(new_n856), .B2(new_n764), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1341gat));
  NOR3_X1   g668(.A1(new_n856), .A2(new_n205), .A3(new_n839), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n866), .A2(new_n554), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n205), .ZN(G1342gat));
  INV_X1    g671(.A(G134gat), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n621), .A2(new_n367), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT117), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n873), .B(new_n875), .C1(new_n860), .C2(new_n861), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n877));
  OAI21_X1  g676(.A(G134gat), .B1(new_n856), .B2(new_n621), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n877), .A2(KEYINPUT118), .A3(new_n878), .A4(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1343gat));
  NAND3_X1  g683(.A1(new_n448), .A2(new_n689), .A3(new_n368), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n835), .A2(KEYINPUT119), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n828), .A2(new_n888), .A3(new_n663), .A4(new_n832), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n644), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n620), .B1(new_n890), .B2(new_n814), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n839), .B1(new_n891), .B2(new_n837), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n482), .B1(new_n892), .B2(new_n854), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n886), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI211_X1 g694(.A(KEYINPUT57), .B(new_n482), .C1(new_n853), .C2(new_n854), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT120), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n888), .B1(new_n850), .B2(new_n663), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n889), .A2(new_n644), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n814), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n621), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n554), .B1(new_n902), .B2(new_n851), .ZN(new_n903));
  INV_X1    g702(.A(new_n854), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n406), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n885), .B1(new_n905), .B2(KEYINPUT57), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n853), .A2(new_n854), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n894), .A3(new_n406), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n898), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n644), .B1(new_n897), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(KEYINPUT121), .A3(G141gat), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n482), .B1(new_n853), .B2(new_n854), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n886), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n225), .A3(new_n644), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT120), .B1(new_n895), .B2(new_n896), .ZN(new_n917));
  INV_X1    g716(.A(new_n814), .ZN(new_n918));
  INV_X1    g717(.A(new_n900), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n887), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n851), .B1(new_n920), .B2(new_n620), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n904), .B1(new_n921), .B2(new_n839), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT57), .B1(new_n922), .B2(new_n482), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n908), .A2(new_n923), .A3(new_n898), .A4(new_n886), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n645), .B1(new_n917), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n916), .B1(new_n925), .B2(new_n225), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n911), .A2(new_n915), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT58), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT58), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n895), .A2(new_n896), .A3(new_n645), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n915), .B(new_n929), .C1(new_n930), .C2(new_n225), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n928), .A2(new_n931), .ZN(G1344gat));
  NAND3_X1  g731(.A1(new_n914), .A2(new_n226), .A3(new_n664), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n897), .A2(new_n909), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  AOI211_X1 g734(.A(KEYINPUT59), .B(new_n226), .C1(new_n935), .C2(new_n664), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT59), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n912), .A2(new_n894), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n854), .B(KEYINPUT122), .Z(new_n939));
  OAI211_X1 g738(.A(new_n894), .B(new_n406), .C1(new_n939), .C2(new_n903), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n938), .A2(new_n940), .A3(new_n664), .A4(new_n886), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n941), .A2(KEYINPUT123), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n226), .B1(new_n941), .B2(KEYINPUT123), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n937), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n933), .B1(new_n936), .B2(new_n944), .ZN(G1345gat));
  AOI21_X1  g744(.A(G155gat), .B1(new_n914), .B2(new_n554), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n554), .A2(G155gat), .ZN(new_n947));
  XOR2_X1   g746(.A(new_n947), .B(KEYINPUT124), .Z(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n935), .B2(new_n948), .ZN(G1346gat));
  OAI21_X1  g748(.A(G162gat), .B1(new_n934), .B2(new_n621), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n719), .A2(new_n280), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n912), .A2(new_n223), .A3(new_n875), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1347gat));
  NOR2_X1   g752(.A1(new_n689), .A2(new_n368), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n483), .ZN(new_n955));
  XOR2_X1   g754(.A(new_n955), .B(KEYINPUT125), .Z(new_n956));
  NAND3_X1  g755(.A1(new_n956), .A2(new_n482), .A3(new_n907), .ZN(new_n957));
  OAI21_X1  g756(.A(G169gat), .B1(new_n957), .B2(new_n645), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n689), .B1(new_n853), .B2(new_n854), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(new_n367), .A3(new_n487), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(new_n289), .A3(new_n644), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n958), .A2(new_n962), .ZN(G1348gat));
  AOI21_X1  g762(.A(G176gat), .B1(new_n961), .B2(new_n664), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n957), .A2(new_n764), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(G176gat), .ZN(G1349gat));
  OAI21_X1  g765(.A(G183gat), .B1(new_n957), .B2(new_n839), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n961), .A2(new_n300), .A3(new_n554), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g769(.A(G190gat), .B1(new_n957), .B2(new_n621), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT61), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n961), .A2(new_n301), .A3(new_n620), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1351gat));
  NAND2_X1  g773(.A1(new_n954), .A2(new_n448), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n938), .A2(new_n940), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n978), .B1(new_n977), .B2(new_n976), .ZN(new_n979));
  OAI21_X1  g778(.A(G197gat), .B1(new_n979), .B2(new_n645), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n959), .A2(new_n367), .A3(new_n406), .A4(new_n448), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n981), .A2(G197gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n980), .B1(new_n645), .B2(new_n982), .ZN(G1352gat));
  OAI21_X1  g782(.A(G204gat), .B1(new_n979), .B2(new_n764), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n981), .A2(G204gat), .A3(new_n764), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT62), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n984), .A2(new_n986), .ZN(G1353gat));
  OR3_X1    g786(.A1(new_n976), .A2(new_n839), .A3(new_n975), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n988), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n989));
  INV_X1    g788(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g789(.A(KEYINPUT63), .B1(new_n988), .B2(G211gat), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n329), .A2(new_n331), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n554), .A2(new_n992), .ZN(new_n993));
  OAI22_X1  g792(.A1(new_n990), .A2(new_n991), .B1(new_n981), .B2(new_n993), .ZN(G1354gat));
  INV_X1    g793(.A(G218gat), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n979), .A2(new_n995), .A3(new_n621), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n995), .B1(new_n981), .B2(new_n621), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT127), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n996), .A2(new_n998), .ZN(G1355gat));
endmodule


