//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G104), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  AOI21_X1  g006(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(G107), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n191), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G101), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n197), .B(new_n191), .C1(new_n193), .C2(new_n194), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT72), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT4), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n196), .A2(new_n198), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT0), .A4(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n205), .A2(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n203), .A2(G143), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT0), .B(G128), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n195), .B(G101), .C1(new_n199), .C2(new_n200), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n202), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT1), .B1(new_n205), .B2(G146), .ZN(new_n216));
  OAI211_X1 g030(.A(G128), .B(new_n216), .C1(new_n208), .C2(new_n209), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n204), .B(new_n206), .C1(KEYINPUT1), .C2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n190), .A2(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n192), .A2(G107), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n197), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n189), .B1(new_n190), .B2(G104), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n192), .A2(KEYINPUT3), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n224), .A2(new_n221), .B1(new_n225), .B2(new_n190), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n223), .B1(new_n226), .B2(new_n197), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n220), .A2(new_n227), .A3(KEYINPUT10), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n215), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT10), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT73), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(new_n220), .B2(new_n227), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n190), .A2(G104), .ZN(new_n233));
  OAI21_X1  g047(.A(G101), .B1(new_n194), .B2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n198), .A2(new_n217), .A3(new_n219), .A4(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(KEYINPUT73), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n230), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT11), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(G137), .ZN(new_n240));
  INV_X1    g054(.A(G137), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(KEYINPUT11), .A3(G134), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(G137), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G131), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n240), .A2(new_n242), .A3(new_n246), .A4(new_n243), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(KEYINPUT74), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT74), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(new_n245), .B2(new_n247), .ZN(new_n251));
  OR2_X1    g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n229), .A2(new_n237), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(G110), .B(G140), .ZN(new_n254));
  INV_X1    g068(.A(G227), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G953), .ZN(new_n256));
  XOR2_X1   g070(.A(new_n254), .B(new_n256), .Z(new_n257));
  NAND2_X1  g071(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT12), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT76), .B1(new_n220), .B2(new_n227), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n198), .A2(new_n234), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n217), .A2(new_n219), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT76), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n260), .B(new_n264), .C1(new_n232), .C2(new_n236), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n248), .A2(KEYINPUT75), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n259), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n263), .B1(new_n261), .B2(new_n262), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n220), .A2(new_n227), .A3(new_n231), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n235), .A2(KEYINPUT73), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI211_X1 g088(.A(KEYINPUT12), .B(new_n266), .C1(new_n271), .C2(new_n274), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n258), .A2(new_n268), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT10), .B1(new_n272), .B2(new_n273), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n215), .A2(new_n228), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n248), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n257), .B1(new_n253), .B2(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n187), .B(new_n188), .C1(new_n276), .C2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n249), .A2(new_n251), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n277), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n257), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n279), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n275), .A2(new_n268), .A3(new_n283), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n286), .B(G469), .C1(new_n287), .C2(new_n257), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n187), .A2(new_n188), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n281), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G221), .ZN(new_n292));
  XOR2_X1   g106(.A(KEYINPUT9), .B(G234), .Z(new_n293));
  AOI21_X1  g107(.A(new_n292), .B1(new_n293), .B2(new_n188), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT16), .ZN(new_n299));
  INV_X1    g113(.A(G140), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n300), .A3(G125), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(G125), .ZN(new_n302));
  INV_X1    g116(.A(G125), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n301), .B1(new_n305), .B2(new_n299), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n203), .ZN(new_n307));
  OAI211_X1 g121(.A(G146), .B(new_n301), .C1(new_n305), .C2(new_n299), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n218), .A2(G119), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n218), .A2(G119), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT67), .ZN(new_n314));
  INV_X1    g128(.A(G119), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(G128), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n314), .B1(new_n316), .B2(KEYINPUT23), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n312), .A2(KEYINPUT67), .A3(new_n311), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n313), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G110), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n316), .A2(new_n310), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT24), .B(G110), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n309), .B(new_n320), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G110), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n313), .B(new_n324), .C1(new_n317), .C2(new_n318), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT68), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n321), .A2(new_n322), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G125), .B(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n203), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n308), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n326), .B1(new_n325), .B2(new_n327), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n323), .B(KEYINPUT69), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT22), .B(G137), .ZN(new_n334));
  INV_X1    g148(.A(G953), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(G221), .A3(G234), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n334), .B(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n323), .B1(new_n331), .B2(new_n332), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT69), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n333), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n339), .B1(new_n343), .B2(new_n337), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT71), .ZN(new_n345));
  INV_X1    g159(.A(G217), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(G234), .B2(new_n188), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(G902), .ZN(new_n348));
  XOR2_X1   g162(.A(new_n348), .B(KEYINPUT70), .Z(new_n349));
  AND3_X1   g163(.A1(new_n344), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n345), .B1(new_n344), .B2(new_n349), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT25), .B1(new_n344), .B2(new_n188), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n338), .B1(new_n342), .B2(new_n333), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n355));
  NOR4_X1   g169(.A1(new_n354), .A2(new_n339), .A3(new_n355), .A4(G902), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n347), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  OR2_X1    g172(.A1(KEYINPUT2), .A2(G113), .ZN(new_n359));
  NAND2_X1  g173(.A1(KEYINPUT2), .A2(G113), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G116), .B(G119), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n359), .A3(new_n360), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(KEYINPUT66), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT66), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n366), .B1(new_n361), .B2(new_n362), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n363), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n213), .A2(new_n248), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n239), .A2(G137), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n241), .A2(G134), .ZN(new_n371));
  OAI21_X1  g185(.A(G131), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n217), .A2(new_n247), .A3(new_n372), .A4(new_n219), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n369), .A2(KEYINPUT30), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n212), .B(KEYINPUT64), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT65), .ZN(new_n376));
  OR2_X1    g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(new_n376), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n375), .A2(new_n248), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n368), .B(new_n374), .C1(new_n379), .C2(KEYINPUT30), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n369), .A2(new_n373), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(new_n368), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(G237), .A2(G953), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G210), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(new_n197), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n386), .B(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n380), .A2(new_n383), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT31), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n382), .A2(KEYINPUT28), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n375), .A2(new_n248), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n377), .A2(new_n378), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n368), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n382), .A2(KEYINPUT28), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n392), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n388), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT31), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n380), .A2(new_n400), .A3(new_n383), .A4(new_n389), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n391), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(G472), .A2(G902), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(KEYINPUT32), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT32), .B1(new_n402), .B2(new_n403), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n374), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n408), .B1(new_n395), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n382), .B1(new_n410), .B2(new_n368), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(new_n389), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT29), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n398), .B2(new_n388), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n381), .A2(new_n368), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n392), .A2(new_n397), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n389), .A2(KEYINPUT29), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n188), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G472), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n358), .B1(new_n407), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n384), .A2(G214), .ZN(new_n423));
  NOR2_X1   g237(.A1(KEYINPUT82), .A2(G143), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n384), .B(G214), .C1(KEYINPUT82), .C2(G143), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n422), .B1(new_n427), .B2(G131), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT17), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(G131), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT83), .A4(new_n246), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n428), .A2(new_n429), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n307), .A2(new_n308), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n427), .A2(KEYINPUT17), .A3(G131), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(G113), .B(G122), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(G104), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n305), .A2(G146), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n330), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT18), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(new_n246), .ZN(new_n442));
  OAI221_X1 g256(.A(new_n440), .B1(new_n427), .B2(new_n442), .C1(new_n430), .C2(new_n441), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n435), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n438), .B1(new_n435), .B2(new_n443), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n188), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g262(.A(KEYINPUT87), .B(new_n188), .C1(new_n444), .C2(new_n445), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(G475), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(G475), .A2(G902), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n451), .B(KEYINPUT86), .Z(new_n452));
  INV_X1    g266(.A(KEYINPUT19), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n305), .B2(KEYINPUT84), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT84), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n329), .A2(new_n455), .A3(KEYINPUT19), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n203), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT85), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT85), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(new_n461), .A3(new_n203), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n459), .A2(new_n460), .A3(new_n308), .A4(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n438), .B1(new_n463), .B2(new_n443), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n452), .B1(new_n444), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT20), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n467), .B(new_n452), .C1(new_n444), .C2(new_n464), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(G116), .B(G122), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(new_n190), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n218), .A2(G143), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT13), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n239), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n205), .A2(G128), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n472), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n476), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n471), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G116), .ZN(new_n480));
  OAI211_X1 g294(.A(KEYINPUT14), .B(G107), .C1(new_n480), .C2(G122), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n471), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n476), .B(G134), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n470), .A2(KEYINPUT14), .A3(G107), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n479), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n293), .A2(G217), .A3(new_n335), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n486), .A2(new_n488), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n188), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G478), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n492), .A2(KEYINPUT15), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n491), .B(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n335), .A2(G952), .ZN(new_n495));
  INV_X1    g309(.A(G234), .ZN(new_n496));
  INV_X1    g310(.A(G237), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(G902), .B(G953), .C1(new_n496), .C2(new_n497), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT88), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT21), .B(G898), .Z(new_n501));
  OAI21_X1  g315(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n450), .A2(new_n469), .A3(new_n494), .A4(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(G210), .B1(G237), .B2(G902), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n368), .A2(new_n214), .A3(new_n202), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n364), .A2(KEYINPUT66), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n361), .A2(new_n366), .A3(new_n362), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(G113), .ZN(new_n511));
  XOR2_X1   g325(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n512));
  AND2_X1   g326(.A1(new_n315), .A2(G116), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n362), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n510), .A2(new_n227), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n507), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g333(.A(G110), .B(G122), .Z(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n520), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n507), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(KEYINPUT6), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n262), .A2(new_n303), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n212), .A2(G125), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G224), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(G953), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n529), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n525), .A2(new_n526), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT6), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n519), .A2(new_n534), .A3(new_n520), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n524), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT80), .B(KEYINPUT8), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n520), .B(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n362), .A2(KEYINPUT5), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n514), .A2(new_n539), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n510), .A2(new_n227), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n227), .B1(new_n510), .B2(new_n517), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n538), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT81), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(KEYINPUT81), .B(new_n538), .C1(new_n541), .C2(new_n542), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT7), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n532), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n525), .A2(new_n526), .B1(KEYINPUT7), .B2(new_n531), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n545), .A2(new_n523), .A3(new_n546), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n188), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n506), .B1(new_n536), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n524), .A2(new_n533), .A3(new_n535), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n554), .A2(new_n188), .A3(new_n505), .A4(new_n551), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G214), .B1(G237), .B2(G902), .ZN(new_n557));
  XOR2_X1   g371(.A(new_n557), .B(KEYINPUT78), .Z(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n298), .A2(new_n421), .A3(new_n504), .A4(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(G101), .ZN(G3));
  OAI21_X1  g376(.A(new_n557), .B1(new_n555), .B2(KEYINPUT89), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n556), .B2(KEYINPUT89), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n298), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n358), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n402), .A2(new_n188), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G472), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n402), .A2(new_n403), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n450), .A2(new_n469), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n491), .A2(new_n492), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT33), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n489), .A2(new_n575), .A3(new_n490), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT91), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n486), .B2(KEYINPUT90), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT90), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n487), .B2(KEYINPUT91), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n578), .A2(new_n487), .B1(new_n486), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n576), .B1(new_n581), .B2(new_n575), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n492), .A2(G902), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n574), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n573), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n586), .A2(new_n502), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n566), .A2(new_n567), .A3(new_n572), .A4(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(KEYINPUT34), .B(G104), .Z(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(G6));
  NAND3_X1  g404(.A1(new_n352), .A2(new_n357), .A3(new_n502), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n469), .A2(KEYINPUT92), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT92), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n466), .A2(new_n593), .A3(new_n468), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n494), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n450), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n566), .A2(new_n572), .A3(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT35), .B(G107), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G9));
  NAND3_X1  g415(.A1(new_n298), .A2(new_n504), .A3(new_n560), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n338), .A2(KEYINPUT36), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT93), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n604), .B(new_n340), .Z(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n349), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n357), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n572), .A2(KEYINPUT94), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT94), .ZN(new_n609));
  INV_X1    g423(.A(new_n607), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(new_n571), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n602), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT37), .B(G110), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G12));
  NOR2_X1   g429(.A1(new_n500), .A2(G900), .ZN(new_n616));
  INV_X1    g430(.A(new_n498), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n618), .B(KEYINPUT95), .Z(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n595), .A2(new_n450), .A3(new_n596), .A4(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n407), .B2(new_n420), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n298), .A2(new_n622), .A3(new_n564), .A4(new_n607), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G128), .ZN(G30));
  XOR2_X1   g438(.A(new_n619), .B(KEYINPUT39), .Z(new_n625));
  AND2_X1   g439(.A1(new_n298), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT97), .B(KEYINPUT40), .Z(new_n627));
  OR2_X1    g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n389), .B1(new_n383), .B2(new_n416), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n630), .B(KEYINPUT96), .Z(new_n631));
  INV_X1    g445(.A(new_n390), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n188), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G472), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n407), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n450), .A2(new_n469), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n607), .A2(new_n636), .A3(new_n494), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n557), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n556), .B(KEYINPUT38), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n628), .A2(new_n629), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(new_n205), .ZN(G45));
  INV_X1    g459(.A(KEYINPUT32), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n570), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n420), .A3(new_n404), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n573), .A2(new_n585), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n619), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n651), .A2(new_n298), .A3(new_n564), .A4(new_n607), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G146), .ZN(G48));
  INV_X1    g467(.A(new_n563), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n553), .A2(KEYINPUT89), .A3(new_n555), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n280), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n265), .A2(new_n267), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT12), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n265), .A2(new_n259), .A3(new_n267), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n659), .A2(new_n257), .A3(new_n253), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n188), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G469), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n295), .A3(new_n281), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n656), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n666), .A2(new_n587), .A3(new_n648), .A4(new_n567), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT41), .B(G113), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G15));
  NAND3_X1  g483(.A1(new_n598), .A2(new_n666), .A3(new_n648), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G116), .ZN(G18));
  AOI21_X1  g485(.A(new_n503), .B1(new_n357), .B2(new_n606), .ZN(new_n672));
  INV_X1    g486(.A(new_n665), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n648), .A2(new_n564), .A3(new_n672), .A4(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT99), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n666), .A2(KEYINPUT99), .A3(new_n648), .A4(new_n672), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G119), .ZN(G21));
  NAND2_X1  g493(.A1(new_n417), .A2(new_n388), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n391), .A2(new_n401), .A3(new_n680), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n568), .A2(G472), .B1(new_n403), .B2(new_n681), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n682), .A2(new_n357), .A3(new_n352), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n573), .A2(new_n502), .A3(new_n596), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n656), .A2(new_n665), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G122), .ZN(G24));
  NAND3_X1  g501(.A1(new_n650), .A2(new_n682), .A3(new_n607), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n688), .A2(new_n656), .A3(new_n665), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT100), .B(G125), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G27));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n296), .A2(KEYINPUT101), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n291), .A2(new_n694), .A3(new_n295), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n553), .A2(new_n555), .A3(new_n557), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  AND4_X1   g511(.A1(KEYINPUT102), .A2(new_n693), .A3(new_n695), .A4(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n696), .B1(new_n296), .B2(KEYINPUT101), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT102), .B1(new_n699), .B2(new_n695), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n421), .B(new_n650), .C1(new_n698), .C2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n692), .B1(new_n701), .B2(KEYINPUT104), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT104), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  AOI211_X1 g519(.A(KEYINPUT104), .B(new_n692), .C1(new_n701), .C2(new_n703), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT105), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n704), .A2(KEYINPUT42), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n708), .B(new_n709), .C1(new_n702), .C2(new_n704), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G131), .ZN(G33));
  INV_X1    g526(.A(new_n621), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n421), .B(new_n713), .C1(new_n698), .C2(new_n700), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G134), .ZN(G36));
  NAND2_X1  g529(.A1(new_n636), .A2(new_n585), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n716), .B1(KEYINPUT106), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n718), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n571), .A3(new_n607), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT107), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n287), .A2(new_n257), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n279), .B2(new_n285), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n726), .A2(KEYINPUT45), .ZN(new_n727));
  OAI21_X1  g541(.A(G469), .B1(new_n726), .B2(KEYINPUT45), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n289), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT46), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n281), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n730), .A2(KEYINPUT46), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n295), .B(new_n625), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n696), .B1(new_n721), .B2(new_n722), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n724), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G137), .ZN(G39));
  OAI21_X1  g552(.A(new_n295), .B1(new_n732), .B2(new_n733), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n739), .A2(KEYINPUT47), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(KEYINPUT47), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n650), .A2(new_n358), .A3(new_n697), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n648), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n740), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G140), .ZN(G42));
  AND3_X1   g559(.A1(new_n720), .A2(new_n617), .A3(new_n683), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n666), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n635), .A2(new_n358), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n665), .A2(new_n498), .A3(new_n696), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n747), .B(new_n495), .C1(new_n649), .C2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n720), .A2(new_n749), .ZN(new_n752));
  INV_X1    g566(.A(new_n421), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT48), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n640), .A2(new_n639), .A3(new_n673), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT112), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n757), .A2(new_n746), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n759), .B1(new_n757), .B2(new_n746), .ZN(new_n760));
  AOI22_X1  g574(.A1(KEYINPUT50), .A2(new_n758), .B1(new_n760), .B2(KEYINPUT114), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(KEYINPUT114), .B2(new_n760), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n750), .A2(new_n573), .A3(new_n585), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n682), .A2(new_n607), .ZN(new_n764));
  INV_X1    g578(.A(new_n752), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n664), .A2(new_n281), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n295), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n740), .B2(new_n741), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n746), .A2(new_n697), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n762), .B(new_n766), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n772));
  AOI211_X1 g586(.A(new_n751), .B(new_n755), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(new_n772), .B2(new_n771), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n450), .A2(new_n469), .A3(new_n494), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n502), .B(new_n775), .C1(new_n636), .C2(new_n585), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n776), .A2(new_n571), .A3(new_n358), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n298), .A3(new_n560), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n561), .B(new_n778), .C1(new_n602), .C2(new_n612), .ZN(new_n779));
  INV_X1    g593(.A(new_n688), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n698), .B2(new_n700), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n595), .A2(new_n450), .A3(new_n494), .A4(new_n620), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n610), .A2(new_n782), .A3(new_n696), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n298), .A3(new_n648), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n676), .A2(new_n677), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n686), .A2(new_n667), .A3(new_n670), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT108), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n587), .A2(new_n567), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n648), .A2(new_n564), .A3(new_n673), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n789), .A2(new_n790), .B1(new_n683), .B2(new_n685), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT108), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n678), .A3(new_n792), .A4(new_n670), .ZN(new_n793));
  AOI211_X1 g607(.A(new_n779), .B(new_n785), .C1(new_n788), .C2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n707), .A2(new_n710), .A3(new_n714), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n780), .A2(new_n666), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n656), .A2(new_n296), .A3(new_n619), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n635), .A3(new_n637), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n652), .A2(new_n623), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT52), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n296), .A2(new_n297), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT77), .B1(new_n291), .B2(new_n295), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n564), .B(new_n607), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n689), .B1(new_n804), .B2(new_n622), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n806), .A3(new_n652), .A4(new_n798), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n800), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT53), .B1(new_n795), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n795), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT110), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n799), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT111), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n799), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n814), .A2(new_n800), .A3(new_n807), .A4(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n799), .A2(new_n812), .A3(new_n815), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n815), .B1(new_n799), .B2(new_n812), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n808), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT53), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n821), .B1(new_n795), .B2(new_n810), .ZN(new_n822));
  OAI211_X1 g636(.A(KEYINPUT54), .B(new_n809), .C1(new_n811), .C2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n795), .B2(new_n808), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n817), .A2(new_n820), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n791), .A2(new_n678), .A3(new_n670), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n714), .A2(KEYINPUT53), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n828), .A2(new_n829), .A3(new_n779), .A4(new_n785), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n827), .B(new_n830), .C1(new_n705), .C2(new_n706), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n825), .A2(new_n826), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n823), .A2(new_n832), .ZN(new_n833));
  OAI22_X1  g647(.A1(new_n774), .A2(new_n833), .B1(G952), .B2(G953), .ZN(new_n834));
  XOR2_X1   g648(.A(new_n767), .B(KEYINPUT49), .Z(new_n835));
  NOR3_X1   g649(.A1(new_n716), .A2(new_n294), .A3(new_n559), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n748), .A2(new_n835), .A3(new_n640), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n834), .A2(new_n837), .ZN(G75));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n825), .A2(new_n831), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(G210), .A3(G902), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT56), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n524), .A2(new_n535), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT115), .ZN(new_n844));
  XOR2_X1   g658(.A(new_n533), .B(KEYINPUT55), .Z(new_n845));
  XNOR2_X1  g659(.A(new_n844), .B(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n841), .A2(new_n842), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n335), .A2(G952), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n847), .B1(new_n841), .B2(new_n842), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n839), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n841), .A2(new_n842), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n846), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(KEYINPUT116), .A3(new_n850), .A4(new_n848), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n853), .A2(new_n856), .ZN(G51));
  XNOR2_X1  g671(.A(new_n289), .B(KEYINPUT57), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n825), .A2(new_n826), .A3(new_n831), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n826), .B1(new_n825), .B2(new_n831), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(KEYINPUT117), .B(new_n858), .C1(new_n859), .C2(new_n860), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n662), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n188), .B1(new_n825), .B2(new_n831), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n729), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n849), .B1(new_n865), .B2(new_n867), .ZN(G54));
  NAND3_X1  g682(.A1(new_n866), .A2(KEYINPUT58), .A3(G475), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n444), .A2(new_n464), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n850), .B1(new_n869), .B2(new_n871), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n870), .B1(new_n869), .B2(new_n871), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G60));
  NAND2_X1  g689(.A1(G478), .A2(G902), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT121), .ZN(new_n877));
  XOR2_X1   g691(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n878));
  XOR2_X1   g692(.A(new_n877), .B(new_n878), .Z(new_n879));
  NAND2_X1  g693(.A1(new_n833), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n582), .B(KEYINPUT119), .Z(new_n882));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n879), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n823), .B2(new_n832), .ZN(new_n885));
  INV_X1    g699(.A(new_n882), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT122), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n859), .A2(new_n860), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n882), .A2(new_n884), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n849), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n883), .A2(new_n887), .A3(new_n890), .ZN(G63));
  NAND2_X1  g705(.A1(G217), .A2(G902), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT60), .Z(new_n893));
  NAND3_X1  g707(.A1(new_n840), .A2(new_n605), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n850), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n344), .B1(new_n840), .B2(new_n893), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n896), .A2(KEYINPUT123), .A3(new_n897), .A4(new_n899), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n897), .A2(KEYINPUT123), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n897), .A2(KEYINPUT123), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n901), .B(new_n902), .C1(new_n895), .C2(new_n898), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n900), .A2(new_n903), .ZN(G66));
  AOI21_X1  g718(.A(new_n335), .B1(new_n501), .B2(G224), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n788), .A2(new_n793), .ZN(new_n906));
  INV_X1    g720(.A(new_n779), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n905), .B1(new_n908), .B2(new_n335), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n844), .B1(G898), .B2(new_n335), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n909), .B(new_n910), .Z(G69));
  NAND3_X1  g725(.A1(new_n564), .A2(new_n573), .A3(new_n596), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n734), .A2(new_n753), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT126), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n805), .A2(new_n652), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT125), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n744), .A2(new_n737), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n914), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(new_n711), .A3(new_n714), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n335), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n457), .B(KEYINPUT124), .Z(new_n921));
  XOR2_X1   g735(.A(new_n410), .B(new_n921), .Z(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n255), .B2(G953), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(G900), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n922), .B2(new_n255), .ZN(new_n926));
  MUX2_X1   g740(.A(new_n596), .B(new_n585), .S(new_n573), .Z(new_n927));
  NAND4_X1  g741(.A1(new_n626), .A2(new_n421), .A3(new_n697), .A4(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n744), .A2(new_n737), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n930));
  OR3_X1    g744(.A1(new_n644), .A2(new_n930), .A3(new_n916), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n930), .B1(new_n644), .B2(new_n916), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n922), .A2(new_n335), .ZN(new_n934));
  OAI221_X1 g748(.A(new_n924), .B1(new_n335), .B2(new_n926), .C1(new_n933), .C2(new_n934), .ZN(G72));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n907), .A3(new_n906), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n937));
  NAND2_X1  g751(.A1(G472), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT63), .Z(new_n939));
  NAND3_X1  g753(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  AOI211_X1 g754(.A(new_n908), .B(new_n929), .C1(new_n931), .C2(new_n932), .ZN(new_n941));
  INV_X1    g755(.A(new_n939), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT127), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n411), .A2(new_n388), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n940), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n412), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n942), .B1(new_n946), .B2(new_n390), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n809), .B(new_n947), .C1(new_n811), .C2(new_n822), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n939), .B1(new_n919), .B2(new_n908), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n411), .A2(new_n388), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n849), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n945), .A2(new_n948), .A3(new_n951), .ZN(G57));
endmodule


