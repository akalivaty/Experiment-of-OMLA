//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT78), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT11), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G137), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT11), .A3(G134), .ZN(new_n195));
  AND2_X1   g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT66), .B1(new_n194), .B2(G134), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n192), .A3(G137), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n196), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n193), .A2(new_n197), .A3(new_n199), .A4(new_n195), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G131), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT64), .A2(G146), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT64), .A2(G146), .ZN(new_n207));
  OAI21_X1  g021(.A(G143), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n208), .A2(new_n209), .A3(G128), .A4(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n214), .B1(new_n208), .B2(KEYINPUT1), .ZN(new_n215));
  INV_X1    g029(.A(G143), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n206), .A2(new_n207), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(new_n216), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n213), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G104), .ZN(new_n221));
  OAI21_X1  g035(.A(G107), .B1(new_n221), .B2(KEYINPUT3), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT79), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(G107), .ZN(new_n227));
  INV_X1    g041(.A(G107), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(KEYINPUT79), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n225), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G101), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n224), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(G104), .A2(G107), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT79), .B(G107), .ZN(new_n234));
  OAI211_X1 g048(.A(G101), .B(new_n233), .C1(new_n234), .C2(G104), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n220), .A2(KEYINPUT10), .A3(new_n232), .A4(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G104), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n228), .A2(KEYINPUT79), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n226), .A2(G107), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n222), .A2(new_n223), .ZN(new_n242));
  OAI21_X1  g056(.A(G101), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n232), .A2(new_n243), .A3(KEYINPUT4), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n245), .B(G101), .C1(new_n241), .C2(new_n242), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT0), .B(G128), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n219), .B2(new_n249), .ZN(new_n250));
  OR2_X1    g064(.A1(KEYINPUT64), .A2(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT64), .A2(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n211), .B1(new_n253), .B2(G143), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT0), .A3(G128), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n251), .A2(new_n216), .A3(new_n252), .ZN(new_n256));
  INV_X1    g070(.A(new_n217), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n249), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(KEYINPUT65), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n250), .A2(new_n255), .A3(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n236), .B1(new_n247), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n232), .A2(new_n235), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n214), .B1(new_n257), .B2(KEYINPUT1), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n213), .B1(new_n254), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT10), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n205), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  AOI211_X1 g082(.A(new_n248), .B(new_n249), .C1(new_n256), .C2(new_n257), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT65), .B1(new_n258), .B2(new_n259), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n271), .A2(new_n255), .A3(new_n246), .A4(new_n244), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n266), .A2(new_n232), .A3(new_n235), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT10), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n205), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n272), .A2(new_n275), .A3(new_n276), .A4(new_n236), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n268), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(G110), .B(G140), .ZN(new_n279));
  INV_X1    g093(.A(G953), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n280), .A2(G227), .ZN(new_n281));
  XOR2_X1   g095(.A(new_n279), .B(new_n281), .Z(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT81), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n278), .A2(KEYINPUT81), .A3(new_n283), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n209), .B1(new_n253), .B2(G143), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n258), .B1(new_n288), .B2(new_n214), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n263), .A2(new_n289), .A3(new_n213), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n273), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n205), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT12), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n276), .B1(new_n290), .B2(new_n273), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT12), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(new_n277), .A3(new_n282), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n286), .A2(new_n287), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G469), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT70), .B(G902), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n277), .A2(new_n282), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT80), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT80), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n277), .A2(new_n306), .A3(new_n282), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n268), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n295), .B(new_n293), .ZN(new_n309));
  INV_X1    g123(.A(new_n277), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n283), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G902), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n300), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n190), .B1(new_n303), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G214), .B1(G237), .B2(G902), .ZN(new_n316));
  OAI21_X1  g130(.A(G210), .B1(G237), .B2(G902), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT83), .B(G224), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n280), .ZN(new_n319));
  XOR2_X1   g133(.A(new_n319), .B(KEYINPUT82), .Z(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(new_n271), .B2(new_n255), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n289), .A2(new_n322), .A3(new_n213), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n321), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n261), .A2(G125), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(new_n324), .A3(new_n320), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(G116), .B(G119), .Z(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT2), .B(G113), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n330), .B(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n244), .A2(new_n332), .A3(new_n246), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT5), .ZN(new_n334));
  INV_X1    g148(.A(G119), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(G116), .ZN(new_n336));
  OAI211_X1 g150(.A(G113), .B(new_n336), .C1(new_n330), .C2(new_n334), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n330), .A2(new_n331), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n232), .A2(new_n337), .A3(new_n338), .A4(new_n235), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  XOR2_X1   g154(.A(G110), .B(G122), .Z(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n341), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n333), .A2(new_n343), .A3(new_n339), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(KEYINPUT6), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT6), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n340), .A2(new_n346), .A3(new_n341), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n329), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT84), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n329), .A2(new_n345), .A3(KEYINPUT84), .A4(new_n347), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n319), .A2(KEYINPUT7), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(new_n323), .B2(new_n325), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n337), .A2(new_n338), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n263), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n339), .ZN(new_n357));
  XOR2_X1   g171(.A(new_n341), .B(KEYINPUT8), .Z(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n327), .A2(KEYINPUT7), .A3(new_n319), .A4(new_n324), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n354), .A2(new_n359), .A3(new_n360), .A4(new_n344), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n313), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n317), .B1(new_n352), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n317), .ZN(new_n365));
  AOI211_X1 g179(.A(new_n365), .B(new_n362), .C1(new_n350), .C2(new_n351), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n316), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n315), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n205), .A2(new_n255), .A3(new_n250), .A4(new_n260), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT30), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n194), .A2(G134), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n192), .A2(G137), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G131), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n220), .A2(new_n202), .A3(new_n374), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n369), .A2(new_n370), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n370), .B1(new_n369), .B2(new_n375), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n332), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(G101), .ZN(new_n380));
  INV_X1    g194(.A(G237), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n280), .A3(G210), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n380), .B(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n332), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n369), .A2(new_n384), .A3(new_n375), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n378), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT31), .ZN(new_n387));
  XOR2_X1   g201(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n388));
  AND3_X1   g202(.A1(new_n369), .A2(new_n384), .A3(new_n375), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n384), .B1(new_n369), .B2(new_n375), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT28), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n385), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n383), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT31), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n378), .A2(new_n397), .A3(new_n383), .A4(new_n385), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n387), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(G472), .A2(G902), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT32), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT32), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n399), .A2(new_n403), .A3(new_n400), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n369), .A2(new_n375), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT30), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n369), .A2(new_n370), .A3(new_n375), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n384), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n395), .B1(new_n409), .B2(new_n389), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT29), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n391), .A2(new_n383), .A3(new_n393), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT68), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n378), .A2(new_n385), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT29), .B1(new_n416), .B2(new_n395), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT68), .A3(new_n412), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT28), .B1(new_n389), .B2(new_n390), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT69), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n406), .A2(new_n332), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n385), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT69), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT28), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n421), .A2(new_n425), .A3(KEYINPUT29), .A4(new_n393), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n302), .B1(new_n426), .B2(new_n395), .ZN(new_n427));
  OAI21_X1  g241(.A(G472), .B1(new_n419), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n405), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G140), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G125), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(KEYINPUT16), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n430), .A2(KEYINPUT72), .A3(G125), .ZN(new_n434));
  XNOR2_X1  g248(.A(G125), .B(G140), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT72), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT16), .ZN(new_n438));
  OAI211_X1 g252(.A(G146), .B(new_n433), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT73), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT24), .B(G110), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n335), .A2(G128), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n214), .A2(G119), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT71), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n444), .B1(new_n442), .B2(new_n443), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n441), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G110), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n443), .A2(KEYINPUT23), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n443), .A2(KEYINPUT23), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n448), .B(new_n442), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n447), .A2(new_n451), .B1(new_n253), .B2(new_n435), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n322), .A2(G140), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n431), .A2(new_n453), .A3(new_n436), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n430), .A2(KEYINPUT72), .A3(G125), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT16), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT73), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n457), .A2(new_n458), .A3(G146), .A4(new_n433), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n440), .A2(new_n452), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT74), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT74), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n440), .A2(new_n452), .A3(new_n462), .A4(new_n459), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n442), .B1(new_n449), .B2(new_n450), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G110), .ZN(new_n466));
  INV_X1    g280(.A(new_n445), .ZN(new_n467));
  INV_X1    g281(.A(new_n446), .ZN(new_n468));
  INV_X1    g282(.A(new_n441), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n457), .A2(new_n433), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n210), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n471), .B1(new_n473), .B2(new_n439), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n464), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n280), .A2(G221), .A3(G234), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT22), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n478), .B(new_n194), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n479), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n464), .A2(new_n475), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n302), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT75), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(KEYINPUT25), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n481), .B1(new_n464), .B2(new_n475), .ZN(new_n488));
  AOI211_X1 g302(.A(new_n479), .B(new_n474), .C1(new_n461), .C2(new_n463), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n302), .A3(new_n485), .ZN(new_n491));
  INV_X1    g305(.A(G217), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n492), .B1(new_n302), .B2(G234), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n487), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n493), .A2(G902), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(KEYINPUT76), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT77), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n494), .A2(new_n498), .A3(KEYINPUT77), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n381), .A2(new_n280), .A3(G214), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT85), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n381), .A2(new_n280), .A3(KEYINPUT85), .A4(G214), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n216), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT86), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n504), .A2(new_n216), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n506), .A2(KEYINPUT86), .A3(new_n216), .A4(new_n507), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G131), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n510), .A2(new_n201), .A3(new_n511), .A4(new_n512), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n473), .A2(new_n439), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n513), .A2(KEYINPUT17), .A3(G131), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(G113), .B(G122), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(new_n221), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n253), .A2(new_n435), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n456), .B2(new_n210), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(new_n201), .ZN(new_n526));
  OAI221_X1 g340(.A(new_n524), .B1(new_n526), .B2(new_n513), .C1(new_n514), .C2(new_n525), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n520), .A2(new_n522), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n522), .B1(new_n520), .B2(new_n527), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n313), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT89), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT89), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n532), .B(new_n313), .C1(new_n528), .C2(new_n529), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(G475), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(G475), .A2(G902), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n514), .A2(new_n516), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT87), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT19), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT88), .B1(new_n435), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n456), .B2(new_n538), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n437), .A2(KEYINPUT88), .A3(KEYINPUT19), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n253), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n543), .A2(new_n440), .A3(new_n459), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT87), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n514), .A2(new_n545), .A3(new_n516), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n537), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n522), .B1(new_n547), .B2(new_n527), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n535), .B1(new_n548), .B2(new_n528), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT20), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT20), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n551), .B(new_n535), .C1(new_n548), .C2(new_n528), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(G128), .B(G143), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(new_n192), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT90), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n554), .A2(new_n192), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT90), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n192), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(G116), .B(G122), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(new_n234), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G116), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(KEYINPUT14), .A3(G122), .ZN(new_n566));
  OAI211_X1 g380(.A(G107), .B(new_n566), .C1(new_n562), .C2(KEYINPUT14), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n556), .A2(new_n560), .A3(new_n564), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n554), .A2(KEYINPUT13), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n216), .A2(G128), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n569), .B(G134), .C1(KEYINPUT13), .C2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n234), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(new_n561), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n571), .B(new_n559), .C1(new_n573), .C2(new_n563), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n187), .A2(new_n492), .A3(G953), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n568), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n575), .B1(new_n568), .B2(new_n574), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n302), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT91), .ZN(new_n580));
  INV_X1    g394(.A(G478), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(KEYINPUT15), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n568), .A2(new_n574), .ZN(new_n583));
  INV_X1    g397(.A(new_n575), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n576), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT91), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n587), .A3(new_n302), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n580), .A2(new_n582), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT92), .ZN(new_n590));
  OR3_X1    g404(.A1(new_n579), .A2(new_n590), .A3(new_n582), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n590), .B1(new_n579), .B2(new_n582), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n589), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT21), .B(G898), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT94), .ZN(new_n596));
  NAND2_X1  g410(.A1(G234), .A2(G237), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n301), .A2(G953), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(KEYINPUT93), .B(G952), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(G953), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n597), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  AND4_X1   g417(.A1(new_n534), .A2(new_n553), .A3(new_n594), .A4(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n368), .A2(new_n429), .A3(new_n503), .A4(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  NAND2_X1  g420(.A1(new_n399), .A2(new_n302), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(G472), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n401), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n315), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n553), .A2(new_n534), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT95), .B(KEYINPUT33), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n586), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n586), .B1(KEYINPUT95), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n613), .A2(G478), .A3(new_n302), .A4(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n580), .A2(new_n581), .A3(new_n588), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n611), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n316), .B(new_n603), .C1(new_n364), .C2(new_n366), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n610), .A2(new_n622), .A3(new_n503), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT34), .B(G104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  INV_X1    g439(.A(KEYINPUT96), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n549), .B2(KEYINPUT20), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n553), .B2(new_n626), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n534), .A2(new_n593), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n621), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(new_n610), .A3(new_n503), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT35), .B(G107), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT97), .B(KEYINPUT98), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  INV_X1    g449(.A(new_n609), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n479), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n476), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n497), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n494), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n368), .A2(new_n604), .A3(new_n636), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT37), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(new_n448), .ZN(G12));
  AND2_X1   g457(.A1(new_n494), .A2(new_n639), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n405), .B2(new_n428), .ZN(new_n645));
  INV_X1    g459(.A(G900), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n598), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n602), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n628), .A2(new_n629), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n368), .A2(new_n645), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  NAND2_X1  g466(.A1(new_n611), .A2(new_n593), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n648), .B(KEYINPUT39), .Z(new_n654));
  NOR2_X1   g468(.A1(new_n315), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n352), .A2(new_n363), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n365), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n352), .A2(new_n317), .A3(new_n363), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT38), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n423), .A2(new_n395), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n386), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n386), .A2(new_n664), .A3(KEYINPUT99), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n313), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(G472), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n640), .B1(new_n405), .B2(new_n670), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n316), .B(new_n671), .C1(new_n655), .C2(new_n656), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n663), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT100), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n663), .A2(new_n676), .A3(new_n673), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n216), .ZN(G45));
  AOI211_X1 g493(.A(new_n649), .B(new_n618), .C1(new_n534), .C2(new_n553), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n368), .A2(new_n645), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  AOI21_X1  g496(.A(KEYINPUT81), .B1(new_n278), .B2(new_n283), .ZN(new_n683));
  AOI211_X1 g497(.A(new_n285), .B(new_n282), .C1(new_n268), .C2(new_n277), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n309), .A2(new_n304), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(G469), .B1(new_n686), .B2(new_n301), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n190), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n622), .A2(new_n429), .A3(new_n503), .A4(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT41), .B(G113), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT101), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n691), .B(new_n693), .ZN(G15));
  NAND4_X1  g508(.A1(new_n630), .A2(new_n429), .A3(new_n503), .A4(new_n690), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  NOR2_X1   g510(.A1(new_n689), .A2(new_n367), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n645), .A2(new_n604), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  NOR2_X1   g513(.A1(new_n653), .A2(new_n621), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n701), .B1(new_n607), .B2(G472), .ZN(new_n702));
  INV_X1    g516(.A(G472), .ZN(new_n703));
  AOI211_X1 g517(.A(KEYINPUT102), .B(new_n703), .C1(new_n399), .C2(new_n302), .ZN(new_n704));
  INV_X1    g518(.A(new_n400), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n387), .A2(new_n398), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n421), .A2(new_n425), .A3(new_n393), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n395), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n705), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n702), .A2(new_n704), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n499), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n700), .A2(new_n710), .A3(new_n711), .A4(new_n690), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  NAND4_X1  g527(.A1(new_n710), .A2(new_n697), .A3(new_n680), .A4(new_n640), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G125), .ZN(G27));
  NAND3_X1  g529(.A1(new_n659), .A2(new_n316), .A3(new_n660), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n315), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(new_n429), .A3(new_n503), .A4(new_n680), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n316), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n364), .A2(new_n366), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n300), .A2(new_n313), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n282), .B1(new_n297), .B2(new_n277), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n277), .A2(new_n306), .A3(new_n282), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n306), .B1(new_n277), .B2(new_n282), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n724), .B1(new_n727), .B2(new_n268), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n723), .B1(new_n728), .B2(G469), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n189), .B1(new_n729), .B2(new_n688), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n618), .B1(new_n553), .B2(new_n534), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n722), .A2(new_n730), .A3(new_n731), .A4(new_n648), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(KEYINPUT42), .A3(new_n429), .A4(new_n711), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n720), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G131), .ZN(G33));
  NAND4_X1  g550(.A1(new_n717), .A2(new_n650), .A3(new_n429), .A4(new_n503), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G134), .ZN(G36));
  AND2_X1   g552(.A1(new_n553), .A2(new_n534), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n619), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT43), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n609), .A3(new_n640), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n716), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n312), .B(KEYINPUT45), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(G469), .ZN(new_n747));
  INV_X1    g561(.A(new_n723), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(KEYINPUT46), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n750), .B(G469), .C1(new_n746), .C2(G902), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n688), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n190), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n654), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n745), .B(new_n754), .C1(new_n744), .C2(new_n743), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G137), .ZN(G39));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n753), .B1(new_n757), .B2(KEYINPUT47), .ZN(new_n758));
  INV_X1    g572(.A(new_n429), .ZN(new_n759));
  XNOR2_X1  g573(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n752), .A2(new_n190), .A3(new_n761), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n503), .A2(new_n620), .A3(new_n649), .A4(new_n716), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n758), .A2(new_n759), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G140), .ZN(G42));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n553), .A2(new_n534), .A3(new_n593), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n721), .B1(new_n659), .B2(new_n660), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT107), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n769), .A2(new_n770), .A3(new_n771), .A4(new_n603), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT107), .B1(new_n621), .B2(new_n768), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n772), .A2(new_n610), .A3(new_n773), .A4(new_n503), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(new_n605), .A3(new_n641), .A4(new_n623), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n695), .A2(new_n691), .A3(new_n712), .A4(new_n698), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n608), .A2(KEYINPUT102), .ZN(new_n779));
  INV_X1    g593(.A(new_n709), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n607), .A2(new_n701), .A3(G472), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n779), .A2(new_n640), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n732), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT68), .B1(new_n417), .B2(new_n412), .ZN(new_n784));
  AND4_X1   g598(.A1(KEYINPUT68), .A2(new_n410), .A3(new_n411), .A4(new_n412), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n427), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n703), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n399), .A2(new_n403), .A3(new_n400), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n403), .B1(new_n399), .B2(new_n400), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n494), .A2(KEYINPUT77), .A3(new_n498), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT77), .B1(new_n494), .B2(new_n498), .ZN(new_n793));
  OAI22_X1  g607(.A1(new_n788), .A2(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n722), .A2(new_n730), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n783), .B1(new_n796), .B2(new_n650), .ZN(new_n797));
  NOR4_X1   g611(.A1(new_n364), .A2(new_n366), .A3(new_n721), .A4(new_n649), .ZN(new_n798));
  INV_X1    g612(.A(new_n628), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n534), .A2(new_n594), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n798), .A2(new_n799), .A3(KEYINPUT108), .A4(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT108), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT96), .B1(new_n550), .B2(new_n552), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n534), .B(new_n594), .C1(new_n803), .C2(new_n627), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n659), .A2(new_n316), .A3(new_n660), .A4(new_n648), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n801), .A2(new_n806), .A3(new_n730), .A4(new_n645), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n778), .B1(new_n797), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n782), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n733), .A2(new_n809), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n778), .A2(new_n807), .A3(new_n737), .A4(new_n810), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n735), .B(new_n777), .C1(new_n808), .C2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n670), .B1(new_n789), .B2(new_n790), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n594), .B1(new_n553), .B2(new_n534), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n770), .A3(new_n644), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n730), .A2(new_n648), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT110), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n653), .A2(new_n367), .ZN(new_n818));
  AOI211_X1 g632(.A(new_n189), .B(new_n649), .C1(new_n729), .C2(new_n688), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT110), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n818), .A2(new_n671), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n368), .B(new_n645), .C1(new_n650), .C2(new_n680), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n714), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT52), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n824), .A2(new_n714), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n822), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n767), .B1(new_n812), .B2(new_n830), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n828), .A2(new_n822), .A3(new_n714), .A4(new_n824), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n828), .B1(new_n827), .B2(new_n822), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n807), .A2(new_n737), .A3(new_n810), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT109), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n797), .A2(new_n778), .A3(new_n807), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n720), .A2(new_n734), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n839), .A2(new_n775), .A3(new_n776), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n834), .A2(KEYINPUT53), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n766), .B1(new_n831), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT111), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n831), .A2(new_n841), .A3(new_n766), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT112), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n831), .A2(new_n841), .A3(new_n847), .A4(new_n766), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n740), .B(KEYINPUT43), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n602), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n689), .A2(new_n716), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n759), .A2(new_n499), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT48), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n852), .A2(new_n503), .ZN(new_n858));
  OR3_X1    g672(.A1(new_n858), .A2(new_n602), .A3(new_n813), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n731), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n710), .A2(new_n711), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n851), .A2(new_n697), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n601), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n861), .A2(KEYINPUT114), .A3(new_n601), .A4(new_n863), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n857), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT115), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n855), .A2(new_n856), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n869), .B1(new_n868), .B2(new_n870), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n758), .A2(new_n762), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n687), .A2(new_n688), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT113), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n874), .B1(new_n190), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(new_n862), .A3(new_n722), .A4(new_n851), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n662), .A2(new_n316), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n851), .A2(new_n690), .A3(new_n862), .A4(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT50), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n880), .B(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n860), .A2(new_n739), .A3(new_n618), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n853), .A2(new_n809), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n878), .A2(new_n882), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT51), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n844), .A2(new_n849), .A3(new_n873), .A4(new_n886), .ZN(new_n887));
  OR2_X1    g701(.A1(G952), .A2(G953), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n740), .A2(new_n499), .A3(new_n189), .A4(new_n721), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT105), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n875), .A2(KEYINPUT49), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n813), .B(new_n662), .C1(new_n893), .C2(KEYINPUT106), .ZN(new_n894));
  OAI221_X1 g708(.A(new_n894), .B1(KEYINPUT106), .B2(new_n893), .C1(KEYINPUT49), .C2(new_n875), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n889), .A2(new_n895), .ZN(G75));
  AOI21_X1  g710(.A(new_n302), .B1(new_n831), .B2(new_n841), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT56), .B1(new_n897), .B2(new_n365), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n345), .A2(new_n347), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(new_n329), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT116), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT55), .Z(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  OR3_X1    g717(.A1(new_n898), .A2(KEYINPUT117), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n280), .A2(G952), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT118), .Z(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n898), .B2(KEYINPUT117), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n903), .B1(new_n898), .B2(KEYINPUT117), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n904), .A2(new_n907), .A3(new_n908), .ZN(G51));
  XOR2_X1   g723(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n723), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n910), .A2(new_n723), .ZN(new_n912));
  INV_X1    g726(.A(new_n845), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n911), .B(new_n912), .C1(new_n913), .C2(new_n842), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n299), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n897), .A2(G469), .A3(new_n746), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n905), .B1(new_n915), .B2(new_n916), .ZN(G54));
  NAND3_X1  g731(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n548), .A2(new_n528), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n905), .ZN(new_n921));
  INV_X1    g735(.A(new_n919), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .A4(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(G60));
  AND2_X1   g740(.A1(new_n613), .A2(new_n615), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n831), .A2(new_n841), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT54), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n843), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n842), .A2(KEYINPUT111), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n930), .A2(new_n931), .A3(new_n846), .A4(new_n848), .ZN(new_n932));
  NAND2_X1  g746(.A1(G478), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT59), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n927), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n927), .B(new_n934), .C1(new_n913), .C2(new_n842), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n935), .A2(new_n906), .A3(new_n937), .ZN(G63));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT60), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n928), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n490), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n906), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OR2_X1    g757(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n638), .B(KEYINPUT121), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n928), .A2(new_n940), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G66));
  INV_X1    g763(.A(new_n318), .ZN(new_n950));
  OAI21_X1  g764(.A(G953), .B1(new_n596), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n777), .B2(G953), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n899), .B1(G898), .B2(new_n280), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(G69));
  NAND2_X1  g768(.A1(new_n407), .A2(new_n408), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(new_n542), .Z(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(G900), .B2(G953), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n754), .A2(new_n854), .A3(new_n818), .ZN(new_n958));
  AOI22_X1  g772(.A1(new_n958), .A2(KEYINPUT125), .B1(new_n650), .B2(new_n796), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(KEYINPUT125), .ZN(new_n960));
  INV_X1    g774(.A(new_n764), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n960), .A2(new_n961), .A3(new_n839), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT124), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n755), .A2(new_n963), .A3(new_n827), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n963), .B1(new_n755), .B2(new_n827), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n959), .B(new_n962), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n957), .B1(new_n966), .B2(G953), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n280), .B1(G227), .B2(G900), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n654), .B1(new_n620), .B2(new_n768), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n796), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT123), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n972), .A2(KEYINPUT123), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n755), .A2(new_n764), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n678), .B2(new_n825), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n675), .A2(KEYINPUT62), .A3(new_n677), .A4(new_n827), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n956), .B1(new_n979), .B2(G953), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n967), .A2(new_n970), .A3(new_n980), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n968), .A2(new_n969), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(G72));
  NAND2_X1  g797(.A1(new_n416), .A2(new_n383), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n416), .A2(new_n383), .ZN(new_n985));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n928), .A2(new_n984), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n988), .B1(new_n979), .B2(new_n777), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n921), .B(new_n990), .C1(new_n991), .C2(new_n984), .ZN(new_n992));
  INV_X1    g806(.A(new_n777), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n987), .B1(new_n966), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT127), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n992), .B1(new_n996), .B2(new_n985), .ZN(G57));
endmodule


