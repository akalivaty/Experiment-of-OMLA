//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997, new_n998;
  AND2_X1   g000(.A1(KEYINPUT87), .A2(G36gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(KEYINPUT87), .A2(G36gat), .ZN(new_n203));
  OAI21_X1  g002(.A(G29gat), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT88), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT14), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT88), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n213), .B(G29gat), .C1(new_n202), .C2(new_n203), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n205), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G43gat), .A2(G50gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(G43gat), .A2(G50gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT15), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT90), .ZN(new_n222));
  INV_X1    g021(.A(G43gat), .ZN(new_n223));
  INV_X1    g022(.A(G50gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(new_n216), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT89), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n211), .A2(new_n222), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n212), .A2(KEYINPUT90), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n225), .A2(KEYINPUT89), .A3(new_n226), .A4(new_n216), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n205), .A2(new_n219), .A3(new_n214), .A4(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n221), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT17), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G22gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G15gat), .ZN(new_n238));
  INV_X1    g037(.A(G15gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G22gat), .ZN(new_n240));
  INV_X1    g039(.A(G1gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT16), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n238), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT91), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G15gat), .B(G22gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(G1gat), .ZN(new_n247));
  OAI21_X1  g046(.A(G8gat), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n238), .A2(new_n240), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n241), .ZN(new_n250));
  INV_X1    g049(.A(G8gat), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n250), .A2(new_n244), .A3(new_n251), .A4(new_n243), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT87), .B(G36gat), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n213), .B1(new_n255), .B2(G29gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n214), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n219), .A2(new_n232), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n258), .A2(new_n230), .A3(new_n229), .A4(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(KEYINPUT17), .A3(new_n221), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n236), .A2(new_n254), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G229gat), .A2(G233gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n234), .A2(new_n253), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n263), .B(KEYINPUT13), .Z(new_n266));
  NOR2_X1   g065(.A1(new_n234), .A2(new_n253), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n260), .A2(new_n221), .B1(new_n248), .B2(new_n252), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT93), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n260), .A3(new_n221), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n264), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT93), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n273), .A3(new_n266), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n265), .A2(KEYINPUT18), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT18), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G113gat), .B(G141gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(G197gat), .ZN(new_n280));
  XOR2_X1   g079(.A(KEYINPUT11), .B(G169gat), .Z(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT12), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n275), .B(new_n278), .C1(KEYINPUT92), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n270), .A2(new_n274), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n262), .A2(KEYINPUT18), .A3(new_n263), .A4(new_n264), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n278), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n273), .B1(new_n272), .B2(new_n266), .ZN(new_n288));
  INV_X1    g087(.A(new_n266), .ZN(new_n289));
  AOI211_X1 g088(.A(KEYINPUT93), .B(new_n289), .C1(new_n271), .C2(new_n264), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n286), .B(KEYINPUT92), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n283), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n287), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n284), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G227gat), .ZN(new_n295));
  INV_X1    g094(.A(G233gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(KEYINPUT64), .B(G190gat), .Z(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT27), .B(G183gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT28), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT66), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n300), .B(new_n302), .Z(new_n303));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  NOR3_X1   g106(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT26), .ZN(new_n308));
  AOI211_X1 g107(.A(new_n305), .B(new_n308), .C1(KEYINPUT26), .C2(new_n307), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n304), .B(KEYINPUT24), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n311), .B1(G183gat), .B2(G190gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n313), .B1(G169gat), .B2(G176gat), .ZN(new_n314));
  MUX2_X1   g113(.A(new_n314), .B(new_n313), .S(new_n307), .Z(new_n315));
  NAND2_X1  g114(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT25), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G183gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n298), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n311), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(new_n315), .A3(KEYINPUT25), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(KEYINPUT65), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT65), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(new_n318), .B2(new_n322), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n310), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT1), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n328), .B1(G113gat), .B2(G120gat), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(G113gat), .B2(G120gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(G127gat), .B(G134gat), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n329), .ZN(new_n333));
  XOR2_X1   g132(.A(KEYINPUT67), .B(G113gat), .Z(new_n334));
  INV_X1    g133(.A(G120gat), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n331), .B(new_n333), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n327), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n337), .B(new_n310), .C1(new_n324), .C2(new_n326), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n297), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n340), .ZN(new_n344));
  INV_X1    g143(.A(new_n297), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n345), .A3(new_n342), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n339), .A2(new_n297), .A3(new_n340), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT32), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT33), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G15gat), .B(G43gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT68), .ZN(new_n353));
  INV_X1    g152(.A(G71gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G99gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n349), .A2(new_n351), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n357), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n348), .B(KEYINPUT32), .C1(new_n350), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n347), .A2(new_n361), .A3(KEYINPUT70), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n347), .B1(new_n361), .B2(KEYINPUT70), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT36), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT36), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n343), .A2(new_n346), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n361), .A2(new_n367), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G155gat), .B(G162gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT75), .ZN(new_n375));
  XNOR2_X1  g174(.A(G141gat), .B(G148gat), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT76), .B(G162gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G155gat), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT2), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n377), .B(new_n381), .C1(new_n375), .C2(new_n376), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n374), .B1(KEYINPUT2), .B2(new_n376), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n338), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT4), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT77), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n338), .B1(new_n384), .B2(new_n387), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n382), .A2(new_n383), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT77), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT3), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n388), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(KEYINPUT78), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT78), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n337), .B1(new_n390), .B2(KEYINPUT3), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n391), .B1(new_n390), .B2(KEYINPUT3), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n395), .B1(new_n398), .B2(new_n392), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n372), .B(new_n386), .C1(new_n394), .C2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n390), .B(new_n338), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT5), .B1(new_n401), .B2(new_n372), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n385), .B(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n393), .A2(KEYINPUT78), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n398), .A2(new_n395), .A3(new_n392), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(KEYINPUT5), .A3(new_n372), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G1gat), .B(G29gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT0), .ZN(new_n412));
  XNOR2_X1  g211(.A(G57gat), .B(G85gat), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n412), .B(new_n413), .Z(new_n414));
  NAND2_X1  g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT80), .ZN(new_n416));
  XOR2_X1   g215(.A(KEYINPUT79), .B(KEYINPUT6), .Z(new_n417));
  INV_X1    g216(.A(new_n414), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n418), .A3(new_n409), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n415), .A2(new_n416), .A3(new_n417), .A4(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G8gat), .B(G36gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(G64gat), .B(G92gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n421), .B(new_n422), .Z(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT71), .B(G197gat), .ZN(new_n425));
  INV_X1    g224(.A(G204gat), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n425), .A2(new_n426), .ZN(new_n428));
  INV_X1    g227(.A(G211gat), .ZN(new_n429));
  INV_X1    g228(.A(G218gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI22_X1  g230(.A1(new_n427), .A2(new_n428), .B1(KEYINPUT22), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT72), .ZN(new_n433));
  XOR2_X1   g232(.A(G211gat), .B(G218gat), .Z(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n433), .A2(new_n435), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n310), .A2(new_n323), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT73), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G226gat), .A2(G233gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n443), .A2(KEYINPUT29), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n310), .A2(KEYINPUT73), .A3(new_n323), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n443), .B(new_n310), .C1(new_n324), .C2(new_n326), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n438), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT74), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n327), .A2(new_n444), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n441), .A2(new_n445), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n438), .B(new_n451), .C1(new_n452), .C2(new_n442), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n448), .A2(new_n449), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n424), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n446), .A2(new_n447), .ZN(new_n457));
  INV_X1    g256(.A(new_n438), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT74), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n460), .A2(new_n450), .A3(new_n453), .A4(new_n423), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n456), .A2(KEYINPUT30), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n454), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT30), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n463), .A2(new_n464), .A3(new_n460), .A4(new_n423), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n403), .A2(new_n418), .A3(new_n409), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n418), .B1(new_n403), .B2(new_n409), .ZN(new_n468));
  INV_X1    g267(.A(new_n417), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n403), .A2(new_n409), .A3(new_n418), .A4(new_n469), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT80), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n420), .B(new_n466), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT29), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n436), .A2(new_n437), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n387), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n390), .ZN(new_n477));
  NAND2_X1  g276(.A1(G228gat), .A2(G233gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n474), .B1(new_n390), .B2(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n438), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n384), .B1(new_n475), .B2(new_n387), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n438), .A2(new_n480), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n478), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n485), .A3(new_n237), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT81), .ZN(new_n487));
  XOR2_X1   g286(.A(G78gat), .B(G106gat), .Z(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT31), .B(G50gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n482), .A2(new_n485), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G22gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n486), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT81), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n493), .A2(new_n496), .A3(new_n486), .A4(new_n490), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n473), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n371), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT82), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n371), .A2(new_n499), .A3(KEYINPUT82), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT86), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n410), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n403), .A2(KEYINPUT86), .A3(new_n409), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n418), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n468), .A2(new_n469), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n507), .A2(new_n508), .B1(new_n469), .B2(new_n467), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT37), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n460), .A2(new_n510), .A3(new_n450), .A4(new_n453), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n457), .B2(new_n438), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n458), .B(new_n451), .C1(new_n452), .C2(new_n442), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT38), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n424), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n461), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT37), .B1(new_n454), .B2(new_n455), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(new_n424), .A3(new_n511), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n516), .B1(KEYINPUT38), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n509), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n497), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n487), .A2(new_n490), .B1(new_n493), .B2(new_n486), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n408), .A2(new_n372), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT83), .B(KEYINPUT39), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n418), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(KEYINPUT85), .A2(KEYINPUT40), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n401), .A2(new_n372), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT39), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n529), .A2(KEYINPUT84), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(KEYINPUT84), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n530), .B(new_n531), .C1(new_n372), .C2(new_n408), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n526), .A2(new_n527), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n527), .B1(new_n526), .B2(new_n532), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n507), .A2(new_n465), .A3(new_n462), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n520), .B(new_n523), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n502), .A2(new_n503), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n361), .A2(KEYINPUT70), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n367), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n495), .A2(new_n497), .A3(new_n540), .A4(new_n362), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT35), .B1(new_n473), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n507), .A2(new_n508), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n471), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT35), .ZN(new_n545));
  INV_X1    g344(.A(new_n369), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n361), .A2(new_n367), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n546), .A2(new_n547), .B1(new_n462), .B2(new_n465), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n544), .A2(new_n545), .A3(new_n523), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n542), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n294), .B1(new_n538), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G183gat), .B(G211gat), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n553));
  INV_X1    g352(.A(G57gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(G64gat), .ZN(new_n555));
  INV_X1    g354(.A(G64gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(G57gat), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n553), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(G71gat), .A2(G78gat), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT94), .ZN(new_n561));
  NAND2_X1  g360(.A1(G71gat), .A2(G78gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n562), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT94), .B1(new_n564), .B2(new_n559), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n558), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n560), .A2(new_n562), .ZN(new_n567));
  XNOR2_X1  g366(.A(G57gat), .B(G64gat), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n567), .B(KEYINPUT94), .C1(new_n568), .C2(new_n553), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT21), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(G127gat), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n566), .A2(new_n569), .A3(new_n570), .A4(new_n572), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n575), .B1(new_n574), .B2(new_n576), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n552), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n574), .A2(new_n576), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(G127gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n552), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n582), .A2(new_n583), .A3(new_n577), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(new_n380), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n570), .B1(new_n566), .B2(new_n569), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT95), .B1(new_n253), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n253), .A2(new_n587), .A3(KEYINPUT95), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n566), .A2(new_n569), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n254), .B(new_n592), .C1(new_n570), .C2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n586), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n588), .A3(new_n596), .ZN(new_n597));
  AND4_X1   g396(.A1(new_n580), .A2(new_n584), .A3(new_n591), .A4(new_n597), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n580), .A2(new_n584), .B1(new_n591), .B2(new_n597), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n605));
  XOR2_X1   g404(.A(G99gat), .B(G106gat), .Z(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT96), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(KEYINPUT7), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(KEYINPUT7), .ZN(new_n610));
  AND2_X1   g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT97), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n612), .B1(new_n610), .B2(new_n611), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n609), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT7), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n616), .A2(KEYINPUT96), .ZN(new_n617));
  NAND2_X1  g416(.A1(G85gat), .A2(G92gat), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT97), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n609), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G99gat), .A2(G106gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT8), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(G85gat), .B2(G92gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n607), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  AOI211_X1 g427(.A(new_n606), .B(new_n626), .C1(new_n615), .C2(new_n622), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n605), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n620), .B1(new_n619), .B2(new_n621), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n627), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n606), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n623), .A2(new_n607), .A3(new_n627), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(KEYINPUT98), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n630), .A2(new_n636), .A3(new_n261), .A4(new_n236), .ZN(new_n637));
  XNOR2_X1  g436(.A(G190gat), .B(G218gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT99), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AND3_X1   g439(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n628), .A2(new_n629), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n641), .B1(new_n642), .B2(new_n234), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n637), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n640), .B1(new_n637), .B2(new_n643), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n604), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n637), .A2(new_n643), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n639), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n637), .A2(new_n640), .A3(new_n643), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(new_n603), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n600), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n653), .B(new_n654), .Z(new_n655));
  OAI21_X1  g454(.A(new_n594), .B1(new_n628), .B2(new_n629), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n634), .A2(new_n593), .A3(new_n635), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT100), .B(KEYINPUT10), .Z(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n642), .A2(KEYINPUT10), .A3(new_n593), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(G230gat), .A2(G233gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(new_n656), .B2(new_n657), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n655), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n662), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n667), .B1(new_n659), .B2(new_n660), .ZN(new_n668));
  INV_X1    g467(.A(new_n655), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n668), .A2(new_n664), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n652), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n551), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n420), .B1(new_n470), .B2(new_n472), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(new_n241), .ZN(G1324gat));
  INV_X1    g477(.A(new_n674), .ZN(new_n679));
  INV_X1    g478(.A(new_n466), .ZN(new_n680));
  NOR2_X1   g479(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT16), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n679), .A2(new_n251), .A3(new_n680), .A4(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n551), .A2(new_n680), .A3(new_n673), .ZN(new_n685));
  OAI21_X1  g484(.A(G8gat), .B1(new_n685), .B2(new_n682), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n684), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n684), .A2(KEYINPUT102), .A3(new_n686), .A4(new_n688), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1325gat));
  OAI21_X1  g492(.A(G15gat), .B1(new_n674), .B2(new_n371), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n368), .A2(new_n369), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n239), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n694), .B1(new_n674), .B2(new_n697), .ZN(G1326gat));
  OR3_X1    g497(.A1(new_n674), .A2(KEYINPUT103), .A3(new_n523), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT103), .B1(new_n674), .B2(new_n523), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT43), .B(G22gat), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n699), .B2(new_n700), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(G1327gat));
  INV_X1    g503(.A(new_n600), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n672), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n646), .A2(new_n650), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  AOI211_X1 g510(.A(new_n294), .B(new_n711), .C1(new_n538), .C2(new_n550), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(new_n206), .A3(new_n675), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT45), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n365), .A2(new_n370), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n473), .B2(new_n498), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n537), .B1(new_n717), .B2(KEYINPUT82), .ZN(new_n718));
  INV_X1    g517(.A(new_n503), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n550), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n709), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n509), .A2(new_n519), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n523), .B1(new_n536), .B2(new_n535), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n550), .B1(new_n726), .B2(new_n500), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n708), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n721), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n707), .A2(new_n294), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n723), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n715), .B1(new_n731), .B2(new_n676), .ZN(new_n732));
  INV_X1    g531(.A(new_n722), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n733), .B1(new_n538), .B2(new_n550), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT44), .B1(new_n727), .B2(new_n708), .ZN(new_n735));
  INV_X1    g534(.A(new_n730), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n737), .A2(KEYINPUT104), .A3(new_n675), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n732), .A2(new_n738), .A3(G29gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n714), .A2(new_n739), .ZN(G1328gat));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n466), .A2(new_n255), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n712), .A2(new_n742), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n284), .A2(new_n293), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n720), .A2(new_n746), .A3(new_n710), .A4(new_n744), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT105), .B1(new_n747), .B2(KEYINPUT46), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(KEYINPUT46), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n734), .A2(new_n735), .A3(new_n466), .A4(new_n736), .ZN(new_n751));
  INV_X1    g550(.A(new_n255), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n741), .B1(new_n749), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n745), .A2(new_n748), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n255), .B1(new_n731), .B2(new_n466), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n755), .A2(KEYINPUT106), .A3(new_n756), .A4(new_n750), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(G1329gat));
  OAI21_X1  g557(.A(G43gat), .B1(new_n731), .B2(new_n371), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n712), .A2(new_n223), .A3(new_n696), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n731), .B2(new_n371), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n737), .A2(KEYINPUT107), .A3(new_n716), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n765), .A2(new_n766), .A3(G43gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n760), .A2(KEYINPUT47), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n763), .B1(new_n767), .B2(new_n768), .ZN(G1330gat));
  INV_X1    g568(.A(KEYINPUT48), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n523), .A2(G50gat), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n720), .A2(new_n746), .A3(new_n710), .A4(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n224), .B1(new_n737), .B2(new_n498), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n770), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n731), .B2(new_n523), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n737), .A2(KEYINPUT109), .A3(new_n498), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n778), .A2(new_n779), .A3(G50gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n772), .A2(KEYINPUT48), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(G1331gat));
  NOR3_X1   g581(.A1(new_n652), .A2(new_n746), .A3(new_n671), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n727), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n676), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(new_n554), .ZN(G1332gat));
  INV_X1    g585(.A(KEYINPUT110), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n784), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n680), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n790));
  XOR2_X1   g589(.A(KEYINPUT49), .B(G64gat), .Z(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n789), .B2(new_n791), .ZN(G1333gat));
  NAND3_X1  g591(.A1(new_n788), .A2(G71gat), .A3(new_n716), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n695), .B(KEYINPUT111), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n354), .B1(new_n784), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g596(.A1(new_n788), .A2(new_n498), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g598(.A1(new_n746), .A2(new_n705), .A3(new_n671), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n723), .A2(new_n729), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(G85gat), .B1(new_n801), .B2(new_n676), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n746), .A2(new_n705), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n727), .A2(new_n708), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n727), .A2(KEYINPUT51), .A3(new_n708), .A4(new_n803), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  OR3_X1    g608(.A1(new_n676), .A2(G85gat), .A3(new_n671), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n802), .B1(new_n809), .B2(new_n810), .ZN(G1336gat));
  OAI21_X1  g610(.A(KEYINPUT113), .B1(new_n801), .B2(new_n466), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n734), .A2(new_n735), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n813), .A2(new_n814), .A3(new_n680), .A4(new_n800), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(G92gat), .A3(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n466), .A2(G92gat), .A3(new_n671), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT52), .B1(new_n808), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n806), .A2(new_n820), .A3(new_n807), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n821), .B(new_n817), .C1(new_n820), .C2(new_n806), .ZN(new_n822));
  OAI21_X1  g621(.A(G92gat), .B1(new_n801), .B2(new_n466), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT52), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n819), .A2(new_n825), .ZN(G1337gat));
  OAI21_X1  g625(.A(G99gat), .B1(new_n801), .B2(new_n371), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n695), .A2(G99gat), .A3(new_n671), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT114), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n809), .B2(new_n829), .ZN(G1338gat));
  NOR3_X1   g629(.A1(new_n523), .A2(G106gat), .A3(new_n671), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n821), .B(new_n831), .C1(new_n820), .C2(new_n806), .ZN(new_n832));
  OAI21_X1  g631(.A(G106gat), .B1(new_n801), .B2(new_n523), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT53), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT53), .B1(new_n808), .B2(new_n831), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(G1339gat));
  NAND4_X1  g637(.A1(new_n651), .A2(new_n284), .A3(new_n293), .A4(new_n671), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT115), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n659), .A2(new_n667), .A3(new_n660), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n663), .A2(KEYINPUT54), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n655), .B1(new_n668), .B2(new_n843), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n842), .A2(KEYINPUT55), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT55), .B1(new_n842), .B2(new_n844), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n845), .A2(new_n846), .A3(new_n670), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n271), .A2(new_n264), .A3(new_n289), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n848), .B(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n263), .B1(new_n262), .B2(new_n264), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n282), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n285), .A2(new_n278), .A3(new_n286), .A4(new_n283), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n847), .A2(new_n708), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n853), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n671), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(new_n847), .B2(new_n746), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n855), .B1(new_n858), .B2(new_n708), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n840), .B1(new_n859), .B2(new_n600), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(new_n676), .ZN(new_n861));
  INV_X1    g660(.A(new_n541), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n680), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n334), .A3(new_n746), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n861), .A2(new_n523), .A3(new_n548), .ZN(new_n866));
  OAI21_X1  g665(.A(G113gat), .B1(new_n866), .B2(new_n294), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1340gat));
  NOR3_X1   g667(.A1(new_n866), .A2(new_n335), .A3(new_n671), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n864), .A2(new_n672), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n335), .ZN(G1341gat));
  NAND3_X1  g670(.A1(new_n864), .A2(new_n575), .A3(new_n705), .ZN(new_n872));
  OAI21_X1  g671(.A(G127gat), .B1(new_n866), .B2(new_n600), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1342gat));
  NAND2_X1  g673(.A1(new_n466), .A2(new_n708), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT117), .Z(new_n876));
  NOR3_X1   g675(.A1(new_n863), .A2(G134gat), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT56), .ZN(new_n878));
  OAI21_X1  g677(.A(G134gat), .B1(new_n866), .B2(new_n709), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1343gat));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n842), .A2(new_n844), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT55), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n670), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n842), .A2(KEYINPUT55), .A3(new_n844), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n746), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n672), .A2(new_n854), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n708), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n882), .A2(new_n883), .ZN(new_n889));
  INV_X1    g688(.A(new_n670), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n890), .A3(new_n885), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n854), .A2(new_n708), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n600), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n839), .B(new_n895), .ZN(new_n896));
  AOI211_X1 g695(.A(new_n881), .B(new_n523), .C1(new_n894), .C2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n887), .B1(new_n891), .B2(new_n294), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n893), .B1(new_n900), .B2(new_n709), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n896), .B1(new_n901), .B2(new_n705), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n498), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n899), .B1(new_n903), .B2(new_n881), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n523), .B1(new_n894), .B2(new_n896), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n905), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n898), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n676), .A2(new_n716), .A3(new_n680), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n746), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G141gat), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT58), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n905), .A2(new_n675), .A3(new_n371), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT121), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(new_n680), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n294), .A2(G141gat), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n910), .B(new_n911), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n907), .A2(KEYINPUT119), .A3(new_n908), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT118), .B1(new_n905), .B2(KEYINPUT57), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n899), .B(new_n881), .C1(new_n860), .C2(new_n523), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n897), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n908), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n918), .A2(new_n924), .A3(new_n746), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n925), .A2(new_n926), .A3(G141gat), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n926), .B1(new_n925), .B2(G141gat), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n912), .A2(new_n680), .A3(new_n916), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n917), .B1(new_n930), .B2(new_n911), .ZN(G1344gat));
  INV_X1    g730(.A(KEYINPUT59), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n918), .A2(new_n924), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n932), .B(G148gat), .C1(new_n933), .C2(new_n671), .ZN(new_n934));
  INV_X1    g733(.A(G148gat), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n523), .B1(new_n894), .B2(new_n839), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n898), .B1(KEYINPUT57), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n937), .A2(new_n672), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n935), .B1(new_n938), .B2(new_n908), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n934), .B1(new_n932), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n914), .A2(new_n935), .A3(new_n672), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1345gat));
  OAI21_X1  g741(.A(G155gat), .B1(new_n933), .B2(new_n600), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n914), .A2(new_n380), .A3(new_n705), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1346gat));
  OAI21_X1  g744(.A(new_n378), .B1(new_n933), .B2(new_n709), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n876), .A2(new_n378), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n913), .B2(new_n947), .ZN(G1347gat));
  NOR2_X1   g747(.A1(new_n675), .A2(new_n466), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n949), .A2(new_n902), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n950), .A2(new_n862), .ZN(new_n951));
  AOI21_X1  g750(.A(G169gat), .B1(new_n951), .B2(new_n746), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n794), .A2(new_n498), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(G169gat), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n954), .A2(new_n955), .A3(new_n294), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n952), .A2(new_n956), .ZN(G1348gat));
  NAND2_X1  g756(.A1(new_n672), .A2(G176gat), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT122), .ZN(new_n960));
  AOI21_X1  g759(.A(G176gat), .B1(new_n951), .B2(new_n672), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(G1349gat));
  NAND3_X1  g761(.A1(new_n951), .A2(new_n299), .A3(new_n705), .ZN(new_n963));
  OAI21_X1  g762(.A(G183gat), .B1(new_n954), .B2(new_n600), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(KEYINPUT123), .A3(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n298), .A3(new_n708), .ZN(new_n967));
  OAI21_X1  g766(.A(G190gat), .B1(new_n954), .B2(new_n709), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1351gat));
  NAND2_X1  g770(.A1(new_n371), .A2(new_n949), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n937), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n974), .A2(new_n746), .ZN(new_n975));
  OR2_X1    g774(.A1(new_n975), .A2(KEYINPUT124), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(KEYINPUT124), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n976), .A2(G197gat), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n972), .A2(new_n903), .ZN(new_n979));
  INV_X1    g778(.A(G197gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n979), .A2(new_n980), .A3(new_n746), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n978), .A2(new_n981), .ZN(G1352gat));
  AOI21_X1  g781(.A(new_n426), .B1(new_n938), .B2(new_n973), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n979), .A2(new_n426), .A3(new_n672), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n984), .B(KEYINPUT62), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n983), .A2(new_n985), .ZN(G1353gat));
  NAND2_X1  g785(.A1(new_n974), .A2(new_n705), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT63), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n429), .B1(KEYINPUT125), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT125), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n990), .A2(new_n991), .A3(KEYINPUT63), .ZN(new_n992));
  OAI211_X1 g791(.A(new_n987), .B(new_n989), .C1(KEYINPUT125), .C2(new_n988), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n979), .A2(new_n429), .A3(new_n705), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(G1354gat));
  NAND2_X1  g794(.A1(new_n974), .A2(new_n708), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n709), .A2(G218gat), .ZN(new_n997));
  AOI22_X1  g796(.A1(new_n996), .A2(G218gat), .B1(new_n979), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g797(.A(new_n998), .B(KEYINPUT126), .Z(G1355gat));
endmodule


