

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(G651), .A2(n646), .ZN(n656) );
  NOR2_X1 U551 ( .A1(n775), .A2(n517), .ZN(n776) );
  NOR2_X1 U552 ( .A1(n557), .A2(n556), .ZN(n558) );
  BUF_X1 U553 ( .A(n547), .Z(n529) );
  AND2_X2 U554 ( .A1(n523), .A2(G2104), .ZN(n894) );
  AND2_X1 U555 ( .A1(n757), .A2(n731), .ZN(n733) );
  INV_X1 U556 ( .A(G2105), .ZN(n523) );
  NOR2_X1 U557 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  XNOR2_X1 U558 ( .A(n729), .B(n728), .ZN(n757) );
  INV_X1 U559 ( .A(KEYINPUT96), .ZN(n728) );
  NOR2_X1 U560 ( .A1(n778), .A2(n768), .ZN(n775) );
  INV_X1 U561 ( .A(KEYINPUT23), .ZN(n581) );
  NAND2_X1 U562 ( .A1(n895), .A2(G137), .ZN(n579) );
  NOR2_X1 U563 ( .A1(n774), .A2(n773), .ZN(n517) );
  OR2_X1 U564 ( .A1(G301), .A2(n736), .ZN(n518) );
  NOR2_X1 U565 ( .A1(n745), .A2(n862), .ZN(n699) );
  INV_X1 U566 ( .A(KEYINPUT30), .ZN(n732) );
  INV_X1 U567 ( .A(KEYINPUT29), .ZN(n722) );
  XNOR2_X1 U568 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n740) );
  XOR2_X1 U569 ( .A(n741), .B(n740), .Z(n742) );
  NAND2_X1 U570 ( .A1(n743), .A2(n742), .ZN(n758) );
  INV_X1 U571 ( .A(KEYINPUT32), .ZN(n753) );
  INV_X1 U572 ( .A(n978), .ZN(n766) );
  XNOR2_X1 U573 ( .A(n754), .B(n753), .ZN(n762) );
  NAND2_X1 U574 ( .A1(n767), .A2(n766), .ZN(n768) );
  OR2_X2 U575 ( .A1(n806), .A2(n704), .ZN(n745) );
  OR2_X1 U576 ( .A1(n697), .A2(n696), .ZN(n806) );
  NOR2_X1 U577 ( .A1(G164), .A2(G1384), .ZN(n807) );
  INV_X1 U578 ( .A(KEYINPUT17), .ZN(n519) );
  XNOR2_X1 U579 ( .A(KEYINPUT72), .B(KEYINPUT15), .ZN(n594) );
  NOR2_X2 U580 ( .A1(G2104), .A2(n523), .ZN(n898) );
  XNOR2_X1 U581 ( .A(n595), .B(n594), .ZN(n611) );
  XNOR2_X1 U582 ( .A(n582), .B(n581), .ZN(n584) );
  NAND2_X1 U583 ( .A1(G102), .A2(n894), .ZN(n522) );
  XNOR2_X2 U584 ( .A(n520), .B(n519), .ZN(n895) );
  NAND2_X1 U585 ( .A1(G138), .A2(n895), .ZN(n521) );
  NAND2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n527) );
  AND2_X1 U587 ( .A1(G2104), .A2(G2105), .ZN(n900) );
  NAND2_X1 U588 ( .A1(G114), .A2(n900), .ZN(n525) );
  NAND2_X1 U589 ( .A1(G126), .A2(n898), .ZN(n524) );
  NAND2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(G164) );
  XOR2_X1 U592 ( .A(G543), .B(KEYINPUT0), .Z(n646) );
  INV_X1 U593 ( .A(G651), .ZN(n532) );
  NOR2_X2 U594 ( .A1(n646), .A2(n532), .ZN(n662) );
  NAND2_X1 U595 ( .A1(n662), .A2(G72), .ZN(n531) );
  NOR2_X1 U596 ( .A1(G543), .A2(G651), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n528), .B(KEYINPUT64), .ZN(n547) );
  NAND2_X1 U598 ( .A1(G85), .A2(n529), .ZN(n530) );
  NAND2_X1 U599 ( .A1(n531), .A2(n530), .ZN(n537) );
  NAND2_X1 U600 ( .A1(G47), .A2(n656), .ZN(n535) );
  NOR2_X1 U601 ( .A1(G543), .A2(n532), .ZN(n533) );
  XOR2_X2 U602 ( .A(KEYINPUT1), .B(n533), .Z(n654) );
  NAND2_X1 U603 ( .A1(G60), .A2(n654), .ZN(n534) );
  NAND2_X1 U604 ( .A1(n535), .A2(n534), .ZN(n536) );
  OR2_X1 U605 ( .A1(n537), .A2(n536), .ZN(G290) );
  INV_X1 U606 ( .A(G57), .ZN(G237) );
  XOR2_X1 U607 ( .A(G2443), .B(G2446), .Z(n539) );
  XNOR2_X1 U608 ( .A(G2427), .B(G2451), .ZN(n538) );
  XNOR2_X1 U609 ( .A(n539), .B(n538), .ZN(n545) );
  XOR2_X1 U610 ( .A(G2430), .B(G2454), .Z(n541) );
  XNOR2_X1 U611 ( .A(G1341), .B(G1348), .ZN(n540) );
  XNOR2_X1 U612 ( .A(n541), .B(n540), .ZN(n543) );
  XOR2_X1 U613 ( .A(G2435), .B(G2438), .Z(n542) );
  XNOR2_X1 U614 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U615 ( .A(n545), .B(n544), .Z(n546) );
  AND2_X1 U616 ( .A1(G14), .A2(n546), .ZN(G401) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U618 ( .A(G860), .ZN(n609) );
  NAND2_X1 U619 ( .A1(G68), .A2(n662), .ZN(n551) );
  NAND2_X1 U620 ( .A1(n547), .A2(G81), .ZN(n548) );
  XOR2_X1 U621 ( .A(KEYINPUT12), .B(n548), .Z(n549) );
  XNOR2_X1 U622 ( .A(n549), .B(KEYINPUT69), .ZN(n550) );
  NAND2_X1 U623 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U624 ( .A(n552), .B(KEYINPUT13), .ZN(n554) );
  NAND2_X1 U625 ( .A1(G43), .A2(n656), .ZN(n553) );
  NAND2_X1 U626 ( .A1(n554), .A2(n553), .ZN(n557) );
  NAND2_X1 U627 ( .A1(n654), .A2(G56), .ZN(n555) );
  XOR2_X1 U628 ( .A(KEYINPUT14), .B(n555), .Z(n556) );
  XOR2_X2 U629 ( .A(KEYINPUT70), .B(n558), .Z(n993) );
  OR2_X1 U630 ( .A1(n609), .A2(n993), .ZN(G153) );
  INV_X1 U631 ( .A(G108), .ZN(G238) );
  INV_X1 U632 ( .A(G120), .ZN(G236) );
  INV_X1 U633 ( .A(G132), .ZN(G219) );
  INV_X1 U634 ( .A(G82), .ZN(G220) );
  NAND2_X1 U635 ( .A1(G52), .A2(n656), .ZN(n560) );
  NAND2_X1 U636 ( .A1(G64), .A2(n654), .ZN(n559) );
  NAND2_X1 U637 ( .A1(n560), .A2(n559), .ZN(n565) );
  NAND2_X1 U638 ( .A1(n662), .A2(G77), .ZN(n562) );
  NAND2_X1 U639 ( .A1(G90), .A2(n529), .ZN(n561) );
  NAND2_X1 U640 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U641 ( .A(KEYINPUT9), .B(n563), .Z(n564) );
  NOR2_X1 U642 ( .A1(n565), .A2(n564), .ZN(G171) );
  INV_X1 U643 ( .A(G171), .ZN(G301) );
  NAND2_X1 U644 ( .A1(n529), .A2(G89), .ZN(n566) );
  XOR2_X1 U645 ( .A(KEYINPUT73), .B(n566), .Z(n567) );
  XNOR2_X1 U646 ( .A(n567), .B(KEYINPUT4), .ZN(n569) );
  NAND2_X1 U647 ( .A1(G76), .A2(n662), .ZN(n568) );
  NAND2_X1 U648 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U649 ( .A(n570), .B(KEYINPUT5), .ZN(n576) );
  NAND2_X1 U650 ( .A1(n656), .A2(G51), .ZN(n571) );
  XNOR2_X1 U651 ( .A(n571), .B(KEYINPUT74), .ZN(n573) );
  NAND2_X1 U652 ( .A1(G63), .A2(n654), .ZN(n572) );
  NAND2_X1 U653 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U654 ( .A(KEYINPUT6), .B(n574), .Z(n575) );
  NAND2_X1 U655 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U656 ( .A(n577), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U657 ( .A1(G113), .A2(n900), .ZN(n578) );
  NAND2_X1 U658 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U659 ( .A(n580), .B(KEYINPUT65), .Z(n697) );
  NAND2_X1 U660 ( .A1(G101), .A2(n894), .ZN(n582) );
  NAND2_X1 U661 ( .A1(G125), .A2(n898), .ZN(n583) );
  NAND2_X1 U662 ( .A1(n584), .A2(n583), .ZN(n695) );
  NOR2_X1 U663 ( .A1(n697), .A2(n695), .ZN(G160) );
  NAND2_X1 U664 ( .A1(G7), .A2(G661), .ZN(n585) );
  XNOR2_X1 U665 ( .A(n585), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U666 ( .A(G223), .B(KEYINPUT68), .Z(n844) );
  AND2_X1 U667 ( .A1(n844), .A2(G567), .ZN(n586) );
  XNOR2_X1 U668 ( .A(n586), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U669 ( .A1(n654), .A2(G66), .ZN(n588) );
  NAND2_X1 U670 ( .A1(G92), .A2(n529), .ZN(n587) );
  NAND2_X1 U671 ( .A1(n588), .A2(n587), .ZN(n593) );
  NAND2_X1 U672 ( .A1(G79), .A2(n662), .ZN(n590) );
  NAND2_X1 U673 ( .A1(G54), .A2(n656), .ZN(n589) );
  NAND2_X1 U674 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U675 ( .A(n591), .B(KEYINPUT71), .Z(n592) );
  NOR2_X1 U676 ( .A1(n593), .A2(n592), .ZN(n595) );
  NOR2_X1 U677 ( .A1(n611), .A2(G868), .ZN(n597) );
  INV_X1 U678 ( .A(G868), .ZN(n675) );
  NOR2_X1 U679 ( .A1(n675), .A2(G301), .ZN(n596) );
  NOR2_X1 U680 ( .A1(n597), .A2(n596), .ZN(G284) );
  XOR2_X1 U681 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U682 ( .A1(G53), .A2(n656), .ZN(n599) );
  NAND2_X1 U683 ( .A1(G65), .A2(n654), .ZN(n598) );
  NAND2_X1 U684 ( .A1(n599), .A2(n598), .ZN(n604) );
  NAND2_X1 U685 ( .A1(n662), .A2(G78), .ZN(n601) );
  NAND2_X1 U686 ( .A1(G91), .A2(n529), .ZN(n600) );
  NAND2_X1 U687 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U688 ( .A(KEYINPUT66), .B(n602), .ZN(n603) );
  NOR2_X1 U689 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U690 ( .A(n605), .B(KEYINPUT67), .Z(n976) );
  INV_X1 U691 ( .A(n976), .ZN(G299) );
  XOR2_X1 U692 ( .A(KEYINPUT75), .B(n675), .Z(n606) );
  NOR2_X1 U693 ( .A1(G286), .A2(n606), .ZN(n608) );
  NOR2_X1 U694 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U695 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U696 ( .A1(G559), .A2(n609), .ZN(n610) );
  XNOR2_X1 U697 ( .A(n610), .B(KEYINPUT76), .ZN(n612) );
  INV_X1 U698 ( .A(n611), .ZN(n988) );
  NAND2_X1 U699 ( .A1(n612), .A2(n988), .ZN(n613) );
  XNOR2_X1 U700 ( .A(KEYINPUT16), .B(n613), .ZN(G148) );
  NOR2_X1 U701 ( .A1(n993), .A2(G868), .ZN(n616) );
  NAND2_X1 U702 ( .A1(n988), .A2(G868), .ZN(n614) );
  NOR2_X1 U703 ( .A1(G559), .A2(n614), .ZN(n615) );
  NOR2_X1 U704 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U705 ( .A1(G111), .A2(n900), .ZN(n617) );
  XNOR2_X1 U706 ( .A(n617), .B(KEYINPUT78), .ZN(n620) );
  NAND2_X1 U707 ( .A1(G99), .A2(n894), .ZN(n618) );
  XOR2_X1 U708 ( .A(KEYINPUT79), .B(n618), .Z(n619) );
  NAND2_X1 U709 ( .A1(n620), .A2(n619), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n898), .A2(G123), .ZN(n621) );
  XNOR2_X1 U711 ( .A(n621), .B(KEYINPUT18), .ZN(n623) );
  NAND2_X1 U712 ( .A1(G135), .A2(n895), .ZN(n622) );
  NAND2_X1 U713 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U714 ( .A(KEYINPUT77), .B(n624), .Z(n625) );
  NOR2_X1 U715 ( .A1(n626), .A2(n625), .ZN(n928) );
  XOR2_X1 U716 ( .A(G2096), .B(n928), .Z(n627) );
  NOR2_X1 U717 ( .A1(G2100), .A2(n627), .ZN(n628) );
  XOR2_X1 U718 ( .A(KEYINPUT80), .B(n628), .Z(G156) );
  NAND2_X1 U719 ( .A1(G55), .A2(n656), .ZN(n629) );
  XNOR2_X1 U720 ( .A(n629), .B(KEYINPUT82), .ZN(n631) );
  NAND2_X1 U721 ( .A1(G93), .A2(n529), .ZN(n630) );
  NAND2_X1 U722 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U723 ( .A1(G80), .A2(n662), .ZN(n633) );
  NAND2_X1 U724 ( .A1(G67), .A2(n654), .ZN(n632) );
  NAND2_X1 U725 ( .A1(n633), .A2(n632), .ZN(n634) );
  OR2_X1 U726 ( .A1(n635), .A2(n634), .ZN(n674) );
  NAND2_X1 U727 ( .A1(n988), .A2(G559), .ZN(n636) );
  XOR2_X1 U728 ( .A(KEYINPUT81), .B(n636), .Z(n672) );
  XNOR2_X1 U729 ( .A(n993), .B(n672), .ZN(n637) );
  NOR2_X1 U730 ( .A1(G860), .A2(n637), .ZN(n638) );
  XOR2_X1 U731 ( .A(n674), .B(n638), .Z(G145) );
  NAND2_X1 U732 ( .A1(n656), .A2(G48), .ZN(n640) );
  NAND2_X1 U733 ( .A1(G86), .A2(n529), .ZN(n639) );
  NAND2_X1 U734 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U735 ( .A1(n662), .A2(G73), .ZN(n641) );
  XOR2_X1 U736 ( .A(KEYINPUT2), .B(n641), .Z(n642) );
  NOR2_X1 U737 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U738 ( .A1(n654), .A2(G61), .ZN(n644) );
  NAND2_X1 U739 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U740 ( .A1(n646), .A2(G87), .ZN(n651) );
  NAND2_X1 U741 ( .A1(G49), .A2(n656), .ZN(n648) );
  NAND2_X1 U742 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U743 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U744 ( .A1(n654), .A2(n649), .ZN(n650) );
  NAND2_X1 U745 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U746 ( .A(KEYINPUT83), .B(n652), .Z(G288) );
  NAND2_X1 U747 ( .A1(n529), .A2(G88), .ZN(n653) );
  XOR2_X1 U748 ( .A(KEYINPUT86), .B(n653), .Z(n661) );
  NAND2_X1 U749 ( .A1(n654), .A2(G62), .ZN(n655) );
  XNOR2_X1 U750 ( .A(n655), .B(KEYINPUT84), .ZN(n658) );
  NAND2_X1 U751 ( .A1(G50), .A2(n656), .ZN(n657) );
  NAND2_X1 U752 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U753 ( .A(KEYINPUT85), .B(n659), .Z(n660) );
  NOR2_X1 U754 ( .A1(n661), .A2(n660), .ZN(n664) );
  NAND2_X1 U755 ( .A1(n662), .A2(G75), .ZN(n663) );
  NAND2_X1 U756 ( .A1(n664), .A2(n663), .ZN(G303) );
  INV_X1 U757 ( .A(G303), .ZN(G166) );
  XOR2_X1 U758 ( .A(n674), .B(G305), .Z(n665) );
  XNOR2_X1 U759 ( .A(n665), .B(G288), .ZN(n666) );
  XNOR2_X1 U760 ( .A(KEYINPUT87), .B(n666), .ZN(n668) );
  XNOR2_X1 U761 ( .A(G290), .B(KEYINPUT19), .ZN(n667) );
  XNOR2_X1 U762 ( .A(n668), .B(n667), .ZN(n671) );
  XOR2_X1 U763 ( .A(n993), .B(G299), .Z(n669) );
  XOR2_X1 U764 ( .A(n669), .B(G166), .Z(n670) );
  XNOR2_X1 U765 ( .A(n671), .B(n670), .ZN(n913) );
  XNOR2_X1 U766 ( .A(n672), .B(n913), .ZN(n673) );
  NAND2_X1 U767 ( .A1(n673), .A2(G868), .ZN(n677) );
  NAND2_X1 U768 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U769 ( .A1(n677), .A2(n676), .ZN(G295) );
  NAND2_X1 U770 ( .A1(G2084), .A2(G2078), .ZN(n678) );
  XOR2_X1 U771 ( .A(KEYINPUT20), .B(n678), .Z(n679) );
  NAND2_X1 U772 ( .A1(n679), .A2(G2090), .ZN(n680) );
  XNOR2_X1 U773 ( .A(n680), .B(KEYINPUT88), .ZN(n681) );
  XNOR2_X1 U774 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U775 ( .A1(G2072), .A2(n682), .ZN(G158) );
  XNOR2_X1 U776 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U777 ( .A1(G220), .A2(G219), .ZN(n683) );
  XOR2_X1 U778 ( .A(KEYINPUT22), .B(n683), .Z(n684) );
  NOR2_X1 U779 ( .A1(G218), .A2(n684), .ZN(n685) );
  NAND2_X1 U780 ( .A1(G96), .A2(n685), .ZN(n848) );
  NAND2_X1 U781 ( .A1(G2106), .A2(n848), .ZN(n686) );
  XNOR2_X1 U782 ( .A(n686), .B(KEYINPUT89), .ZN(n690) );
  NOR2_X1 U783 ( .A1(G236), .A2(G238), .ZN(n687) );
  NAND2_X1 U784 ( .A1(G69), .A2(n687), .ZN(n688) );
  OR2_X1 U785 ( .A1(G237), .A2(n688), .ZN(n849) );
  AND2_X1 U786 ( .A1(G567), .A2(n849), .ZN(n689) );
  NOR2_X1 U787 ( .A1(n690), .A2(n689), .ZN(G319) );
  NAND2_X1 U788 ( .A1(G483), .A2(G661), .ZN(n692) );
  INV_X1 U789 ( .A(G319), .ZN(n691) );
  NOR2_X1 U790 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U791 ( .A(n693), .B(KEYINPUT90), .ZN(n847) );
  NAND2_X1 U792 ( .A1(G36), .A2(n847), .ZN(G176) );
  INV_X1 U793 ( .A(G40), .ZN(n694) );
  OR2_X1 U794 ( .A1(n695), .A2(n694), .ZN(n696) );
  INV_X1 U795 ( .A(n807), .ZN(n704) );
  INV_X1 U796 ( .A(G1996), .ZN(n862) );
  INV_X1 U797 ( .A(KEYINPUT26), .ZN(n698) );
  XNOR2_X1 U798 ( .A(n699), .B(n698), .ZN(n701) );
  NAND2_X1 U799 ( .A1(n745), .A2(G1341), .ZN(n700) );
  NAND2_X1 U800 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U801 ( .A1(n702), .A2(n993), .ZN(n710) );
  AND2_X1 U802 ( .A1(n710), .A2(n988), .ZN(n703) );
  XNOR2_X1 U803 ( .A(n703), .B(KEYINPUT97), .ZN(n708) );
  NOR2_X1 U804 ( .A1(n704), .A2(n806), .ZN(n724) );
  NOR2_X1 U805 ( .A1(n724), .A2(G1348), .ZN(n706) );
  NOR2_X1 U806 ( .A1(G2067), .A2(n745), .ZN(n705) );
  NOR2_X1 U807 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U808 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U809 ( .A(n709), .B(KEYINPUT98), .ZN(n712) );
  OR2_X1 U810 ( .A1(n988), .A2(n710), .ZN(n711) );
  NAND2_X1 U811 ( .A1(n712), .A2(n711), .ZN(n717) );
  NAND2_X1 U812 ( .A1(n724), .A2(G2072), .ZN(n713) );
  XNOR2_X1 U813 ( .A(n713), .B(KEYINPUT27), .ZN(n715) );
  INV_X1 U814 ( .A(G1956), .ZN(n859) );
  NOR2_X1 U815 ( .A1(n859), .A2(n724), .ZN(n714) );
  NOR2_X1 U816 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U817 ( .A1(n976), .A2(n718), .ZN(n716) );
  NAND2_X1 U818 ( .A1(n717), .A2(n716), .ZN(n721) );
  NOR2_X1 U819 ( .A1(n976), .A2(n718), .ZN(n719) );
  XOR2_X1 U820 ( .A(n719), .B(KEYINPUT28), .Z(n720) );
  NAND2_X1 U821 ( .A1(n721), .A2(n720), .ZN(n723) );
  XNOR2_X1 U822 ( .A(n723), .B(n722), .ZN(n727) );
  NAND2_X1 U823 ( .A1(G1961), .A2(n745), .ZN(n726) );
  XOR2_X1 U824 ( .A(G2078), .B(KEYINPUT25), .Z(n956) );
  NAND2_X1 U825 ( .A1(n724), .A2(n956), .ZN(n725) );
  NAND2_X1 U826 ( .A1(n726), .A2(n725), .ZN(n736) );
  NAND2_X1 U827 ( .A1(n727), .A2(n518), .ZN(n743) );
  NAND2_X1 U828 ( .A1(G8), .A2(n745), .ZN(n787) );
  NOR2_X1 U829 ( .A1(G1966), .A2(n787), .ZN(n729) );
  INV_X1 U830 ( .A(G8), .ZN(n730) );
  NOR2_X1 U831 ( .A1(G2084), .A2(n745), .ZN(n755) );
  NOR2_X1 U832 ( .A1(n730), .A2(n755), .ZN(n731) );
  XNOR2_X1 U833 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U834 ( .A1(G168), .A2(n734), .ZN(n735) );
  XNOR2_X1 U835 ( .A(n735), .B(KEYINPUT99), .ZN(n739) );
  NAND2_X1 U836 ( .A1(G301), .A2(n736), .ZN(n737) );
  XNOR2_X1 U837 ( .A(KEYINPUT100), .B(n737), .ZN(n738) );
  NAND2_X1 U838 ( .A1(n739), .A2(n738), .ZN(n741) );
  NAND2_X1 U839 ( .A1(n758), .A2(G286), .ZN(n750) );
  NOR2_X1 U840 ( .A1(G1971), .A2(n787), .ZN(n744) );
  XOR2_X1 U841 ( .A(KEYINPUT103), .B(n744), .Z(n747) );
  NOR2_X1 U842 ( .A1(G2090), .A2(n745), .ZN(n746) );
  NOR2_X1 U843 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U844 ( .A1(n748), .A2(G303), .ZN(n749) );
  NAND2_X1 U845 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U846 ( .A(n751), .B(KEYINPUT104), .ZN(n752) );
  NAND2_X1 U847 ( .A1(n752), .A2(G8), .ZN(n754) );
  NAND2_X1 U848 ( .A1(G8), .A2(n755), .ZN(n756) );
  NAND2_X1 U849 ( .A1(n757), .A2(n756), .ZN(n760) );
  XOR2_X1 U850 ( .A(n758), .B(KEYINPUT102), .Z(n759) );
  NOR2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X2 U852 ( .A1(n762), .A2(n761), .ZN(n778) );
  NOR2_X1 U853 ( .A1(G1971), .A2(G303), .ZN(n763) );
  XNOR2_X1 U854 ( .A(n763), .B(KEYINPUT105), .ZN(n765) );
  NOR2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n978) );
  INV_X1 U856 ( .A(n787), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n978), .A2(n771), .ZN(n764) );
  NAND2_X1 U858 ( .A1(n764), .A2(KEYINPUT33), .ZN(n769) );
  AND2_X1 U859 ( .A1(n765), .A2(n769), .ZN(n767) );
  INV_X1 U860 ( .A(n769), .ZN(n774) );
  INV_X1 U861 ( .A(KEYINPUT33), .ZN(n770) );
  NAND2_X1 U862 ( .A1(G1976), .A2(G288), .ZN(n981) );
  AND2_X1 U863 ( .A1(n770), .A2(n981), .ZN(n772) );
  AND2_X1 U864 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U865 ( .A(n776), .B(KEYINPUT106), .ZN(n777) );
  XOR2_X1 U866 ( .A(G1981), .B(G305), .Z(n973) );
  NAND2_X1 U867 ( .A1(n777), .A2(n973), .ZN(n784) );
  INV_X1 U868 ( .A(n778), .ZN(n781) );
  NOR2_X1 U869 ( .A1(G2090), .A2(G303), .ZN(n779) );
  NAND2_X1 U870 ( .A1(G8), .A2(n779), .ZN(n780) );
  NAND2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n782), .A2(n787), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n832) );
  NOR2_X1 U874 ( .A1(G1981), .A2(G305), .ZN(n785) );
  XNOR2_X1 U875 ( .A(n785), .B(KEYINPUT24), .ZN(n786) );
  XNOR2_X1 U876 ( .A(n786), .B(KEYINPUT95), .ZN(n788) );
  NOR2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n830) );
  NAND2_X1 U878 ( .A1(G141), .A2(n895), .ZN(n790) );
  NAND2_X1 U879 ( .A1(G117), .A2(n900), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n894), .A2(G105), .ZN(n791) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(n791), .Z(n792) );
  NOR2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n898), .A2(G129), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n891) );
  NOR2_X1 U886 ( .A1(G1996), .A2(n891), .ZN(n938) );
  NAND2_X1 U887 ( .A1(G131), .A2(n895), .ZN(n797) );
  NAND2_X1 U888 ( .A1(G119), .A2(n898), .ZN(n796) );
  NAND2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n801) );
  NAND2_X1 U890 ( .A1(G95), .A2(n894), .ZN(n799) );
  NAND2_X1 U891 ( .A1(G107), .A2(n900), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U894 ( .A(n802), .B(KEYINPUT93), .ZN(n906) );
  NAND2_X1 U895 ( .A1(G1991), .A2(n906), .ZN(n803) );
  XOR2_X1 U896 ( .A(KEYINPUT94), .B(n803), .Z(n805) );
  AND2_X1 U897 ( .A1(G1996), .A2(n891), .ZN(n804) );
  NOR2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n924) );
  INV_X1 U899 ( .A(n924), .ZN(n808) );
  NOR2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n833) );
  NAND2_X1 U901 ( .A1(n808), .A2(n833), .ZN(n834) );
  INV_X1 U902 ( .A(n834), .ZN(n811) );
  NOR2_X1 U903 ( .A1(G1991), .A2(n906), .ZN(n929) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U905 ( .A1(n929), .A2(n809), .ZN(n810) );
  NOR2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U907 ( .A1(n938), .A2(n812), .ZN(n813) );
  XNOR2_X1 U908 ( .A(n813), .B(KEYINPUT39), .ZN(n825) );
  NAND2_X1 U909 ( .A1(G104), .A2(n894), .ZN(n815) );
  NAND2_X1 U910 ( .A1(G140), .A2(n895), .ZN(n814) );
  NAND2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U912 ( .A(KEYINPUT34), .B(n816), .ZN(n822) );
  NAND2_X1 U913 ( .A1(G116), .A2(n900), .ZN(n818) );
  NAND2_X1 U914 ( .A1(G128), .A2(n898), .ZN(n817) );
  NAND2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U916 ( .A(KEYINPUT35), .B(n819), .ZN(n820) );
  XNOR2_X1 U917 ( .A(KEYINPUT91), .B(n820), .ZN(n821) );
  NOR2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U919 ( .A(KEYINPUT36), .B(n823), .ZN(n880) );
  XNOR2_X1 U920 ( .A(KEYINPUT37), .B(G2067), .ZN(n826) );
  NOR2_X1 U921 ( .A1(n880), .A2(n826), .ZN(n824) );
  XNOR2_X1 U922 ( .A(n824), .B(KEYINPUT92), .ZN(n927) );
  NAND2_X1 U923 ( .A1(n833), .A2(n927), .ZN(n835) );
  NAND2_X1 U924 ( .A1(n825), .A2(n835), .ZN(n827) );
  NAND2_X1 U925 ( .A1(n826), .A2(n880), .ZN(n944) );
  NAND2_X1 U926 ( .A1(n827), .A2(n944), .ZN(n828) );
  NAND2_X1 U927 ( .A1(n828), .A2(n833), .ZN(n839) );
  INV_X1 U928 ( .A(n839), .ZN(n829) );
  OR2_X1 U929 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U930 ( .A1(n832), .A2(n831), .ZN(n841) );
  XNOR2_X1 U931 ( .A(G1986), .B(G290), .ZN(n980) );
  AND2_X1 U932 ( .A1(n980), .A2(n833), .ZN(n837) );
  NAND2_X1 U933 ( .A1(n835), .A2(n834), .ZN(n836) );
  OR2_X1 U934 ( .A1(n837), .A2(n836), .ZN(n838) );
  AND2_X1 U935 ( .A1(n839), .A2(n838), .ZN(n840) );
  NOR2_X2 U936 ( .A1(n841), .A2(n840), .ZN(n843) );
  XOR2_X1 U937 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n842) );
  XNOR2_X1 U938 ( .A(n843), .B(n842), .ZN(G329) );
  NAND2_X1 U939 ( .A1(G2106), .A2(n844), .ZN(G217) );
  AND2_X1 U940 ( .A1(G15), .A2(G2), .ZN(n845) );
  NAND2_X1 U941 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U942 ( .A1(G3), .A2(G1), .ZN(n846) );
  NAND2_X1 U943 ( .A1(n847), .A2(n846), .ZN(G188) );
  NOR2_X1 U944 ( .A1(n849), .A2(n848), .ZN(G325) );
  XOR2_X1 U945 ( .A(KEYINPUT108), .B(G325), .Z(G261) );
  INV_X1 U947 ( .A(G96), .ZN(G221) );
  XOR2_X1 U948 ( .A(KEYINPUT42), .B(G2090), .Z(n851) );
  XNOR2_X1 U949 ( .A(G2078), .B(G2072), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U951 ( .A(n852), .B(G2100), .Z(n854) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2084), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U954 ( .A(G2096), .B(KEYINPUT43), .Z(n856) );
  XNOR2_X1 U955 ( .A(G2678), .B(KEYINPUT109), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U957 ( .A(n858), .B(n857), .Z(G227) );
  XNOR2_X1 U958 ( .A(G1986), .B(G2474), .ZN(n870) );
  XOR2_X1 U959 ( .A(G1976), .B(G1971), .Z(n861) );
  XOR2_X1 U960 ( .A(G1961), .B(n859), .Z(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n866) );
  XOR2_X1 U962 ( .A(G1981), .B(G1966), .Z(n864) );
  XOR2_X1 U963 ( .A(n862), .B(G1991), .Z(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U965 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U966 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(G229) );
  NAND2_X1 U969 ( .A1(G124), .A2(n898), .ZN(n871) );
  XNOR2_X1 U970 ( .A(n871), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G112), .A2(n900), .ZN(n872) );
  XOR2_X1 U972 ( .A(KEYINPUT111), .B(n872), .Z(n873) );
  NAND2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n878) );
  NAND2_X1 U974 ( .A1(G100), .A2(n894), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G136), .A2(n895), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U977 ( .A1(n878), .A2(n877), .ZN(G162) );
  XOR2_X1 U978 ( .A(G160), .B(n928), .Z(n879) );
  XNOR2_X1 U979 ( .A(n880), .B(n879), .ZN(n890) );
  NAND2_X1 U980 ( .A1(G118), .A2(n900), .ZN(n882) );
  NAND2_X1 U981 ( .A1(G130), .A2(n898), .ZN(n881) );
  NAND2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n888) );
  NAND2_X1 U983 ( .A1(G106), .A2(n894), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G142), .A2(n895), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U986 ( .A(KEYINPUT45), .B(n885), .Z(n886) );
  XNOR2_X1 U987 ( .A(KEYINPUT112), .B(n886), .ZN(n887) );
  NOR2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U989 ( .A(n890), .B(n889), .Z(n893) );
  XOR2_X1 U990 ( .A(n891), .B(G162), .Z(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n911) );
  XNOR2_X1 U992 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n908) );
  NAND2_X1 U993 ( .A1(G103), .A2(n894), .ZN(n897) );
  NAND2_X1 U994 ( .A1(G139), .A2(n895), .ZN(n896) );
  NAND2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n905) );
  NAND2_X1 U996 ( .A1(n898), .A2(G127), .ZN(n899) );
  XOR2_X1 U997 ( .A(KEYINPUT113), .B(n899), .Z(n902) );
  NAND2_X1 U998 ( .A1(n900), .A2(G115), .ZN(n901) );
  NAND2_X1 U999 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1000 ( .A(KEYINPUT47), .B(n903), .Z(n904) );
  NOR2_X1 U1001 ( .A1(n905), .A2(n904), .ZN(n933) );
  XNOR2_X1 U1002 ( .A(n906), .B(n933), .ZN(n907) );
  XNOR2_X1 U1003 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1004 ( .A(G164), .B(n909), .Z(n910) );
  XNOR2_X1 U1005 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n912), .ZN(G395) );
  XOR2_X1 U1007 ( .A(n988), .B(G286), .Z(n914) );
  XNOR2_X1 U1008 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1009 ( .A(n915), .B(G301), .Z(n916) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n916), .ZN(G397) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n917) );
  XOR2_X1 U1012 ( .A(KEYINPUT49), .B(n917), .Z(n918) );
  XNOR2_X1 U1013 ( .A(KEYINPUT114), .B(n918), .ZN(n923) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n919) );
  XOR2_X1 U1015 ( .A(KEYINPUT115), .B(n919), .Z(n920) );
  NAND2_X1 U1016 ( .A1(G319), .A2(n920), .ZN(n921) );
  NOR2_X1 U1017 ( .A1(G401), .A2(n921), .ZN(n922) );
  NAND2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1021 ( .A(G160), .B(G2084), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n931) );
  NOR2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1026 ( .A(KEYINPUT116), .B(n932), .ZN(n943) );
  XOR2_X1 U1027 ( .A(G2072), .B(n933), .Z(n935) );
  XOR2_X1 U1028 ( .A(G164), .B(G2078), .Z(n934) );
  NOR2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1030 ( .A(KEYINPUT50), .B(n936), .ZN(n941) );
  XOR2_X1 U1031 ( .A(G2090), .B(G162), .Z(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1033 ( .A(KEYINPUT51), .B(n939), .Z(n940) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n945) );
  NAND2_X1 U1036 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n946), .ZN(n947) );
  NAND2_X1 U1038 ( .A1(n947), .A2(G29), .ZN(n1028) );
  XNOR2_X1 U1039 ( .A(G1991), .B(G25), .ZN(n949) );
  XNOR2_X1 U1040 ( .A(G33), .B(G2072), .ZN(n948) );
  NOR2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n955) );
  XOR2_X1 U1042 ( .A(G2067), .B(G26), .Z(n950) );
  NAND2_X1 U1043 ( .A1(n950), .A2(G28), .ZN(n953) );
  XNOR2_X1 U1044 ( .A(KEYINPUT118), .B(G1996), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(G32), .B(n951), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n958) );
  XNOR2_X1 U1048 ( .A(G27), .B(n956), .ZN(n957) );
  NOR2_X1 U1049 ( .A1(n958), .A2(n957), .ZN(n961) );
  XNOR2_X1 U1050 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(n959), .B(KEYINPUT53), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(n961), .B(n960), .ZN(n968) );
  XOR2_X1 U1053 ( .A(KEYINPUT121), .B(G34), .Z(n963) );
  XNOR2_X1 U1054 ( .A(G2084), .B(KEYINPUT54), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(n963), .B(n962), .ZN(n966) );
  XOR2_X1 U1056 ( .A(KEYINPUT117), .B(G2090), .Z(n964) );
  XNOR2_X1 U1057 ( .A(G35), .B(n964), .ZN(n965) );
  NOR2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1060 ( .A(KEYINPUT122), .B(n969), .Z(n970) );
  NOR2_X1 U1061 ( .A1(G29), .A2(n970), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(KEYINPUT55), .B(n971), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(n972), .A2(G11), .ZN(n1026) );
  INV_X1 U1064 ( .A(G16), .ZN(n1022) );
  XOR2_X1 U1065 ( .A(n1022), .B(KEYINPUT56), .Z(n999) );
  XNOR2_X1 U1066 ( .A(G1966), .B(G168), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n975), .B(KEYINPUT57), .ZN(n997) );
  XOR2_X1 U1069 ( .A(G1956), .B(n976), .Z(n977) );
  XNOR2_X1 U1070 ( .A(n977), .B(KEYINPUT123), .ZN(n986) );
  XNOR2_X1 U1071 ( .A(KEYINPUT124), .B(n978), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n984) );
  XOR2_X1 U1074 ( .A(G1971), .B(G166), .Z(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(KEYINPUT125), .B(n987), .ZN(n992) );
  XOR2_X1 U1078 ( .A(G171), .B(G1961), .Z(n990) );
  XOR2_X1 U1079 ( .A(n988), .B(G1348), .Z(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(G1341), .B(n993), .ZN(n994) );
  NOR2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1024) );
  XNOR2_X1 U1086 ( .A(G1966), .B(G21), .ZN(n1001) );
  XNOR2_X1 U1087 ( .A(G5), .B(G1961), .ZN(n1000) );
  NOR2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1012) );
  XOR2_X1 U1089 ( .A(KEYINPUT126), .B(G4), .Z(n1003) );
  XNOR2_X1 U1090 ( .A(G1348), .B(KEYINPUT59), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(n1003), .B(n1002), .ZN(n1009) );
  XOR2_X1 U1092 ( .A(G20), .B(G1956), .Z(n1007) );
  XNOR2_X1 U1093 ( .A(G1341), .B(G19), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(G1981), .B(G6), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(n1010), .B(KEYINPUT60), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1019) );
  XNOR2_X1 U1100 ( .A(G1971), .B(G22), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(G23), .B(G1976), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(G1986), .B(G24), .Z(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(KEYINPUT58), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1020), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1112 ( .A(n1029), .B(KEYINPUT62), .ZN(n1030) );
  XOR2_X1 U1113 ( .A(KEYINPUT127), .B(n1030), .Z(G150) );
  INV_X1 U1114 ( .A(G150), .ZN(G311) );
endmodule

