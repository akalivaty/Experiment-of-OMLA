

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U320 ( .A(n412), .B(KEYINPUT48), .ZN(n550) );
  NOR2_X2 U321 ( .A1(n405), .A2(n578), .ZN(n407) );
  XNOR2_X1 U322 ( .A(n445), .B(KEYINPUT122), .ZN(n564) );
  XNOR2_X1 U323 ( .A(n575), .B(KEYINPUT41), .ZN(n552) );
  XNOR2_X2 U324 ( .A(n342), .B(n341), .ZN(n575) );
  XNOR2_X1 U325 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U326 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U327 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U328 ( .A(n401), .B(n400), .Z(n565) );
  XOR2_X1 U329 ( .A(n366), .B(n335), .Z(n288) );
  XNOR2_X1 U330 ( .A(n379), .B(KEYINPUT66), .ZN(n380) );
  XOR2_X1 U331 ( .A(G155GAT), .B(G22GAT), .Z(n345) );
  XNOR2_X1 U332 ( .A(n408), .B(KEYINPUT47), .ZN(n409) );
  XNOR2_X1 U333 ( .A(n393), .B(G113GAT), .ZN(n394) );
  INV_X1 U334 ( .A(n345), .ZN(n302) );
  NOR2_X1 U335 ( .A1(n464), .A2(n568), .ZN(n430) );
  XNOR2_X1 U336 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U337 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U338 ( .A(n473), .B(KEYINPUT99), .ZN(n474) );
  XNOR2_X1 U339 ( .A(n355), .B(n354), .ZN(n357) );
  XNOR2_X1 U340 ( .A(n475), .B(n474), .ZN(n519) );
  XNOR2_X1 U341 ( .A(n476), .B(KEYINPUT38), .ZN(n477) );
  NOR2_X1 U342 ( .A1(n564), .A2(n561), .ZN(n482) );
  XOR2_X1 U343 ( .A(KEYINPUT101), .B(n477), .Z(n504) );
  XNOR2_X1 U344 ( .A(n450), .B(KEYINPUT124), .ZN(n451) );
  XNOR2_X1 U345 ( .A(n452), .B(n451), .ZN(G1350GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT84), .B(KEYINPUT22), .Z(n290) );
  XNOR2_X1 U347 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n289) );
  XNOR2_X1 U348 ( .A(n290), .B(n289), .ZN(n307) );
  XOR2_X1 U349 ( .A(KEYINPUT83), .B(KEYINPUT86), .Z(n292) );
  NAND2_X1 U350 ( .A1(G228GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U351 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U352 ( .A(n293), .B(KEYINPUT24), .Z(n299) );
  XOR2_X1 U353 ( .A(G197GAT), .B(KEYINPUT21), .Z(n295) );
  XNOR2_X1 U354 ( .A(G218GAT), .B(G211GAT), .ZN(n294) );
  XNOR2_X1 U355 ( .A(n295), .B(n294), .ZN(n423) );
  XOR2_X1 U356 ( .A(KEYINPUT77), .B(G78GAT), .Z(n297) );
  XNOR2_X1 U357 ( .A(G148GAT), .B(G106GAT), .ZN(n296) );
  XNOR2_X1 U358 ( .A(n297), .B(n296), .ZN(n338) );
  XNOR2_X1 U359 ( .A(n423), .B(n338), .ZN(n298) );
  XNOR2_X1 U360 ( .A(n299), .B(n298), .ZN(n305) );
  XOR2_X1 U361 ( .A(KEYINPUT85), .B(KEYINPUT3), .Z(n301) );
  XNOR2_X1 U362 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n300) );
  XNOR2_X1 U363 ( .A(n301), .B(n300), .ZN(n319) );
  XOR2_X1 U364 ( .A(G162GAT), .B(G50GAT), .Z(n363) );
  XNOR2_X1 U365 ( .A(n319), .B(n363), .ZN(n303) );
  XNOR2_X1 U366 ( .A(n307), .B(n306), .ZN(n464) );
  XOR2_X1 U367 ( .A(KEYINPUT1), .B(KEYINPUT88), .Z(n309) );
  XNOR2_X1 U368 ( .A(KEYINPUT4), .B(KEYINPUT89), .ZN(n308) );
  XNOR2_X1 U369 ( .A(n309), .B(n308), .ZN(n326) );
  XOR2_X1 U370 ( .A(G148GAT), .B(G1GAT), .Z(n311) );
  XNOR2_X1 U371 ( .A(G85GAT), .B(G162GAT), .ZN(n310) );
  XNOR2_X1 U372 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U373 ( .A(KEYINPUT87), .B(KEYINPUT5), .Z(n313) );
  XNOR2_X1 U374 ( .A(G57GAT), .B(G155GAT), .ZN(n312) );
  XNOR2_X1 U375 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U376 ( .A(n315), .B(n314), .Z(n324) );
  XOR2_X1 U377 ( .A(G113GAT), .B(G134GAT), .Z(n317) );
  XNOR2_X1 U378 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U380 ( .A(G120GAT), .B(n318), .Z(n443) );
  XOR2_X1 U381 ( .A(n319), .B(KEYINPUT6), .Z(n321) );
  NAND2_X1 U382 ( .A1(G225GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n443), .B(n322), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U386 ( .A(n326), .B(n325), .ZN(n478) );
  XNOR2_X1 U387 ( .A(G29GAT), .B(n478), .ZN(n548) );
  XOR2_X1 U388 ( .A(KEYINPUT75), .B(KEYINPUT13), .Z(n328) );
  XNOR2_X1 U389 ( .A(KEYINPUT74), .B(G71GAT), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U391 ( .A(G57GAT), .B(n329), .ZN(n356) );
  XOR2_X1 U392 ( .A(G204GAT), .B(KEYINPUT78), .Z(n331) );
  XNOR2_X1 U393 ( .A(G92GAT), .B(G176GAT), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U395 ( .A(G64GAT), .B(n332), .Z(n414) );
  XOR2_X1 U396 ( .A(n356), .B(n414), .Z(n342) );
  XOR2_X1 U397 ( .A(G85GAT), .B(G99GAT), .Z(n366) );
  XOR2_X1 U398 ( .A(KEYINPUT76), .B(KEYINPUT31), .Z(n334) );
  XNOR2_X1 U399 ( .A(G120GAT), .B(KEYINPUT79), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n334), .B(n333), .ZN(n335) );
  NAND2_X1 U401 ( .A1(G230GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U402 ( .A(n288), .B(n336), .ZN(n337) );
  XOR2_X1 U403 ( .A(n337), .B(KEYINPUT32), .Z(n340) );
  XNOR2_X1 U404 ( .A(n338), .B(KEYINPUT33), .ZN(n339) );
  XNOR2_X1 U405 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U406 ( .A(KEYINPUT81), .B(KEYINPUT14), .Z(n344) );
  XNOR2_X1 U407 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n349) );
  XOR2_X1 U409 ( .A(G64GAT), .B(G8GAT), .Z(n347) );
  XOR2_X1 U410 ( .A(G1GAT), .B(G15GAT), .Z(n392) );
  XNOR2_X1 U411 ( .A(n392), .B(n345), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U413 ( .A(n349), .B(n348), .Z(n355) );
  XOR2_X1 U414 ( .A(G78GAT), .B(G183GAT), .Z(n351) );
  XNOR2_X1 U415 ( .A(G127GAT), .B(G211GAT), .ZN(n350) );
  XNOR2_X1 U416 ( .A(n351), .B(n350), .ZN(n353) );
  NAND2_X1 U417 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XOR2_X1 U418 ( .A(n357), .B(n356), .Z(n558) );
  INV_X1 U419 ( .A(n558), .ZN(n578) );
  XOR2_X1 U420 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n359) );
  XNOR2_X1 U421 ( .A(KEYINPUT64), .B(G106GAT), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n377) );
  XOR2_X1 U423 ( .A(KEYINPUT67), .B(G92GAT), .Z(n361) );
  XNOR2_X1 U424 ( .A(KEYINPUT11), .B(KEYINPUT80), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n362), .B(G218GAT), .ZN(n365) );
  XOR2_X1 U427 ( .A(G134GAT), .B(n363), .Z(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n370) );
  XOR2_X1 U429 ( .A(n366), .B(KEYINPUT10), .Z(n368) );
  NAND2_X1 U430 ( .A1(G232GAT), .A2(G233GAT), .ZN(n367) );
  XOR2_X1 U431 ( .A(n368), .B(n367), .Z(n369) );
  XNOR2_X1 U432 ( .A(n370), .B(n369), .ZN(n375) );
  XOR2_X1 U433 ( .A(KEYINPUT8), .B(KEYINPUT72), .Z(n372) );
  XNOR2_X1 U434 ( .A(G43GAT), .B(G29GAT), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U436 ( .A(KEYINPUT7), .B(n373), .Z(n401) );
  XOR2_X1 U437 ( .A(G190GAT), .B(G36GAT), .Z(n418) );
  XNOR2_X1 U438 ( .A(n401), .B(n418), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U440 ( .A(n377), .B(n376), .Z(n406) );
  XNOR2_X1 U441 ( .A(n406), .B(KEYINPUT97), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n378), .B(KEYINPUT36), .ZN(n471) );
  AND2_X1 U443 ( .A1(n578), .A2(n471), .ZN(n381) );
  INV_X1 U444 ( .A(KEYINPUT45), .ZN(n379) );
  NOR2_X1 U445 ( .A1(n575), .A2(n382), .ZN(n383) );
  XNOR2_X1 U446 ( .A(KEYINPUT112), .B(n383), .ZN(n402) );
  XOR2_X1 U447 ( .A(KEYINPUT30), .B(KEYINPUT73), .Z(n385) );
  XNOR2_X1 U448 ( .A(G141GAT), .B(G22GAT), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n399) );
  XOR2_X1 U450 ( .A(KEYINPUT29), .B(G197GAT), .Z(n387) );
  XNOR2_X1 U451 ( .A(G36GAT), .B(G50GAT), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U453 ( .A(KEYINPUT68), .B(KEYINPUT71), .Z(n389) );
  XNOR2_X1 U454 ( .A(KEYINPUT70), .B(KEYINPUT69), .ZN(n388) );
  XNOR2_X1 U455 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U456 ( .A(n391), .B(n390), .Z(n397) );
  XOR2_X1 U457 ( .A(G8GAT), .B(G169GAT), .Z(n413) );
  XOR2_X1 U458 ( .A(n413), .B(n392), .Z(n395) );
  NAND2_X1 U459 ( .A1(G229GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U460 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U461 ( .A(n399), .B(n398), .Z(n400) );
  NAND2_X1 U462 ( .A1(n402), .A2(n565), .ZN(n411) );
  NOR2_X1 U463 ( .A1(n565), .A2(n552), .ZN(n404) );
  XNOR2_X1 U464 ( .A(KEYINPUT46), .B(KEYINPUT110), .ZN(n403) );
  XNOR2_X1 U465 ( .A(n404), .B(n403), .ZN(n405) );
  BUF_X1 U466 ( .A(n406), .Z(n561) );
  NAND2_X1 U467 ( .A1(n407), .A2(n561), .ZN(n408) );
  XNOR2_X1 U468 ( .A(n409), .B(KEYINPUT111), .ZN(n410) );
  NAND2_X1 U469 ( .A1(n411), .A2(n410), .ZN(n412) );
  XOR2_X1 U470 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n416) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U473 ( .A(n418), .B(n417), .Z(n420) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n425) );
  XOR2_X1 U476 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n422) );
  XNOR2_X1 U477 ( .A(G183GAT), .B(KEYINPUT17), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n437) );
  XNOR2_X1 U479 ( .A(n437), .B(n423), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n458) );
  INV_X1 U481 ( .A(n458), .ZN(n497) );
  NAND2_X1 U482 ( .A1(n550), .A2(n497), .ZN(n427) );
  XNOR2_X1 U483 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n426) );
  XOR2_X1 U484 ( .A(n427), .B(n426), .Z(n428) );
  NAND2_X1 U485 ( .A1(n548), .A2(n428), .ZN(n568) );
  XNOR2_X1 U486 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n444) );
  XOR2_X1 U488 ( .A(G169GAT), .B(G99GAT), .Z(n432) );
  XNOR2_X1 U489 ( .A(G43GAT), .B(G190GAT), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U491 ( .A(KEYINPUT20), .B(G176GAT), .Z(n434) );
  XNOR2_X1 U492 ( .A(G71GAT), .B(G15GAT), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n441) );
  XOR2_X1 U495 ( .A(n437), .B(KEYINPUT82), .Z(n439) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U497 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U499 ( .A(n443), .B(n442), .Z(n500) );
  NAND2_X1 U500 ( .A1(n444), .A2(n500), .ZN(n445) );
  XNOR2_X1 U501 ( .A(KEYINPUT104), .B(n552), .ZN(n535) );
  NOR2_X1 U502 ( .A1(n564), .A2(n535), .ZN(n449) );
  XOR2_X1 U503 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n447) );
  XNOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(G1349GAT) );
  NOR2_X1 U507 ( .A1(n558), .A2(n564), .ZN(n452) );
  INV_X1 U508 ( .A(G183GAT), .ZN(n450) );
  INV_X1 U509 ( .A(KEYINPUT27), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n453), .B(n458), .ZN(n465) );
  XNOR2_X1 U511 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n454), .B(KEYINPUT26), .ZN(n457) );
  INV_X1 U513 ( .A(n464), .ZN(n455) );
  NOR2_X1 U514 ( .A1(n500), .A2(n455), .ZN(n456) );
  XOR2_X1 U515 ( .A(n457), .B(n456), .Z(n567) );
  NAND2_X1 U516 ( .A1(n465), .A2(n567), .ZN(n547) );
  XNOR2_X1 U517 ( .A(n547), .B(KEYINPUT94), .ZN(n462) );
  INV_X1 U518 ( .A(n500), .ZN(n532) );
  NOR2_X1 U519 ( .A1(n458), .A2(n532), .ZN(n459) );
  NOR2_X1 U520 ( .A1(n464), .A2(n459), .ZN(n460) );
  XNOR2_X1 U521 ( .A(KEYINPUT25), .B(n460), .ZN(n461) );
  NAND2_X1 U522 ( .A1(n462), .A2(n461), .ZN(n463) );
  NAND2_X1 U523 ( .A1(n463), .A2(n548), .ZN(n468) );
  XOR2_X1 U524 ( .A(n464), .B(KEYINPUT28), .Z(n527) );
  NAND2_X1 U525 ( .A1(n465), .A2(n527), .ZN(n466) );
  NOR2_X1 U526 ( .A1(n548), .A2(n466), .ZN(n530) );
  NAND2_X1 U527 ( .A1(n530), .A2(n532), .ZN(n467) );
  NAND2_X1 U528 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U529 ( .A(KEYINPUT95), .B(n469), .ZN(n487) );
  NOR2_X1 U530 ( .A1(n487), .A2(n578), .ZN(n470) );
  XNOR2_X1 U531 ( .A(KEYINPUT98), .B(n470), .ZN(n472) );
  NAND2_X1 U532 ( .A1(n472), .A2(n471), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT100), .B(KEYINPUT37), .Z(n473) );
  NOR2_X1 U534 ( .A1(n565), .A2(n575), .ZN(n488) );
  NAND2_X1 U535 ( .A1(n519), .A2(n488), .ZN(n476) );
  INV_X1 U536 ( .A(n504), .ZN(n501) );
  NOR2_X1 U537 ( .A1(G29GAT), .A2(n501), .ZN(n480) );
  NOR2_X1 U538 ( .A1(n504), .A2(n478), .ZN(n479) );
  OR2_X1 U539 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(KEYINPUT39), .ZN(G1328GAT) );
  INV_X1 U541 ( .A(G190GAT), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n482), .B(KEYINPUT58), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(G1351GAT) );
  NAND2_X1 U544 ( .A1(n561), .A2(n578), .ZN(n485) );
  XNOR2_X1 U545 ( .A(KEYINPUT16), .B(n485), .ZN(n486) );
  NOR2_X1 U546 ( .A1(n487), .A2(n486), .ZN(n507) );
  NAND2_X1 U547 ( .A1(n488), .A2(n507), .ZN(n495) );
  NOR2_X1 U548 ( .A1(n548), .A2(n495), .ZN(n489) );
  XOR2_X1 U549 ( .A(KEYINPUT34), .B(n489), .Z(n490) );
  XNOR2_X1 U550 ( .A(G1GAT), .B(n490), .ZN(G1324GAT) );
  INV_X1 U551 ( .A(n497), .ZN(n523) );
  NOR2_X1 U552 ( .A1(n523), .A2(n495), .ZN(n491) );
  XOR2_X1 U553 ( .A(KEYINPUT96), .B(n491), .Z(n492) );
  XNOR2_X1 U554 ( .A(G8GAT), .B(n492), .ZN(G1325GAT) );
  NOR2_X1 U555 ( .A1(n532), .A2(n495), .ZN(n494) );
  XNOR2_X1 U556 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NOR2_X1 U558 ( .A1(n527), .A2(n495), .ZN(n496) );
  XOR2_X1 U559 ( .A(G22GAT), .B(n496), .Z(G1327GAT) );
  NAND2_X1 U560 ( .A1(n501), .A2(n497), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n498), .B(KEYINPUT102), .ZN(n499) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n499), .ZN(G1329GAT) );
  NAND2_X1 U563 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n502), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NOR2_X1 U566 ( .A1(n504), .A2(n527), .ZN(n506) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(KEYINPUT103), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(G1331GAT) );
  INV_X1 U569 ( .A(n565), .ZN(n570) );
  NOR2_X1 U570 ( .A1(n535), .A2(n570), .ZN(n520) );
  NAND2_X1 U571 ( .A1(n520), .A2(n507), .ZN(n514) );
  NOR2_X1 U572 ( .A1(n548), .A2(n514), .ZN(n508) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n508), .Z(n509) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(n509), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n523), .A2(n514), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(KEYINPUT105), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1333GAT) );
  NOR2_X1 U578 ( .A1(n532), .A2(n514), .ZN(n512) );
  XOR2_X1 U579 ( .A(KEYINPUT106), .B(n512), .Z(n513) );
  XNOR2_X1 U580 ( .A(G71GAT), .B(n513), .ZN(G1334GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n527), .ZN(n518) );
  XOR2_X1 U582 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n516) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT108), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n526) );
  NOR2_X1 U587 ( .A1(n548), .A2(n526), .ZN(n522) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(G1336GAT) );
  NOR2_X1 U590 ( .A1(n523), .A2(n526), .ZN(n524) );
  XOR2_X1 U591 ( .A(G92GAT), .B(n524), .Z(G1337GAT) );
  NOR2_X1 U592 ( .A1(n532), .A2(n526), .ZN(n525) );
  XOR2_X1 U593 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  NOR2_X1 U594 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U595 ( .A(KEYINPUT44), .B(n528), .Z(n529) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NAND2_X1 U597 ( .A1(n530), .A2(n550), .ZN(n531) );
  NOR2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U599 ( .A(KEYINPUT113), .B(n533), .ZN(n544) );
  INV_X1 U600 ( .A(n544), .ZN(n540) );
  NAND2_X1 U601 ( .A1(n570), .A2(n540), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n534), .B(G113GAT), .ZN(G1340GAT) );
  NOR2_X1 U603 ( .A1(n544), .A2(n535), .ZN(n539) );
  XOR2_X1 U604 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n537) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n536) );
  XNOR2_X1 U606 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n542) );
  NAND2_X1 U609 ( .A1(n540), .A2(n578), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U611 ( .A(G127GAT), .B(n543), .Z(G1342GAT) );
  NOR2_X1 U612 ( .A1(n561), .A2(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NOR2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n560) );
  NOR2_X1 U617 ( .A1(n565), .A2(n560), .ZN(n551) );
  XOR2_X1 U618 ( .A(G141GAT), .B(n551), .Z(G1344GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n560), .ZN(n557) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n554) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(KEYINPUT117), .B(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n558), .A2(n560), .ZN(n559) );
  XOR2_X1 U626 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1347GAT) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U631 ( .A(G169GAT), .B(n566), .Z(G1348GAT) );
  INV_X1 U632 ( .A(n567), .ZN(n569) );
  NOR2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n581) );
  AND2_X1 U634 ( .A1(n581), .A2(n570), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n572) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U640 ( .A1(n581), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U642 ( .A1(n578), .A2(n581), .ZN(n579) );
  XNOR2_X1 U643 ( .A(n579), .B(KEYINPUT126), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n580), .ZN(G1354GAT) );
  NAND2_X1 U645 ( .A1(n581), .A2(n471), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

