//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(new_n202), .A2(G50), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(new_n208), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G87), .A2(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G116), .ZN(new_n214));
  INV_X1    g0014(.A(G270), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI211_X1 g0022(.A(new_n216), .B(new_n222), .C1(G107), .C2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT65), .B(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n212), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT1), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n210), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(G13), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n212), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT64), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT0), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n229), .B(new_n235), .C1(new_n228), .C2(new_n227), .ZN(G361));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n219), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n207), .ZN(new_n254));
  OAI21_X1  g0054(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n255), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n208), .A2(new_n256), .A3(KEYINPUT68), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT68), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G20), .B2(G33), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G150), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n254), .B1(new_n260), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G50), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n269), .A2(new_n254), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT69), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT69), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(new_n269), .B2(new_n254), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n211), .A2(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n267), .B(new_n271), .C1(new_n278), .C2(new_n270), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G1), .A3(G13), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(new_n284), .A3(G274), .ZN(new_n285));
  INV_X1    g0085(.A(G226), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G222), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(G1698), .ZN(new_n293));
  XOR2_X1   g0093(.A(KEYINPUT67), .B(G223), .Z(new_n294));
  OAI221_X1 g0094(.A(new_n292), .B1(new_n220), .B2(new_n290), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n207), .B1(G33), .B2(G41), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n289), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n279), .B1(new_n297), .B2(G169), .ZN(new_n298));
  INV_X1    g0098(.A(G179), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(new_n297), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n279), .B(KEYINPUT9), .ZN(new_n301));
  INV_X1    g0101(.A(G200), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(G190), .B2(new_n297), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n301), .A2(new_n307), .A3(new_n304), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n300), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G33), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n310), .A2(new_n312), .A3(G232), .A4(G1698), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n310), .A2(new_n312), .A3(G226), .A4(new_n291), .ZN(new_n314));
  NAND2_X1  g0114(.A1(G33), .A2(G97), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n296), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n284), .A2(G238), .A3(new_n287), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n285), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(KEYINPUT72), .A3(KEYINPUT13), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT72), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n319), .B1(new_n296), .B2(new_n316), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT13), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n325), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n322), .A2(new_n326), .A3(G179), .A4(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT14), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n317), .A2(new_n320), .A3(new_n325), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n325), .B1(new_n317), .B2(new_n320), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n329), .B(G169), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT74), .ZN(new_n334));
  INV_X1    g0134(.A(G169), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n321), .A2(KEYINPUT13), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(new_n327), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n334), .B1(new_n337), .B2(new_n329), .ZN(new_n338));
  OAI21_X1  g0138(.A(G169), .B1(new_n330), .B2(new_n331), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(KEYINPUT74), .A3(KEYINPUT14), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n333), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n253), .A2(new_n207), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n261), .A2(new_n263), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G50), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n257), .A2(G77), .B1(G20), .B2(new_n225), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n342), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n346), .A2(KEYINPUT11), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n230), .A2(G1), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n348), .A2(KEYINPUT70), .A3(G20), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT70), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n268), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n352), .A2(G68), .A3(new_n342), .A4(new_n277), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n346), .A2(KEYINPUT11), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT12), .B1(new_n352), .B2(G68), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT12), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n348), .A2(new_n356), .A3(G20), .A4(new_n225), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n347), .A2(new_n353), .A3(new_n354), .A4(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n341), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n264), .A2(new_n259), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT15), .B(G87), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n364), .A2(new_n258), .B1(new_n208), .B2(new_n220), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n254), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AND4_X1   g0167(.A1(G77), .A2(new_n352), .A3(new_n342), .A4(new_n277), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n352), .A2(G77), .ZN(new_n369));
  OR3_X1    g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n285), .B1(new_n221), .B2(new_n288), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n290), .A2(G232), .A3(new_n291), .ZN(new_n372));
  INV_X1    g0172(.A(G107), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n372), .B1(new_n373), .B2(new_n290), .C1(new_n293), .C2(new_n224), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n371), .B1(new_n374), .B2(new_n296), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n370), .B1(G190), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n302), .B2(new_n375), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n299), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n370), .B(new_n378), .C1(G169), .C2(new_n375), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n309), .A2(new_n362), .A3(new_n377), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n343), .A2(G159), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n218), .A2(new_n225), .ZN(new_n382));
  OAI21_X1  g0182(.A(G20), .B1(new_n382), .B2(new_n201), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n290), .B2(G20), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n310), .A2(new_n312), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n388), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n387), .A2(new_n389), .A3(KEYINPUT75), .ZN(new_n390));
  OAI21_X1  g0190(.A(G68), .B1(new_n387), .B2(KEYINPUT75), .ZN(new_n391));
  OAI211_X1 g0191(.A(KEYINPUT16), .B(new_n385), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n225), .B1(new_n387), .B2(new_n389), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(new_n384), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(new_n254), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n259), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(new_n269), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n273), .A2(new_n275), .B1(new_n211), .B2(G20), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n399), .B1(new_n400), .B2(new_n259), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n284), .A2(G232), .A3(new_n287), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT76), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT76), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n284), .A2(new_n287), .A3(new_n405), .A4(G232), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n284), .A2(G274), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n404), .A2(new_n406), .B1(new_n407), .B2(new_n282), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n310), .A2(new_n312), .A3(G226), .A4(G1698), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n310), .A2(new_n312), .A3(G223), .A4(new_n291), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G87), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n296), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n335), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n404), .A2(new_n406), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n416), .A3(new_n285), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n415), .B1(new_n299), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n402), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n417), .A2(new_n302), .ZN(new_n422));
  INV_X1    g0222(.A(G190), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n408), .A2(new_n423), .A3(new_n413), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n396), .A2(new_n425), .A3(new_n401), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT17), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n421), .A2(KEYINPUT77), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT77), .B1(new_n421), .B2(new_n427), .ZN(new_n429));
  OAI21_X1  g0229(.A(G200), .B1(new_n330), .B2(new_n331), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT71), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(KEYINPUT71), .B(G200), .C1(new_n330), .C2(new_n331), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n322), .A2(new_n326), .A3(G190), .A4(new_n327), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n360), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT73), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n435), .A2(new_n360), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n432), .A2(new_n433), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT73), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NOR4_X1   g0243(.A1(new_n380), .A2(new_n428), .A3(new_n429), .A4(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT89), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n310), .A2(new_n312), .A3(new_n208), .A4(G87), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(KEYINPUT88), .B2(KEYINPUT22), .ZN(new_n447));
  NOR2_X1   g0247(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n290), .A2(new_n208), .A3(G87), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT23), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n208), .B2(G107), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n373), .A2(KEYINPUT23), .A3(G20), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n453), .A2(new_n454), .B1(new_n257), .B2(G116), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT24), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT24), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n451), .A2(new_n458), .A3(new_n455), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n342), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n211), .A2(G33), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n272), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT25), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n268), .B2(G107), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n268), .A2(new_n463), .A3(G107), .ZN(new_n466));
  OAI22_X1  g0266(.A1(new_n462), .A2(new_n373), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n445), .B1(new_n460), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n281), .A2(G1), .ZN(new_n469));
  OR2_X1    g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n296), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  NOR2_X1   g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n473), .A2(G264), .B1(new_n477), .B2(new_n407), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n310), .A2(new_n312), .A3(G257), .A4(G1698), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n310), .A2(new_n312), .A3(G250), .A4(new_n291), .ZN(new_n480));
  INV_X1    g0280(.A(G294), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n479), .B(new_n480), .C1(new_n256), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n296), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n478), .A2(new_n483), .A3(G179), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT91), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n478), .A2(new_n483), .A3(KEYINPUT91), .A4(G179), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n478), .A2(new_n483), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT90), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(G169), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n490), .B1(new_n489), .B2(G169), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n451), .A2(new_n458), .A3(new_n455), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n458), .B1(new_n451), .B2(new_n455), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n254), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n467), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(KEYINPUT89), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n468), .A2(new_n494), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT92), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n478), .A2(new_n483), .A3(G190), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n489), .A2(G200), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n497), .A2(new_n498), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n500), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n501), .B1(new_n500), .B2(new_n504), .ZN(new_n506));
  OR2_X1    g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(G97), .A2(G107), .ZN(new_n508));
  NOR2_X1   g0308(.A1(G97), .A2(G107), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n508), .A2(new_n509), .B1(KEYINPUT78), .B2(KEYINPUT6), .ZN(new_n510));
  NOR2_X1   g0310(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g0311(.A(G97), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n511), .B1(KEYINPUT6), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g0313(.A(G97), .B(G107), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI22_X1  g0315(.A1(new_n515), .A2(new_n208), .B1(new_n220), .B2(new_n264), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT79), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT79), .ZN(new_n518));
  OAI221_X1 g0318(.A(new_n518), .B1(new_n220), .B2(new_n264), .C1(new_n515), .C2(new_n208), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n387), .A2(new_n389), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G107), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n517), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n254), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n310), .A2(new_n312), .A3(G250), .A4(G1698), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT81), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT81), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n290), .A2(new_n526), .A3(G250), .A4(G1698), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n310), .A2(new_n312), .A3(G244), .A4(new_n291), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT80), .ZN(new_n530));
  OR2_X1    g0330(.A1(new_n530), .A2(KEYINPUT4), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n290), .A2(G244), .A3(new_n531), .A4(new_n291), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G283), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n296), .B1(new_n528), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G274), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n476), .A2(new_n296), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT82), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n476), .A2(new_n284), .ZN(new_n541));
  INV_X1    g0341(.A(G257), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n476), .A2(KEYINPUT82), .A3(G257), .A4(new_n284), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n539), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n537), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G200), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n269), .A2(new_n512), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n462), .B2(new_n512), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n537), .A2(new_n545), .A3(G190), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n523), .A2(new_n547), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n537), .A2(new_n545), .A3(new_n299), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT83), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n537), .A2(new_n545), .A3(KEYINPUT83), .A4(new_n299), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n516), .A2(KEYINPUT79), .B1(G107), .B2(new_n520), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n342), .B1(new_n558), .B2(new_n519), .ZN(new_n559));
  INV_X1    g0359(.A(new_n546), .ZN(new_n560));
  OAI22_X1  g0360(.A1(new_n559), .A2(new_n549), .B1(new_n560), .B2(G169), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n552), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n214), .B1(new_n211), .B2(G33), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n352), .A2(new_n342), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n349), .A2(new_n214), .A3(new_n351), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n253), .A2(new_n207), .B1(G20), .B2(new_n214), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n535), .B(new_n208), .C1(G33), .C2(new_n512), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT20), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n566), .A2(KEYINPUT20), .A3(new_n567), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n564), .B(new_n565), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G179), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n311), .A2(G33), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n573));
  OAI21_X1  g0373(.A(G303), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n310), .A2(new_n312), .A3(G264), .A4(G1698), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n310), .A2(new_n312), .A3(G257), .A4(new_n291), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n296), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT87), .B1(new_n541), .B2(new_n215), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n477), .A2(new_n407), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT87), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n476), .A2(new_n581), .A3(G270), .A4(new_n284), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n571), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(G169), .A3(new_n570), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT21), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT21), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n583), .A2(new_n587), .A3(new_n570), .A4(G169), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n584), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n570), .B1(new_n583), .B2(G200), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n423), .B2(new_n583), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n310), .A2(new_n312), .A3(G238), .A4(new_n291), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n310), .A2(new_n312), .A3(G244), .A4(G1698), .ZN(new_n593));
  NAND2_X1  g0393(.A1(G33), .A2(G116), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n296), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n284), .A2(G274), .A3(new_n469), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n211), .A2(G45), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n284), .A2(G250), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n335), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n602), .A2(G179), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  XNOR2_X1  g0405(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n258), .B2(new_n512), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n290), .A2(new_n208), .A3(G68), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT19), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT84), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT84), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT19), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n315), .ZN(new_n615));
  AOI21_X1  g0415(.A(G20), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(G87), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n616), .A2(KEYINPUT85), .B1(new_n617), .B2(new_n509), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n208), .B1(new_n606), .B2(new_n315), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT85), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n609), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n364), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n622), .A2(new_n342), .B1(new_n352), .B2(new_n623), .ZN(new_n624));
  OR3_X1    g0424(.A1(new_n462), .A2(KEYINPUT86), .A3(new_n364), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT86), .B1(new_n462), .B2(new_n364), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n603), .B(new_n605), .C1(new_n624), .C2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n352), .A2(new_n623), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n462), .A2(new_n617), .ZN(new_n630));
  INV_X1    g0430(.A(new_n609), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n509), .A2(new_n617), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n619), .B2(new_n620), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n616), .A2(KEYINPUT85), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI211_X1 g0435(.A(new_n629), .B(new_n630), .C1(new_n635), .C2(new_n254), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n602), .A2(G200), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n600), .B1(new_n296), .B2(new_n595), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G190), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n589), .A2(new_n591), .A3(new_n628), .A4(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n562), .A2(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n444), .A2(new_n507), .A3(new_n643), .ZN(G372));
  INV_X1    g0444(.A(new_n379), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n361), .B1(new_n442), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n427), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n421), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n306), .A2(new_n308), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n300), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n444), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n557), .A2(new_n561), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n595), .A2(KEYINPUT93), .A3(new_n296), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT93), .B1(new_n595), .B2(new_n296), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n601), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G200), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n636), .A2(new_n639), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n335), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n658), .B(new_n605), .C1(new_n624), .C2(new_n627), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n652), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n523), .A2(new_n550), .B1(new_n335), .B2(new_n546), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n555), .A2(new_n556), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n628), .A2(new_n641), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT26), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n662), .A2(new_n659), .A3(new_n667), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n657), .A2(new_n659), .A3(new_n504), .ZN(new_n669));
  INV_X1    g0469(.A(new_n493), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n670), .A2(new_n491), .B1(new_n486), .B2(new_n487), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n460), .A2(new_n467), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n589), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AND4_X1   g0473(.A1(new_n665), .A2(new_n669), .A3(new_n552), .A4(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n650), .B1(new_n651), .B2(new_n675), .ZN(G369));
  NAND2_X1  g0476(.A1(new_n348), .A2(new_n208), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n468), .A2(new_n499), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n507), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n500), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n682), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n682), .A2(new_n570), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n589), .A2(new_n591), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n589), .B2(new_n689), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n671), .A2(new_n672), .ZN(new_n695));
  INV_X1    g0495(.A(new_n682), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n589), .A2(new_n682), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n507), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n694), .A2(new_n697), .A3(new_n699), .ZN(G399));
  NOR2_X1   g0500(.A1(new_n231), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n632), .A2(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n205), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n696), .B1(new_n668), .B2(new_n674), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT97), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT97), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n710), .B(new_n696), .C1(new_n668), .C2(new_n674), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n669), .A2(new_n665), .A3(new_n552), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n500), .A2(new_n589), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT98), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n657), .A2(new_n659), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT26), .B1(new_n665), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n629), .B1(new_n635), .B2(new_n254), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n625), .A2(new_n626), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n604), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n721), .A2(new_n603), .B1(new_n640), .B2(new_n636), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n722), .A2(new_n661), .A3(new_n664), .A4(new_n663), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n718), .A2(new_n659), .A3(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n562), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT98), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n726), .A3(new_n714), .A4(new_n669), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n716), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(KEYINPUT29), .A3(new_n696), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n712), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n643), .B(new_n696), .C1(new_n505), .C2(new_n506), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT94), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(KEYINPUT30), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n638), .A2(new_n578), .A3(new_n579), .A4(new_n582), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n484), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n734), .B1(new_n560), .B2(new_n736), .ZN(new_n737));
  NOR4_X1   g0537(.A1(new_n546), .A2(new_n735), .A3(new_n484), .A4(new_n733), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(G179), .B1(new_n478), .B2(new_n483), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n546), .A2(new_n583), .A3(new_n655), .A4(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT95), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n740), .A2(new_n583), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(KEYINPUT95), .A3(new_n546), .A4(new_n655), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n739), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n682), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n739), .A2(new_n741), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n696), .A2(new_n749), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n748), .A2(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n731), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(KEYINPUT96), .B1(new_n753), .B2(G330), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT96), .ZN(new_n755));
  INV_X1    g0555(.A(G330), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n755), .B(new_n756), .C1(new_n731), .C2(new_n752), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n730), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n706), .B1(new_n759), .B2(G1), .ZN(G364));
  INV_X1    g0560(.A(new_n692), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n230), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n211), .B1(new_n762), .B2(G45), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n702), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(G330), .B2(new_n691), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n232), .A2(new_n290), .ZN(new_n768));
  INV_X1    g0568(.A(G355), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n768), .A2(new_n769), .B1(G116), .B2(new_n232), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n248), .A2(new_n281), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n232), .A2(new_n388), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n281), .B2(new_n206), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n770), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n207), .B1(G20), .B2(new_n335), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n765), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n208), .A2(G179), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G190), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(G20), .A2(G179), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n783), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G329), .A2(new_n785), .B1(new_n789), .B2(G311), .ZN(new_n790));
  INV_X1    g0590(.A(G322), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n786), .A2(new_n423), .A3(G200), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n790), .B(new_n388), .C1(new_n791), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n787), .A2(G200), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G190), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(KEYINPUT33), .B(G317), .Z(new_n798));
  NAND3_X1  g0598(.A1(new_n782), .A2(G190), .A3(G200), .ZN(new_n799));
  INV_X1    g0599(.A(G303), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n797), .A2(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n794), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n795), .A2(new_n423), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G326), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n423), .A2(G179), .A3(G200), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n208), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n804), .B1(new_n481), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n782), .A2(new_n423), .A3(G200), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT99), .Z(new_n809));
  AOI22_X1  g0609(.A1(KEYINPUT100), .A2(new_n807), .B1(new_n809), .B2(G283), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n802), .B(new_n810), .C1(KEYINPUT100), .C2(new_n807), .ZN(new_n811));
  INV_X1    g0611(.A(new_n803), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n785), .A2(G159), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n812), .A2(new_n270), .B1(new_n813), .B2(KEYINPUT32), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n797), .A2(new_n225), .B1(new_n617), .B2(new_n799), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n809), .A2(G107), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n290), .B1(new_n793), .B2(new_n218), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G77), .B2(new_n789), .ZN(new_n819));
  INV_X1    g0619(.A(new_n806), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n813), .A2(KEYINPUT32), .B1(new_n820), .B2(G97), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n816), .A2(new_n817), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n811), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n781), .B1(new_n823), .B2(new_n778), .ZN(new_n824));
  INV_X1    g0624(.A(new_n777), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n691), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n767), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  NAND2_X1  g0628(.A1(new_n645), .A2(KEYINPUT102), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT102), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n379), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n829), .A2(new_n377), .A3(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n696), .B(new_n833), .C1(new_n668), .C2(new_n674), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n708), .A2(new_n711), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n370), .A2(new_n682), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n832), .A2(new_n838), .B1(new_n379), .B2(new_n696), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n834), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n765), .B1(new_n840), .B2(new_n758), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n758), .B2(new_n840), .ZN(new_n842));
  INV_X1    g0642(.A(new_n778), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n776), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n765), .B1(G77), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(G311), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n793), .A2(new_n481), .B1(new_n784), .B2(new_n846), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n290), .B(new_n847), .C1(G116), .C2(new_n789), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n809), .A2(G87), .ZN(new_n849));
  INV_X1    g0649(.A(new_n799), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n820), .A2(G97), .B1(new_n850), .B2(G107), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G283), .A2(new_n796), .B1(new_n803), .B2(G303), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n848), .A2(new_n849), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n789), .A2(G159), .B1(G143), .B2(new_n792), .ZN(new_n854));
  INV_X1    g0654(.A(G137), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n854), .B1(new_n797), .B2(new_n265), .C1(new_n855), .C2(new_n812), .ZN(new_n856));
  XNOR2_X1  g0656(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n809), .A2(G68), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n799), .A2(new_n270), .ZN(new_n860));
  INV_X1    g0660(.A(G132), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n290), .B1(new_n784), .B2(new_n861), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n860), .B(new_n862), .C1(G58), .C2(new_n820), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n858), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n856), .A2(new_n857), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n853), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n845), .B1(new_n866), .B2(new_n778), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n839), .B2(new_n776), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n842), .A2(new_n868), .ZN(G384));
  INV_X1    g0669(.A(KEYINPUT35), .ZN(new_n870));
  OAI211_X1 g0670(.A(G116), .B(new_n209), .C1(new_n515), .C2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n870), .B2(new_n515), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT36), .ZN(new_n873));
  OR3_X1    g0673(.A1(new_n205), .A2(new_n220), .A3(new_n382), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n270), .A2(G68), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n211), .B(G13), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n392), .A2(new_n254), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT7), .B1(new_n388), .B2(new_n208), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT75), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n225), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n387), .A2(new_n389), .A3(KEYINPUT75), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n384), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n883), .A2(KEYINPUT16), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n401), .B1(new_n878), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n680), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n421), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n888), .B1(new_n889), .B2(new_n647), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT105), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT104), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n398), .B1(new_n278), .B2(new_n397), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n342), .B1(new_n883), .B2(KEYINPUT16), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n385), .B1(new_n390), .B2(new_n391), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n393), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n893), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n417), .A2(new_n299), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n898), .A2(new_n414), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n426), .B(new_n892), .C1(new_n897), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n887), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n885), .A2(new_n418), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n892), .B1(new_n902), .B2(new_n426), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n891), .B(KEYINPUT37), .C1(new_n901), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n402), .A2(new_n886), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n419), .A2(new_n905), .A3(new_n426), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n906), .A2(KEYINPUT37), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n894), .A2(new_n896), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n899), .B1(new_n909), .B2(new_n401), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n396), .A2(new_n425), .A3(new_n401), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT104), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(new_n887), .A3(new_n900), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n891), .B1(new_n913), .B2(KEYINPUT37), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n890), .B1(new_n908), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(KEYINPUT38), .B(new_n890), .C1(new_n908), .C2(new_n914), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n917), .A2(KEYINPUT39), .A3(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n906), .B(KEYINPUT37), .Z(new_n920));
  AOI21_X1  g0720(.A(new_n905), .B1(new_n421), .B2(new_n427), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT103), .B1(new_n341), .B2(new_n360), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n328), .A2(new_n332), .ZN(new_n927));
  INV_X1    g0727(.A(new_n340), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT74), .B1(new_n339), .B2(KEYINPUT14), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT103), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n930), .A2(new_n931), .A3(new_n359), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n682), .B1(new_n926), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n919), .A2(new_n925), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n917), .A2(new_n918), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n926), .A2(new_n932), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n359), .A2(new_n682), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n440), .B1(new_n438), .B2(new_n439), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n930), .B1(new_n437), .B2(new_n441), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n936), .A2(new_n940), .B1(new_n941), .B2(new_n937), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n829), .A2(new_n831), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n696), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n943), .B1(new_n834), .B2(new_n945), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n935), .A2(new_n946), .B1(new_n889), .B2(new_n680), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n934), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n650), .B1(new_n730), .B2(new_n651), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n918), .A2(new_n922), .ZN(new_n951));
  NOR2_X1   g0751(.A1(KEYINPUT106), .A2(KEYINPUT31), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n747), .B2(new_n682), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n696), .B(new_n952), .C1(new_n739), .C2(new_n746), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n731), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n957), .A2(new_n839), .A3(new_n942), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT40), .B1(new_n951), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT40), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n957), .A2(new_n960), .A3(new_n942), .A4(new_n839), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n935), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n444), .A2(new_n957), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n756), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n965), .B2(new_n964), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n950), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n211), .B2(new_n762), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n950), .A2(new_n967), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n877), .B1(new_n969), .B2(new_n970), .ZN(G367));
  AND3_X1   g0771(.A1(new_n240), .A2(new_n232), .A3(new_n388), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n779), .B1(new_n232), .B2(new_n364), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n765), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(G143), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n812), .A2(new_n975), .B1(new_n799), .B2(new_n218), .ZN(new_n976));
  INV_X1    g0776(.A(new_n808), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n976), .B1(G77), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n388), .B1(G150), .B2(new_n792), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G137), .A2(new_n785), .B1(new_n789), .B2(G50), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n820), .A2(G68), .B1(new_n796), .B2(G159), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n978), .A2(new_n979), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G294), .A2(new_n796), .B1(new_n977), .B2(G97), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n373), .B2(new_n806), .C1(new_n846), .C2(new_n812), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n850), .A2(KEYINPUT46), .A3(G116), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n789), .A2(G283), .B1(G303), .B2(new_n792), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n290), .B1(new_n785), .B2(G317), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT46), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n799), .B2(new_n214), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n985), .A2(new_n986), .A3(new_n987), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n982), .B1(new_n984), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT115), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT47), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n974), .B1(new_n993), .B2(new_n778), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n636), .A2(new_n696), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n995), .A2(new_n721), .A3(new_n658), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n717), .B2(new_n995), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n994), .B1(new_n825), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n763), .B(KEYINPUT114), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n652), .A2(new_n682), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(KEYINPUT107), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(KEYINPUT107), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n682), .B1(new_n559), .B2(new_n549), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n1002), .A2(new_n1003), .B1(new_n725), .B2(new_n1004), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n507), .A2(new_n698), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n697), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT44), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n725), .A2(new_n1004), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1012), .A2(new_n697), .A3(new_n699), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT112), .Z(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1013), .B(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n693), .B1(new_n1009), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT44), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1008), .B(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1013), .B(new_n1015), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(new_n1021), .A3(new_n694), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1006), .B1(KEYINPUT113), .B2(new_n692), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT113), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n761), .A2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1023), .B(new_n1025), .C1(new_n687), .C2(new_n698), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n687), .A2(new_n698), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1024), .B(new_n761), .C1(new_n1027), .C2(new_n1006), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1018), .A2(new_n1022), .A3(new_n759), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n759), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(KEYINPUT110), .B(KEYINPUT41), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n701), .B(new_n1032), .Z(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1000), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(KEYINPUT42), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n652), .B1(new_n1012), .B2(new_n685), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1038), .B1(new_n682), .B2(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1040), .A2(KEYINPUT108), .B1(KEYINPUT42), .B2(new_n1037), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1040), .A2(KEYINPUT108), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1036), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n687), .A2(new_n761), .A3(new_n1012), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1044), .A2(KEYINPUT109), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(KEYINPUT109), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1045), .B(new_n1046), .C1(KEYINPUT43), .C2(new_n997), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1043), .B(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n998), .B1(new_n1035), .B2(new_n1052), .ZN(G387));
  NOR2_X1   g0853(.A1(new_n1029), .A2(new_n759), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1029), .A2(new_n759), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n701), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1054), .B1(new_n1056), .B2(KEYINPUT118), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(KEYINPUT118), .B2(new_n1056), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n768), .A2(new_n703), .B1(G107), .B2(new_n232), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n772), .B1(new_n244), .B2(G45), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n281), .B1(new_n225), .B2(new_n220), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n703), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1061), .B1(new_n1062), .B2(KEYINPUT116), .ZN(new_n1063));
  AND3_X1   g0863(.A1(new_n397), .A2(KEYINPUT50), .A3(new_n270), .ZN(new_n1064));
  AOI21_X1  g0864(.A(KEYINPUT50), .B1(new_n397), .B2(new_n270), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1063), .B1(KEYINPUT116), .B2(new_n1062), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1059), .B1(new_n1060), .B2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n789), .A2(G68), .B1(G50), .B2(new_n792), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1068), .B(new_n290), .C1(new_n265), .C2(new_n784), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n806), .A2(new_n364), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G159), .B2(new_n803), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n220), .B2(new_n799), .C1(new_n259), .C2(new_n797), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1069), .B(new_n1072), .C1(G97), .C2(new_n809), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n789), .A2(G303), .B1(G317), .B2(new_n792), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n797), .B2(new_n846), .C1(new_n791), .C2(new_n812), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT117), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT48), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n820), .A2(G283), .B1(new_n850), .B2(G294), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1082), .A2(KEYINPUT49), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n290), .B1(new_n785), .B2(G326), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n214), .B2(new_n808), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n1082), .B2(KEYINPUT49), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1073), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n765), .B1(new_n780), .B2(new_n1067), .C1(new_n1087), .C2(new_n843), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n688), .B2(new_n777), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n1029), .B2(new_n1000), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1058), .A2(new_n1090), .ZN(G393));
  NAND2_X1  g0891(.A1(new_n1018), .A2(new_n1022), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT119), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1018), .A2(new_n1022), .A3(KEYINPUT119), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n1000), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1092), .A2(new_n1055), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(new_n701), .A3(new_n1030), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n779), .B1(new_n512), .B2(new_n232), .C1(new_n251), .C2(new_n772), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n765), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n799), .A2(new_n225), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n806), .A2(new_n220), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(G50), .C2(new_n796), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n290), .B1(new_n784), .B2(new_n975), .C1(new_n259), .C2(new_n788), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1103), .A2(new_n849), .A3(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n803), .A2(G150), .B1(G159), .B2(new_n792), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT51), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n388), .B1(new_n788), .B2(new_n481), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G322), .B2(new_n785), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n820), .A2(G116), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G303), .A2(new_n796), .B1(new_n850), .B2(G283), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n817), .A2(new_n1110), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n803), .A2(G317), .B1(G311), .B2(new_n792), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT52), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1106), .A2(new_n1108), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1100), .B1(new_n1116), .B2(new_n778), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n1012), .B2(new_n825), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1096), .A2(new_n1098), .A3(new_n1118), .ZN(G390));
  AOI21_X1  g0919(.A(new_n776), .B1(new_n919), .B2(new_n925), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n793), .A2(new_n214), .B1(new_n784), .B2(new_n481), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n290), .B(new_n1121), .C1(G97), .C2(new_n789), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1102), .B1(G87), .B2(new_n850), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(G107), .A2(new_n796), .B1(new_n803), .B2(G283), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1122), .A2(new_n859), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT54), .B(G143), .ZN(new_n1126));
  INV_X1    g0926(.A(G125), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n788), .A2(new_n1126), .B1(new_n784), .B2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n388), .B(new_n1128), .C1(G132), .C2(new_n792), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n799), .A2(new_n265), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT53), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n820), .A2(G159), .B1(new_n796), .B2(G137), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G128), .A2(new_n803), .B1(new_n977), .B2(G50), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n843), .B1(new_n1125), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n765), .B1(new_n397), .B2(new_n844), .ZN(new_n1136));
  OR3_X1    g0936(.A1(new_n1120), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n834), .A2(new_n945), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n933), .B1(new_n1138), .B2(new_n942), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n917), .A2(KEYINPUT39), .A3(new_n918), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT39), .B1(new_n918), .B2(new_n922), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n728), .A2(new_n696), .A3(new_n833), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n943), .B1(new_n1144), .B2(new_n945), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n933), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n923), .A2(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n839), .B(new_n942), .C1(new_n754), .C2(new_n757), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1143), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n756), .B1(new_n956), .B2(new_n731), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1151), .A2(new_n839), .A3(new_n942), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1139), .B1(new_n919), .B2(new_n925), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1150), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1137), .B1(new_n1157), .B2(new_n999), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1144), .A2(new_n945), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n942), .B1(new_n1151), .B2(new_n839), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n1149), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n839), .B1(new_n754), .B2(new_n757), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1153), .B1(new_n1163), .B2(new_n943), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1138), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1162), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n444), .A2(new_n1151), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1167), .B(new_n650), .C1(new_n730), .C2(new_n651), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n702), .B1(new_n1170), .B2(new_n1157), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1166), .A2(new_n1150), .A3(new_n1156), .A4(new_n1169), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1158), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(G378));
  NAND2_X1  g0974(.A1(new_n279), .A2(new_n886), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n309), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n309), .A2(new_n1175), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1179), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n964), .B2(G330), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n957), .A2(new_n839), .A3(new_n942), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n960), .B1(new_n1184), .B2(new_n923), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n961), .B1(new_n918), .B2(new_n917), .ZN(new_n1186));
  OAI211_X1 g0986(.A(G330), .B(new_n1182), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n948), .B1(new_n1183), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1182), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1190), .B1(new_n1191), .B2(new_n756), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n948), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1192), .A2(new_n1193), .A3(new_n1187), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1189), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1190), .A2(new_n775), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n765), .B1(G50), .B2(new_n844), .ZN(new_n1197));
  INV_X1    g0997(.A(G128), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n793), .A2(new_n1198), .B1(new_n788), .B2(new_n855), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n803), .A2(G125), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n799), .B2(new_n1126), .C1(new_n797), .C2(new_n861), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1199), .B(new_n1201), .C1(G150), .C2(new_n820), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n977), .A2(G159), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G33), .B(G41), .C1(new_n785), .C2(G124), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n812), .A2(new_n214), .B1(new_n808), .B2(new_n218), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n388), .A2(new_n280), .ZN(new_n1210));
  INV_X1    g1010(.A(G283), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n793), .A2(new_n373), .B1(new_n784), .B2(new_n1211), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1210), .B(new_n1212), .C1(new_n623), .C2(new_n789), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n820), .A2(G68), .B1(new_n850), .B2(G77), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1209), .B(new_n1215), .C1(G97), .C2(new_n796), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT58), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1210), .B(new_n270), .C1(G33), .C2(G41), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1216), .A2(KEYINPUT58), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1208), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1197), .B1(new_n1220), .B2(new_n778), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1195), .A2(new_n1000), .B1(new_n1196), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1163), .A2(new_n943), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n1152), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1224), .A2(new_n1138), .B1(new_n1149), .B2(new_n1161), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1169), .B1(new_n1157), .B2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1195), .A2(KEYINPUT57), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n701), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1226), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1222), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT120), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(KEYINPUT120), .B(new_n1222), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(G375));
  OAI211_X1 g1035(.A(new_n1168), .B(new_n1162), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1170), .A2(new_n1034), .A3(new_n1236), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT121), .Z(new_n1238));
  NAND2_X1  g1038(.A1(new_n943), .A2(new_n775), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n765), .B1(G68), .B2(new_n844), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n812), .A2(new_n481), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1070), .B(new_n1241), .C1(G116), .C2(new_n796), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n799), .A2(new_n512), .B1(new_n784), .B2(new_n800), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT122), .Z(new_n1244));
  NAND2_X1  g1044(.A1(new_n809), .A2(G77), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n388), .B1(new_n793), .B2(new_n1211), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G107), .B2(new_n789), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1242), .A2(new_n1244), .A3(new_n1245), .A4(new_n1247), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n806), .A2(new_n270), .B1(new_n788), .B2(new_n265), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1249), .B(KEYINPUT123), .Z(new_n1250));
  OAI22_X1  g1050(.A1(new_n812), .A2(new_n861), .B1(new_n808), .B2(new_n218), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n850), .A2(G159), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n797), .B2(new_n1126), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n290), .B1(new_n784), .B2(new_n1198), .C1(new_n793), .C2(new_n855), .ZN(new_n1254));
  OR3_X1    g1054(.A1(new_n1251), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1248), .B1(new_n1250), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1240), .B1(new_n1256), .B2(new_n778), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1166), .A2(new_n1000), .B1(new_n1239), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1238), .A2(new_n1258), .ZN(G381));
  AND3_X1   g1059(.A1(new_n1096), .A2(new_n1098), .A3(new_n1118), .ZN(new_n1260));
  INV_X1    g1060(.A(G384), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1043), .A2(new_n1051), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1043), .A2(new_n1051), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1033), .B1(new_n1030), .B2(new_n759), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1262), .B(new_n1263), .C1(new_n1264), .C2(new_n1000), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1260), .A2(new_n1261), .A3(new_n1265), .A4(new_n998), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1058), .A2(new_n827), .A3(new_n1090), .ZN(new_n1267));
  NOR4_X1   g1067(.A1(new_n1266), .A2(G381), .A3(G378), .A4(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1234), .ZN(G407));
  INV_X1    g1069(.A(G213), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1270), .A2(G343), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1234), .A2(new_n1173), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT124), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1272), .B(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(G213), .A3(G407), .ZN(G409));
  NAND2_X1  g1075(.A1(G393), .A2(G396), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1267), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(G387), .A2(new_n1260), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G390), .B1(new_n1265), .B2(new_n998), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1277), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G387), .A2(new_n1260), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1265), .A2(G390), .A3(new_n998), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1267), .A3(new_n1276), .A4(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1195), .A2(new_n1034), .A3(new_n1226), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT125), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT125), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1195), .A2(new_n1226), .A3(new_n1287), .A4(new_n1034), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1286), .A2(new_n1222), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1173), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G378), .B(new_n1222), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1271), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1236), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(KEYINPUT60), .B2(new_n1170), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1225), .A2(KEYINPUT60), .A3(new_n1168), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n701), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1258), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1261), .ZN(new_n1300));
  OAI211_X1 g1100(.A(G384), .B(new_n1258), .C1(new_n1296), .C2(new_n1298), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1292), .A2(new_n1293), .A3(new_n1294), .A4(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1271), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1271), .A2(G2897), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1302), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(G2897), .A3(new_n1271), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1303), .B(new_n1304), .C1(new_n1305), .C2(new_n1310), .ZN(new_n1311));
  AOI211_X1 g1111(.A(new_n1271), .B(new_n1308), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1312), .A2(new_n1293), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1284), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1280), .A2(new_n1304), .A3(new_n1283), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1315), .B1(new_n1312), .B2(KEYINPUT63), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT126), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1317), .A2(new_n1318), .A3(new_n1307), .A4(new_n1309), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT63), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1320), .B1(new_n1317), .B2(new_n1308), .ZN(new_n1321));
  OAI21_X1  g1121(.A(KEYINPUT126), .B1(new_n1310), .B2(new_n1305), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1316), .A2(new_n1319), .A3(new_n1321), .A4(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1314), .A2(new_n1323), .ZN(G405));
  NAND2_X1  g1124(.A1(new_n1302), .A2(KEYINPUT127), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1232), .A2(new_n1233), .A3(new_n1173), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1284), .A2(new_n1291), .A3(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1284), .B1(new_n1291), .B2(new_n1326), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1325), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1326), .A2(new_n1291), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1331), .A2(new_n1283), .A3(new_n1280), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1332), .A2(KEYINPUT127), .A3(new_n1302), .A4(new_n1327), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1330), .A2(new_n1333), .ZN(G402));
endmodule


