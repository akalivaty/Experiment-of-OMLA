//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G116), .A2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  INV_X1    g0008(.A(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n202), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n212), .B(new_n217), .C1(G97), .C2(G257), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G1), .B2(G20), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n220));
  XNOR2_X1  g0020(.A(new_n219), .B(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NOR3_X1   g0029(.A1(new_n221), .A2(new_n225), .A3(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G87), .B(G116), .ZN(new_n239));
  INV_X1    g0039(.A(G107), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G97), .ZN(new_n241));
  INV_X1    g0041(.A(G97), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G107), .ZN(new_n243));
  NAND3_X1  g0043(.A1(new_n239), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G97), .B(G107), .ZN(new_n245));
  OAI21_X1  g0045(.A(new_n244), .B1(new_n239), .B2(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n246), .B(KEYINPUT66), .Z(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G1698), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n252), .A2(G222), .A3(new_n255), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n254), .A2(G223), .B1(new_n256), .B2(KEYINPUT69), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n257), .B1(KEYINPUT69), .B2(new_n256), .C1(new_n208), .C2(new_n252), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT67), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G45), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n263), .B(G274), .C1(new_n268), .C2(G41), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT68), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n260), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n270), .B1(new_n260), .B2(new_n271), .ZN(new_n273));
  OAI21_X1  g0073(.A(G226), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n262), .A2(new_n269), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G200), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT74), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n262), .A2(G190), .A3(new_n269), .A4(new_n274), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT10), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n276), .A2(new_n278), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT9), .ZN(new_n283));
  INV_X1    g0083(.A(G13), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n284), .A2(new_n223), .A3(G1), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n202), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT70), .B1(new_n226), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT70), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n290), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n263), .A2(G20), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n289), .A2(new_n224), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n287), .B1(new_n294), .B2(new_n202), .ZN(new_n295));
  XOR2_X1   g0095(.A(new_n295), .B(KEYINPUT73), .Z(new_n296));
  NAND2_X1  g0096(.A1(new_n203), .A2(G20), .ZN(new_n297));
  INV_X1    g0097(.A(G150), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G58), .ZN(new_n301));
  AOI21_X1  g0101(.A(KEYINPUT71), .B1(new_n301), .B2(KEYINPUT8), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT71), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT8), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n302), .A2(new_n305), .B1(KEYINPUT72), .B2(new_n301), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT72), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n307), .B(G58), .C1(new_n303), .C2(new_n304), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n223), .A2(G33), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n297), .B1(new_n298), .B2(new_n300), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n289), .A2(new_n224), .A3(new_n291), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n283), .B1(new_n296), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n296), .B1(new_n312), .B2(new_n311), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT9), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n281), .A2(new_n282), .A3(new_n315), .A4(new_n317), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n317), .A2(new_n276), .A3(new_n278), .A4(new_n315), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(new_n280), .A3(new_n279), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n316), .B1(new_n321), .B2(new_n275), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(G179), .B2(new_n275), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n318), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT11), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n310), .A2(new_n208), .B1(new_n223), .B2(G68), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT75), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT75), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n328), .B1(new_n223), .B2(G68), .C1(new_n310), .C2(new_n208), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n327), .B(new_n329), .C1(new_n202), .C2(new_n300), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT76), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(new_n331), .A3(new_n312), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n331), .B1(new_n330), .B2(new_n312), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n325), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n334), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT11), .A3(new_n332), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n284), .A2(G1), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(G20), .A3(new_n215), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n340), .A2(KEYINPUT12), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n294), .A2(G68), .B1(KEYINPUT12), .B2(new_n340), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n335), .A2(new_n337), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT77), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT14), .ZN(new_n345));
  OAI21_X1  g0145(.A(G238), .B1(new_n272), .B2(new_n273), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n288), .A2(KEYINPUT3), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n214), .A2(new_n255), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT3), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G33), .ZN(new_n350));
  INV_X1    g0150(.A(G232), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G1698), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n347), .A2(new_n348), .A3(new_n350), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n261), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n346), .A2(new_n356), .A3(new_n269), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT13), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT13), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n346), .A2(new_n356), .A3(new_n359), .A4(new_n269), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n345), .B1(new_n361), .B2(G169), .ZN(new_n362));
  AOI211_X1 g0162(.A(KEYINPUT14), .B(new_n321), .C1(new_n358), .C2(new_n360), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n358), .A2(G179), .A3(new_n360), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n344), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NOR4_X1   g0167(.A1(new_n362), .A2(new_n363), .A3(KEYINPUT77), .A4(new_n365), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n343), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n347), .A2(new_n350), .A3(new_n255), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n253), .A2(new_n216), .B1(new_n351), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n252), .A2(new_n240), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n261), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(G244), .B1(new_n272), .B2(new_n273), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n269), .A3(new_n374), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n375), .A2(G179), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n321), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT8), .B(G58), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT15), .B(G87), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n300), .A2(new_n378), .B1(new_n379), .B2(new_n310), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n223), .A2(new_n208), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n312), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n285), .A2(new_n208), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n294), .A2(G77), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n376), .A2(new_n377), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n375), .A2(G200), .ZN(new_n387));
  INV_X1    g0187(.A(new_n385), .ZN(new_n388));
  INV_X1    g0188(.A(G190), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n387), .B(new_n388), .C1(new_n389), .C2(new_n375), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n369), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n324), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n309), .A2(new_n286), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n306), .A2(new_n308), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n293), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT80), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT80), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(new_n398), .A3(new_n395), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n301), .A2(new_n215), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n401), .A2(new_n201), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(G20), .B1(G159), .B2(new_n299), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n347), .A2(new_n350), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT78), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT7), .B1(new_n404), .B2(new_n223), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT7), .ZN(new_n410));
  OAI211_X1 g0210(.A(KEYINPUT78), .B(new_n410), .C1(new_n252), .C2(G20), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G68), .ZN(new_n412));
  OAI211_X1 g0212(.A(KEYINPUT16), .B(new_n403), .C1(new_n409), .C2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT16), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n404), .A2(new_n223), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n410), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT79), .B1(new_n349), .B2(G33), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT79), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(new_n288), .A3(KEYINPUT3), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n419), .A3(new_n350), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n215), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n403), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n414), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n413), .A2(new_n424), .A3(new_n312), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n400), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n252), .B1(G223), .B2(G1698), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n255), .A2(G226), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n427), .A2(new_n428), .B1(new_n288), .B2(new_n210), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n261), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n260), .A2(G232), .A3(new_n271), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n430), .A2(new_n431), .A3(new_n269), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G190), .ZN(new_n433));
  AOI21_X1  g0233(.A(G41), .B1(new_n265), .B2(new_n267), .ZN(new_n434));
  INV_X1    g0234(.A(G274), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n434), .A2(G1), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(new_n429), .B2(new_n261), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n431), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G200), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n426), .A2(KEYINPUT17), .A3(new_n433), .A4(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n400), .A2(new_n433), .A3(new_n425), .A4(new_n439), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT17), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n400), .A2(new_n425), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n438), .A2(G169), .ZN(new_n445));
  INV_X1    g0245(.A(G179), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n445), .B1(new_n446), .B2(new_n438), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n444), .A2(new_n447), .A3(KEYINPUT18), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT18), .B1(new_n444), .B2(new_n447), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n440), .B(new_n443), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n361), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G190), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n343), .B1(G200), .B2(new_n361), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n392), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n286), .A2(G97), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n288), .A2(G1), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n312), .A2(new_n285), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n456), .B1(new_n458), .B2(G97), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT6), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n241), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n462), .B1(new_n461), .B2(new_n245), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(new_n223), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n300), .A2(new_n208), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n416), .A2(new_n421), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n465), .B(new_n467), .C1(new_n468), .C2(new_n240), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n460), .B1(new_n469), .B2(new_n312), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n264), .A2(G1), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  AND2_X1   g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n471), .B(G274), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n471), .B1(new_n473), .B2(new_n472), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n260), .ZN(new_n476));
  INV_X1    g0276(.A(G257), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT4), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(KEYINPUT81), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT81), .ZN(new_n482));
  OAI21_X1  g0282(.A(G244), .B1(new_n482), .B2(KEYINPUT4), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n481), .B1(new_n370), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n252), .A2(G250), .A3(G1698), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n209), .B1(KEYINPUT81), .B2(new_n479), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n252), .A2(new_n487), .A3(new_n255), .A4(new_n480), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n478), .B1(new_n489), .B2(new_n261), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G190), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n261), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT82), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT82), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n489), .A2(new_n494), .A3(new_n261), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n478), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G200), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n470), .B(new_n491), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n458), .A2(G87), .ZN(new_n499));
  NOR2_X1   g0299(.A1(G97), .A2(G107), .ZN(new_n500));
  AND2_X1   g0300(.A1(KEYINPUT84), .A2(G87), .ZN(new_n501));
  NOR2_X1   g0301(.A1(KEYINPUT84), .A2(G87), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n354), .A2(new_n223), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n503), .A2(KEYINPUT19), .A3(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n347), .A2(new_n350), .A3(new_n223), .A4(G68), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n354), .A2(G20), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n506), .B1(KEYINPUT19), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n312), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n379), .A2(new_n285), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n499), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n209), .A2(G1698), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(G238), .B2(G1698), .ZN(new_n513));
  INV_X1    g0313(.A(G116), .ZN(new_n514));
  OAI22_X1  g0314(.A1(new_n513), .A2(new_n404), .B1(new_n288), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n261), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n260), .A2(G250), .ZN(new_n517));
  INV_X1    g0317(.A(new_n471), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n264), .A2(G1), .A3(G274), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT83), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n471), .B1(new_n260), .B2(G250), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT83), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n523), .A2(new_n524), .A3(new_n520), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n516), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G200), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n519), .A2(KEYINPUT83), .A3(new_n521), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n524), .B1(new_n523), .B2(new_n520), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n528), .A2(new_n529), .B1(new_n261), .B2(new_n515), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G190), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n511), .A2(new_n527), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n379), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n458), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(new_n509), .A3(new_n510), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n516), .B(new_n446), .C1(new_n522), .C2(new_n525), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n535), .B(new_n536), .C1(new_n530), .C2(G169), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n478), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n489), .A2(new_n494), .A3(new_n261), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n494), .B1(new_n489), .B2(new_n261), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n446), .B(new_n539), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n240), .B1(new_n416), .B2(new_n421), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n543), .A2(new_n464), .A3(new_n466), .ZN(new_n544));
  INV_X1    g0344(.A(new_n312), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n459), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n490), .A2(G169), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n542), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n240), .A2(G20), .ZN(new_n549));
  XNOR2_X1  g0349(.A(new_n549), .B(KEYINPUT23), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n347), .A2(new_n350), .A3(new_n223), .A4(G87), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT22), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT22), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n252), .A2(new_n553), .A3(new_n223), .A4(G87), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n550), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT24), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n223), .A2(G33), .A3(G116), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n556), .B1(new_n555), .B2(new_n557), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n312), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT86), .B1(new_n370), .B2(new_n211), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n252), .A2(G257), .A3(G1698), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT86), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n252), .A2(new_n564), .A3(G250), .A4(new_n255), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G294), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n562), .A2(new_n563), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n261), .ZN(new_n568));
  INV_X1    g0368(.A(new_n476), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G264), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n474), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G200), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n567), .A2(new_n261), .B1(G264), .B2(new_n569), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(G190), .A3(new_n474), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n458), .A2(G107), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n338), .A2(G20), .A3(new_n240), .ZN(new_n576));
  XNOR2_X1  g0376(.A(new_n576), .B(KEYINPUT25), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n561), .A2(new_n572), .A3(new_n574), .A4(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n498), .A2(new_n538), .A3(new_n548), .A4(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n485), .B(new_n223), .C1(G33), .C2(new_n242), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n514), .A2(G20), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n312), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT20), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n312), .A2(KEYINPUT20), .A3(new_n581), .A4(new_n582), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n263), .A2(new_n514), .A3(G13), .A4(G20), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n588), .B(KEYINPUT85), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n458), .B2(G116), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n255), .A2(G257), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G264), .A2(G1698), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n347), .A2(new_n350), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n594), .B(new_n261), .C1(G303), .C2(new_n252), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n475), .A2(G270), .A3(new_n260), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n474), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n597), .A2(G169), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n591), .A2(new_n598), .A3(KEYINPUT21), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT21), .B1(new_n591), .B2(new_n598), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n571), .A2(new_n321), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n573), .A2(new_n446), .A3(new_n474), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n552), .A2(new_n554), .ZN(new_n604));
  INV_X1    g0404(.A(new_n550), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n557), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT24), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n545), .B1(new_n607), .B2(new_n558), .ZN(new_n608));
  INV_X1    g0408(.A(new_n578), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n602), .B(new_n603), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n597), .A2(new_n446), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n591), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n597), .A2(G200), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n389), .B2(new_n597), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n614), .A2(new_n591), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n601), .A2(new_n610), .A3(new_n612), .A4(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n455), .A2(new_n580), .A3(new_n616), .ZN(G372));
  INV_X1    g0417(.A(new_n323), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n441), .B(KEYINPUT17), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n453), .A2(new_n452), .ZN(new_n620));
  INV_X1    g0420(.A(new_n377), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n385), .B1(new_n375), .B2(G179), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT88), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT88), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n376), .A2(new_n624), .A3(new_n377), .A4(new_n385), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n369), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n619), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT18), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n321), .B1(new_n437), .B2(new_n431), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(G179), .B2(new_n432), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n630), .B1(new_n426), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n444), .A2(new_n447), .A3(KEYINPUT18), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n318), .A2(new_n320), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n618), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n532), .A2(new_n537), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT26), .B1(new_n548), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n542), .A2(new_n547), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT87), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT87), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n542), .A2(new_n643), .A3(new_n547), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n642), .A2(new_n546), .A3(new_n538), .A4(new_n644), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n537), .B(new_n640), .C1(new_n645), .C2(KEYINPUT26), .ZN(new_n646));
  INV_X1    g0446(.A(new_n610), .ZN(new_n647));
  INV_X1    g0447(.A(new_n600), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n591), .A2(new_n598), .A3(KEYINPUT21), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(new_n612), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n579), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n498), .A2(new_n538), .A3(new_n548), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n638), .B1(new_n455), .B2(new_n654), .ZN(G369));
  NOR2_X1   g0455(.A1(new_n284), .A2(G20), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(new_n263), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n263), .A2(new_n223), .A3(G13), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n658), .A2(new_n660), .A3(G213), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT89), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT89), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n658), .A2(new_n660), .A3(new_n663), .A4(G213), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT90), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT90), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n610), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n608), .B2(new_n609), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n579), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n671), .B1(new_n673), .B2(new_n610), .ZN(new_n674));
  AOI211_X1 g0474(.A(new_n446), .B(new_n597), .C1(new_n587), .C2(new_n590), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n599), .A2(new_n600), .A3(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(new_n670), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n671), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT91), .Z(new_n679));
  NAND2_X1  g0479(.A1(new_n670), .A2(new_n591), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n676), .B(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n681), .A2(new_n615), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n674), .A2(new_n677), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n674), .A2(new_n677), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n679), .A2(new_n686), .ZN(G399));
  OR2_X1    g0487(.A1(new_n501), .A2(new_n502), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(new_n514), .A3(new_n500), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT92), .ZN(new_n690));
  INV_X1    g0490(.A(new_n227), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G41), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n690), .A2(new_n263), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n222), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n692), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT28), .Z(new_n696));
  INV_X1    g0496(.A(KEYINPUT29), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n561), .A2(new_n574), .A3(new_n578), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n676), .A2(new_n610), .B1(new_n698), .B2(new_n572), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT98), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n498), .A2(new_n700), .A3(new_n548), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n700), .B1(new_n498), .B2(new_n548), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n699), .B(new_n532), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT26), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n548), .B2(new_n639), .ZN(new_n705));
  OAI211_X1 g0505(.A(KEYINPUT97), .B(new_n705), .C1(new_n645), .C2(new_n704), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n542), .A2(new_n643), .A3(new_n547), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n643), .B1(new_n542), .B2(new_n547), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n707), .A2(new_n708), .A3(new_n470), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT97), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n709), .A2(new_n710), .A3(KEYINPUT26), .A4(new_n538), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n703), .A2(new_n706), .A3(new_n537), .A4(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n670), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n697), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n646), .B2(new_n653), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT96), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g0517(.A(KEYINPUT96), .B(new_n713), .C1(new_n646), .C2(new_n653), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n714), .B1(new_n719), .B2(new_n697), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n580), .A2(new_n616), .A3(new_n670), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n526), .A2(new_n446), .A3(new_n597), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(new_n724), .A3(new_n571), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT95), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n573), .A2(new_n611), .A3(new_n490), .A4(new_n530), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  OAI21_X1  g0529(.A(KEYINPUT94), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n728), .A2(KEYINPUT94), .A3(new_n729), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n670), .B1(new_n727), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n721), .B1(new_n722), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n713), .A2(new_n722), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n728), .A2(new_n729), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(new_n725), .A3(new_n731), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT93), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n736), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G330), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n720), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n696), .B1(new_n746), .B2(G1), .ZN(G364));
  XOR2_X1   g0547(.A(new_n683), .B(KEYINPUT99), .Z(new_n748));
  NOR3_X1   g0548(.A1(new_n284), .A2(new_n264), .A3(G20), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(KEYINPUT100), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(KEYINPUT100), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(G1), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n692), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n748), .B(new_n754), .C1(G330), .C2(new_n682), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT101), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n223), .A2(new_n446), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(G190), .A3(new_n497), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT104), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(G190), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n497), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n759), .A2(G58), .B1(G50), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G190), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n757), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n762), .B1(new_n208), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT105), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n223), .A2(G179), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(new_n389), .A3(G200), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT106), .Z(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n240), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n446), .A2(new_n497), .A3(G190), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n242), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n757), .A2(new_n389), .A3(G200), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n767), .A2(G190), .A3(G200), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n252), .B1(new_n775), .B2(new_n215), .C1(new_n688), .C2(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n770), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n767), .A2(new_n763), .ZN(new_n779));
  INV_X1    g0579(.A(G159), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT32), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n766), .A2(new_n778), .A3(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G311), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n764), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n769), .ZN(new_n786));
  INV_X1    g0586(.A(new_n761), .ZN(new_n787));
  INV_X1    g0587(.A(G326), .ZN(new_n788));
  INV_X1    g0588(.A(G294), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n787), .A2(new_n788), .B1(new_n789), .B2(new_n773), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n786), .A2(G283), .B1(new_n790), .B2(KEYINPUT107), .ZN(new_n791));
  XOR2_X1   g0591(.A(KEYINPUT33), .B(G317), .Z(new_n792));
  NOR2_X1   g0592(.A1(new_n775), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n779), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n793), .B1(G329), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n758), .ZN(new_n796));
  INV_X1    g0596(.A(new_n776), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G322), .A2(new_n796), .B1(new_n797), .B2(G303), .ZN(new_n798));
  AND3_X1   g0598(.A1(new_n795), .A2(new_n404), .A3(new_n798), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n791), .B(new_n799), .C1(KEYINPUT107), .C2(new_n790), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n783), .B1(new_n785), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n224), .B1(G20), .B2(new_n321), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n802), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT102), .Z(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT103), .Z(new_n808));
  NOR2_X1   g0608(.A1(new_n691), .A2(new_n252), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n809), .B1(new_n222), .B2(new_n268), .C1(new_n250), .C2(new_n264), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n252), .A2(G355), .A3(new_n227), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n810), .B(new_n811), .C1(G116), .C2(new_n227), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n801), .A2(new_n802), .B1(new_n808), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n805), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n682), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n756), .B1(new_n754), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT108), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  AOI21_X1  g0618(.A(new_n388), .B1(new_n668), .B2(new_n669), .ZN(new_n819));
  AND3_X1   g0619(.A1(new_n623), .A2(new_n625), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(new_n386), .B2(new_n390), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n717), .A2(new_n718), .A3(new_n823), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n822), .B(new_n713), .C1(new_n646), .C2(new_n653), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n744), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n826), .A2(new_n744), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n827), .A2(new_n828), .A3(new_n754), .ZN(new_n829));
  INV_X1    g0629(.A(G283), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n404), .B1(new_n779), .B2(new_n784), .C1(new_n775), .C2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n774), .B1(G303), .B2(new_n761), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n789), .B2(new_n758), .ZN(new_n833));
  INV_X1    g0633(.A(new_n764), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n831), .B(new_n833), .C1(G116), .C2(new_n834), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n835), .B1(new_n210), .B2(new_n769), .C1(new_n240), .C2(new_n776), .ZN(new_n836));
  INV_X1    g0636(.A(new_n775), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G137), .A2(new_n761), .B1(new_n837), .B2(G150), .ZN(new_n838));
  INV_X1    g0638(.A(new_n759), .ZN(new_n839));
  INV_X1    g0639(.A(G143), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n838), .B1(new_n780), .B2(new_n764), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT34), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n252), .B1(new_n776), .B2(new_n202), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n769), .A2(new_n215), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n845), .B(new_n846), .C1(G58), .C2(new_n772), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n843), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G132), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n779), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n836), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n754), .B1(new_n851), .B2(new_n802), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n802), .A2(new_n803), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n208), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n852), .B(new_n854), .C1(new_n822), .C2(new_n804), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n829), .A2(new_n855), .ZN(G384));
  INV_X1    g0656(.A(KEYINPUT35), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n223), .B(new_n224), .C1(new_n463), .C2(new_n857), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n858), .B(G116), .C1(new_n857), .C2(new_n463), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT36), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n401), .A2(new_n222), .A3(new_n208), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT109), .Z(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(G50), .B2(new_n215), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(G1), .A3(new_n284), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT40), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n735), .A2(new_n722), .ZN(new_n866));
  INV_X1    g0666(.A(new_n721), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n737), .B1(new_n727), .B2(new_n734), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n343), .A2(new_n670), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n620), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n369), .A2(KEYINPUT110), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n361), .A2(G169), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT14), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n361), .A2(new_n345), .A3(G169), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(new_n366), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT77), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n364), .A2(new_n344), .A3(new_n366), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT110), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n880), .A3(new_n343), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n871), .B1(new_n872), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n369), .B1(new_n620), .B2(new_n870), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n822), .B(new_n869), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT37), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n416), .A2(new_n405), .A3(new_n406), .ZN(new_n887));
  INV_X1    g0687(.A(new_n412), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n423), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n889), .A2(KEYINPUT16), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n413), .A2(new_n312), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n400), .ZN(new_n893));
  INV_X1    g0693(.A(new_n665), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n892), .A2(new_n893), .B1(new_n447), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n886), .B1(new_n895), .B2(new_n441), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n665), .B(KEYINPUT111), .Z(new_n897));
  OAI21_X1  g0697(.A(new_n444), .B1(new_n447), .B2(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n898), .A2(new_n886), .A3(new_n441), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n890), .A2(new_n891), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n665), .B1(new_n901), .B2(new_n400), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n619), .B2(new_n635), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n885), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n450), .A2(new_n902), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n901), .A2(new_n400), .B1(new_n632), .B2(new_n665), .ZN(new_n907));
  INV_X1    g0707(.A(new_n441), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT37), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n898), .A2(new_n886), .A3(new_n441), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n906), .A2(new_n911), .A3(KEYINPUT38), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n905), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n865), .B1(new_n884), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n871), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n880), .B1(new_n879), .B2(new_n343), .ZN(new_n916));
  INV_X1    g0716(.A(new_n343), .ZN(new_n917));
  AOI211_X1 g0717(.A(KEYINPUT110), .B(new_n917), .C1(new_n877), .C2(new_n878), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n915), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n628), .A2(new_n871), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(KEYINPUT112), .B(KEYINPUT38), .Z(new_n922));
  INV_X1    g0722(.A(new_n897), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n426), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n619), .B2(new_n635), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n886), .B1(new_n898), .B2(new_n441), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n899), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n922), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n865), .B1(new_n929), .B2(new_n912), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n921), .A2(new_n930), .A3(new_n822), .A4(new_n869), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n914), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n455), .B1(new_n736), .B2(new_n868), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(G330), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n720), .A2(new_n455), .ZN(new_n936));
  INV_X1    g0736(.A(new_n638), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT39), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n906), .A2(new_n911), .A3(KEYINPUT38), .ZN(new_n940));
  INV_X1    g0740(.A(new_n922), .ZN(new_n941));
  INV_X1    g0741(.A(new_n927), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n910), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n450), .A2(new_n924), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n939), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n872), .A2(new_n713), .A3(new_n881), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n905), .A2(KEYINPUT39), .A3(new_n912), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n633), .A2(new_n634), .A3(new_n923), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n905), .A2(new_n912), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n386), .A2(new_n670), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n825), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n921), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n950), .A2(new_n951), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n938), .B(new_n957), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n935), .A2(new_n958), .B1(new_n263), .B2(new_n656), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT113), .Z(new_n960));
  AND2_X1   g0760(.A1(new_n935), .A2(new_n958), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n860), .B(new_n864), .C1(new_n960), .C2(new_n961), .ZN(G367));
  NOR2_X1   g0762(.A1(new_n713), .A2(new_n511), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT114), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(new_n639), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n701), .A2(new_n702), .B1(new_n470), .B2(new_n713), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n709), .A2(new_n670), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(new_n684), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT42), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n647), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n670), .B1(new_n973), .B2(new_n548), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n966), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n686), .A2(new_n970), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n980), .B1(new_n977), .B2(new_n978), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n679), .A2(new_n969), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT44), .Z(new_n984));
  NAND2_X1  g0784(.A1(new_n679), .A2(new_n969), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT45), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n686), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n685), .A2(new_n684), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n988), .B1(new_n748), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n746), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n746), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n692), .B(KEYINPUT41), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n981), .B(new_n982), .C1(new_n994), .C2(new_n752), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n758), .A2(new_n298), .B1(new_n776), .B2(new_n301), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n773), .A2(new_n215), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n252), .B1(new_n764), .B2(new_n202), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G159), .B2(new_n837), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n794), .A2(G137), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n768), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n761), .A2(G143), .B1(new_n1002), .B2(G77), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n773), .A2(new_n240), .B1(new_n768), .B2(new_n242), .ZN(new_n1005));
  INV_X1    g0805(.A(G317), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n404), .B1(new_n779), .B2(new_n1006), .C1(new_n830), .C2(new_n764), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1005), .B(new_n1007), .C1(G294), .C2(new_n837), .ZN(new_n1008));
  INV_X1    g0808(.A(G303), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1008), .B1(new_n1009), .B2(new_n839), .C1(new_n784), .C2(new_n787), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n776), .A2(new_n514), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT46), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1004), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT47), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n802), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n807), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n809), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1016), .B1(new_n227), .B2(new_n379), .C1(new_n237), .C2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1015), .A2(new_n753), .A3(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT115), .Z(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n814), .B2(new_n965), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n995), .A2(new_n1021), .ZN(G387));
  OR2_X1    g0822(.A1(new_n990), .A2(new_n746), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1023), .A2(new_n692), .A3(new_n991), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n404), .B1(new_n768), .B2(new_n514), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G322), .A2(new_n761), .B1(new_n837), .B2(G311), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n1009), .B2(new_n764), .C1(new_n839), .C2(new_n1006), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT48), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n830), .B2(new_n773), .C1(new_n789), .C2(new_n776), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT49), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1025), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n1030), .B2(new_n1029), .C1(new_n788), .C2(new_n779), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n252), .B1(new_n215), .B2(new_n764), .C1(new_n309), .C2(new_n775), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n776), .A2(new_n208), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n787), .A2(new_n780), .B1(new_n202), .B2(new_n758), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n773), .A2(new_n379), .ZN(new_n1036));
  NOR4_X1   g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n242), .B2(new_n769), .C1(new_n298), .C2(new_n779), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1032), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n754), .B1(new_n1039), .B2(new_n802), .ZN(new_n1040));
  OR3_X1    g0840(.A1(new_n378), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT50), .B1(new_n378), .B2(G50), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1041), .A2(new_n264), .A3(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1043), .B(new_n690), .C1(G68), .C2(G77), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n268), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n809), .B1(new_n234), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n690), .A2(new_n227), .A3(new_n252), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n227), .A2(G107), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n808), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1040), .B(new_n1050), .C1(new_n674), .C2(new_n814), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT116), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n990), .A2(new_n752), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1024), .A2(new_n1052), .A3(new_n1053), .ZN(G393));
  NOR2_X1   g0854(.A1(new_n987), .A2(new_n686), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n984), .A2(new_n988), .A3(new_n986), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n991), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1057), .B(new_n692), .C1(new_n991), .C2(new_n987), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1016), .B1(new_n242), .B2(new_n227), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n246), .B2(new_n809), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n787), .A2(new_n1006), .B1(new_n784), .B2(new_n758), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT52), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n404), .B1(new_n764), .B2(new_n789), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n773), .A2(new_n514), .B1(new_n776), .B2(new_n830), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(G322), .C2(new_n794), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1062), .B(new_n1065), .C1(new_n240), .C2(new_n769), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n775), .A2(new_n1009), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n776), .A2(new_n215), .B1(new_n779), .B2(new_n840), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT117), .Z(new_n1069));
  OAI22_X1  g0869(.A1(new_n769), .A2(new_n210), .B1(new_n208), .B2(new_n773), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n252), .B1(new_n764), .B2(new_n378), .C1(new_n202), .C2(new_n775), .ZN(new_n1071));
  OR3_X1    g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G150), .A2(new_n761), .B1(new_n796), .B2(G159), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT51), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n1066), .A2(new_n1067), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1060), .B1(new_n1075), .B2(new_n802), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n969), .B2(new_n814), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(new_n754), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1078), .B1(new_n1079), .B2(new_n752), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1058), .A2(new_n1080), .ZN(G390));
  NAND2_X1  g0881(.A1(new_n872), .A2(new_n881), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n883), .B1(new_n1082), .B2(new_n915), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n822), .A2(G330), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n869), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(KEYINPUT119), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT119), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1084), .B1(new_n736), .B2(new_n868), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n921), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n743), .A2(new_n1085), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n1083), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1087), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n954), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n712), .A2(new_n713), .A3(new_n822), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n953), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n921), .A2(new_n743), .A3(new_n1085), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1094), .A2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n392), .A2(G330), .A3(new_n454), .A4(new_n869), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n638), .B(new_n1102), .C1(new_n720), .C2(new_n455), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n954), .B1(new_n882), .B2(new_n883), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1106), .A2(new_n947), .B1(new_n946), .B2(new_n949), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1098), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT118), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1096), .A2(new_n921), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n929), .A2(new_n912), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n947), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1110), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1095), .A2(new_n953), .B1(new_n919), .B2(new_n920), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1116), .A2(KEYINPUT118), .A3(new_n1113), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1108), .B(new_n1109), .C1(new_n1115), .C2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1111), .A2(new_n1110), .A3(new_n1114), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT118), .B1(new_n1116), .B2(new_n1113), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1107), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1105), .B(new_n1118), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1103), .B1(new_n1094), .B2(new_n1100), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1098), .B(new_n1107), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1124), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1123), .A2(new_n692), .A3(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1118), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n946), .A2(new_n949), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n803), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n309), .A2(new_n853), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT54), .B(G143), .Z(new_n1133));
  AOI21_X1  g0933(.A(new_n404), .B1(new_n834), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(G125), .ZN(new_n1135));
  INV_X1    g0935(.A(G137), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1134), .B1(new_n1135), .B2(new_n779), .C1(new_n1136), .C2(new_n775), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n797), .A2(G150), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT53), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1002), .A2(G50), .B1(new_n772), .B2(G159), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n849), .B2(new_n758), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1137), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(G128), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1142), .B1(new_n1143), .B2(new_n787), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n846), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n775), .A2(new_n240), .B1(new_n779), .B2(new_n789), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(G97), .B2(new_n834), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n796), .A2(G116), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n761), .A2(G283), .B1(G77), .B2(new_n772), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n404), .B1(new_n776), .B2(new_n210), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT120), .Z(new_n1152));
  OAI21_X1  g0952(.A(new_n1144), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n754), .B1(new_n1153), .B2(new_n802), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1131), .A2(new_n1132), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT121), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1129), .A2(new_n752), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1128), .A2(new_n1159), .ZN(G378));
  NAND2_X1  g0960(.A1(new_n1127), .A2(new_n1104), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n914), .A2(G330), .A3(new_n931), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n324), .A2(KEYINPUT55), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT55), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n318), .A2(new_n1164), .A3(new_n320), .A4(new_n323), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n316), .A2(new_n665), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT56), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT122), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1163), .A2(new_n1165), .A3(new_n1168), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1162), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1175), .A2(new_n914), .A3(G330), .A4(new_n931), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n957), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT123), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n956), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1174), .A2(KEYINPUT123), .A3(new_n957), .A4(new_n1176), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1179), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT57), .B1(new_n1161), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1177), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n957), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT57), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1103), .B1(new_n1129), .B2(new_n1124), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n692), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1184), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1170), .A2(new_n803), .A3(new_n1172), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n853), .A2(new_n202), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n775), .A2(new_n242), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n764), .A2(new_n379), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n779), .A2(new_n830), .ZN(new_n1195));
  OR4_X1    g0995(.A1(G41), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  NOR4_X1   g0996(.A1(new_n1196), .A2(new_n252), .A3(new_n997), .A4(new_n1034), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G116), .A2(new_n761), .B1(new_n796), .B2(G107), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n301), .C2(new_n768), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT58), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n787), .A2(new_n1135), .B1(new_n1143), .B2(new_n758), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n837), .A2(G132), .B1(G150), .B2(new_n772), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n1136), .B2(new_n764), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(new_n797), .C2(new_n1133), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT59), .ZN(new_n1205));
  AOI21_X1  g1005(.A(G41), .B1(new_n1002), .B2(G159), .ZN(new_n1206));
  AOI21_X1  g1006(.A(G33), .B1(new_n794), .B2(G124), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1200), .B(new_n1208), .C1(G50), .C2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n754), .B1(new_n1210), .B2(new_n802), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1191), .A2(new_n1192), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1183), .B2(new_n752), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1190), .A2(new_n1214), .ZN(G375));
  OAI22_X1  g1015(.A1(new_n787), .A2(new_n849), .B1(new_n301), .B2(new_n768), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n404), .B1(new_n837), .B2(new_n1133), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n1143), .B2(new_n779), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n298), .B2(new_n764), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1216), .B(new_n1220), .C1(G50), .C2(new_n772), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n1136), .B2(new_n839), .C1(new_n780), .C2(new_n776), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n404), .B1(new_n779), .B2(new_n1009), .C1(new_n240), .C2(new_n764), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1036), .B1(G294), .B2(new_n761), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n242), .B2(new_n776), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(G116), .C2(new_n837), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n208), .B2(new_n769), .C1(new_n830), .C2(new_n758), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1222), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n754), .B1(new_n1228), .B2(new_n802), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n921), .B2(new_n804), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n215), .B2(new_n853), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1101), .B2(new_n752), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1094), .A2(new_n1103), .A3(new_n1100), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n993), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1232), .B1(new_n1234), .B2(new_n1124), .ZN(G381));
  NAND4_X1  g1035(.A1(new_n995), .A2(new_n1058), .A3(new_n1021), .A4(new_n1080), .ZN(new_n1236));
  OR2_X1    g1036(.A1(G381), .A2(G384), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(new_n1236), .A2(G396), .A3(G393), .A4(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(G378), .ZN(new_n1239));
  INV_X1    g1039(.A(G375), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(G407));
  NOR2_X1   g1041(.A1(new_n1238), .A2(new_n666), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1240), .A2(new_n1239), .ZN(new_n1243));
  OAI21_X1  g1043(.A(G213), .B1(new_n1242), .B2(new_n1243), .ZN(G409));
  NAND3_X1  g1044(.A1(new_n1161), .A2(new_n1183), .A3(new_n993), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n752), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1245), .A2(new_n1212), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1239), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G378), .B(new_n1214), .C1(new_n1184), .C2(new_n1189), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT124), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT60), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1233), .A2(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1094), .A2(KEYINPUT60), .A3(new_n1103), .A4(new_n1100), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1254), .A2(new_n1105), .A3(new_n692), .A4(new_n1255), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1256), .A2(G384), .A3(new_n1232), .ZN(new_n1257));
  AOI21_X1  g1057(.A(G384), .B1(new_n1256), .B2(new_n1232), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n666), .A2(G213), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1248), .A2(new_n1249), .A3(KEYINPUT124), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1252), .A2(new_n1259), .A3(new_n1260), .A4(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1262), .A2(KEYINPUT62), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1250), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT62), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT61), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1250), .A2(new_n1260), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n666), .A2(G213), .A3(G2897), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT125), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1097), .A2(new_n1271), .B1(new_n1093), .B2(new_n954), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1255), .B(new_n692), .C1(new_n1103), .C2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT60), .B1(new_n1272), .B2(new_n1103), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1232), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(G384), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT125), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1256), .A2(G384), .A3(new_n1232), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1269), .B1(new_n1270), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1268), .B1(new_n1259), .B2(new_n1278), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1267), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1265), .A2(new_n1266), .A3(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(KEYINPUT126), .B1(new_n1263), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G387), .A2(G390), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n817), .B(G393), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n1288), .A3(new_n1236), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1288), .B1(new_n1287), .B2(new_n1236), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1248), .A2(new_n1249), .A3(KEYINPUT124), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT124), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT62), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1295), .A2(new_n1296), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT126), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT61), .B1(new_n1264), .B2(KEYINPUT62), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1297), .A2(new_n1298), .A3(new_n1284), .A4(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1286), .A2(new_n1292), .A3(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1291), .ZN(new_n1302));
  AOI21_X1  g1102(.A(KEYINPUT61), .B1(new_n1302), .B2(new_n1289), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  OR2_X1    g1104(.A1(new_n1264), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1262), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1252), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1304), .B1(new_n1307), .B2(new_n1283), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1303), .B(new_n1305), .C1(new_n1306), .C2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1301), .A2(new_n1309), .ZN(G405));
  NAND2_X1  g1110(.A1(new_n1249), .A2(KEYINPUT127), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1311), .B(new_n1259), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(G375), .A2(new_n1239), .ZN(new_n1313));
  OR2_X1    g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1314), .A2(new_n1292), .A3(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1292), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(G402));
endmodule


