

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n618), .A2(n983), .ZN(n612) );
  NAND2_X2 U553 ( .A1(n586), .A2(n684), .ZN(n656) );
  XOR2_X2 U554 ( .A(n568), .B(KEYINPUT17), .Z(n691) );
  NAND2_X1 U555 ( .A1(n582), .A2(n581), .ZN(n758) );
  NOR2_X2 U556 ( .A1(n548), .A2(n522), .ZN(n518) );
  NOR2_X1 U557 ( .A1(n656), .A2(n947), .ZN(n588) );
  INV_X1 U558 ( .A(KEYINPUT84), .ZN(n611) );
  INV_X1 U559 ( .A(KEYINPUT29), .ZN(n637) );
  XNOR2_X1 U560 ( .A(n638), .B(n637), .ZN(n645) );
  NAND2_X1 U561 ( .A1(n674), .A2(n673), .ZN(n737) );
  NOR2_X1 U562 ( .A1(G651), .A2(n548), .ZN(n786) );
  XNOR2_X1 U563 ( .A(KEYINPUT40), .B(KEYINPUT95), .ZN(n754) );
  XOR2_X1 U564 ( .A(G543), .B(KEYINPUT0), .Z(n548) );
  NAND2_X1 U565 ( .A1(n786), .A2(G52), .ZN(n521) );
  XOR2_X1 U566 ( .A(KEYINPUT66), .B(G651), .Z(n522) );
  NOR2_X1 U567 ( .A1(G543), .A2(n522), .ZN(n519) );
  XOR2_X2 U568 ( .A(KEYINPUT1), .B(n519), .Z(n787) );
  NAND2_X1 U569 ( .A1(G64), .A2(n787), .ZN(n520) );
  NAND2_X1 U570 ( .A1(n521), .A2(n520), .ZN(n528) );
  NOR2_X1 U571 ( .A1(G651), .A2(G543), .ZN(n783) );
  NAND2_X1 U572 ( .A1(G90), .A2(n783), .ZN(n524) );
  NAND2_X1 U573 ( .A1(G77), .A2(n518), .ZN(n523) );
  NAND2_X1 U574 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U575 ( .A(KEYINPUT67), .B(n525), .ZN(n526) );
  XNOR2_X1 U576 ( .A(KEYINPUT9), .B(n526), .ZN(n527) );
  NOR2_X1 U577 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U578 ( .A(KEYINPUT68), .B(n529), .ZN(G171) );
  NAND2_X1 U579 ( .A1(n783), .A2(G89), .ZN(n530) );
  XNOR2_X1 U580 ( .A(n530), .B(KEYINPUT4), .ZN(n532) );
  NAND2_X1 U581 ( .A1(G76), .A2(n518), .ZN(n531) );
  NAND2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U583 ( .A(n533), .B(KEYINPUT5), .ZN(n538) );
  NAND2_X1 U584 ( .A1(n786), .A2(G51), .ZN(n535) );
  NAND2_X1 U585 ( .A1(G63), .A2(n787), .ZN(n534) );
  NAND2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U587 ( .A(KEYINPUT6), .B(n536), .Z(n537) );
  NAND2_X1 U588 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U589 ( .A(n539), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U590 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U591 ( .A1(G88), .A2(n783), .ZN(n541) );
  NAND2_X1 U592 ( .A1(G75), .A2(n518), .ZN(n540) );
  NAND2_X1 U593 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U594 ( .A(KEYINPUT75), .B(n542), .ZN(n547) );
  NAND2_X1 U595 ( .A1(n786), .A2(G50), .ZN(n544) );
  NAND2_X1 U596 ( .A1(G62), .A2(n787), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U598 ( .A(KEYINPUT74), .B(n545), .Z(n546) );
  NAND2_X1 U599 ( .A1(n547), .A2(n546), .ZN(G303) );
  NAND2_X1 U600 ( .A1(G87), .A2(n548), .ZN(n550) );
  NAND2_X1 U601 ( .A1(G74), .A2(G651), .ZN(n549) );
  NAND2_X1 U602 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U603 ( .A1(n787), .A2(n551), .ZN(n553) );
  NAND2_X1 U604 ( .A1(n786), .A2(G49), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n553), .A2(n552), .ZN(G288) );
  NAND2_X1 U606 ( .A1(G86), .A2(n783), .ZN(n555) );
  NAND2_X1 U607 ( .A1(G48), .A2(n786), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U609 ( .A1(n518), .A2(G73), .ZN(n556) );
  XNOR2_X1 U610 ( .A(n556), .B(KEYINPUT2), .ZN(n557) );
  XNOR2_X1 U611 ( .A(n557), .B(KEYINPUT73), .ZN(n558) );
  NOR2_X1 U612 ( .A1(n559), .A2(n558), .ZN(n561) );
  NAND2_X1 U613 ( .A1(G61), .A2(n787), .ZN(n560) );
  NAND2_X1 U614 ( .A1(n561), .A2(n560), .ZN(G305) );
  NAND2_X1 U615 ( .A1(G85), .A2(n783), .ZN(n563) );
  NAND2_X1 U616 ( .A1(G72), .A2(n518), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U618 ( .A1(n786), .A2(G47), .ZN(n565) );
  NAND2_X1 U619 ( .A1(G60), .A2(n787), .ZN(n564) );
  NAND2_X1 U620 ( .A1(n565), .A2(n564), .ZN(n566) );
  OR2_X1 U621 ( .A1(n567), .A2(n566), .ZN(G290) );
  NOR2_X1 U622 ( .A1(G2104), .A2(G2105), .ZN(n568) );
  NAND2_X1 U623 ( .A1(n691), .A2(G137), .ZN(n757) );
  INV_X1 U624 ( .A(G2105), .ZN(n571) );
  AND2_X1 U625 ( .A1(n571), .A2(G2104), .ZN(n578) );
  NAND2_X1 U626 ( .A1(n578), .A2(G101), .ZN(n569) );
  XNOR2_X1 U627 ( .A(KEYINPUT23), .B(n569), .ZN(n575) );
  NAND2_X1 U628 ( .A1(G2104), .A2(G2105), .ZN(n570) );
  XNOR2_X2 U629 ( .A(n570), .B(KEYINPUT65), .ZN(n875) );
  NAND2_X1 U630 ( .A1(G113), .A2(n875), .ZN(n573) );
  NOR2_X2 U631 ( .A1(n571), .A2(G2104), .ZN(n876) );
  NAND2_X1 U632 ( .A1(G125), .A2(n876), .ZN(n572) );
  NAND2_X1 U633 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U634 ( .A1(n575), .A2(n574), .ZN(n756) );
  AND2_X1 U635 ( .A1(n756), .A2(G40), .ZN(n576) );
  NAND2_X1 U636 ( .A1(n757), .A2(n576), .ZN(n685) );
  INV_X1 U637 ( .A(n685), .ZN(n586) );
  INV_X1 U638 ( .A(G1384), .ZN(n583) );
  AND2_X1 U639 ( .A1(G138), .A2(n583), .ZN(n577) );
  AND2_X1 U640 ( .A1(n691), .A2(n577), .ZN(n585) );
  NAND2_X1 U641 ( .A1(G126), .A2(n876), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G102), .A2(n578), .ZN(n579) );
  AND2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U644 ( .A1(n875), .A2(G114), .ZN(n581) );
  AND2_X1 U645 ( .A1(n583), .A2(n758), .ZN(n584) );
  OR2_X1 U646 ( .A1(n585), .A2(n584), .ZN(n684) );
  INV_X1 U647 ( .A(G1996), .ZN(n947) );
  XOR2_X1 U648 ( .A(KEYINPUT26), .B(KEYINPUT82), .Z(n587) );
  XNOR2_X1 U649 ( .A(n588), .B(n587), .ZN(n590) );
  NAND2_X1 U650 ( .A1(n656), .A2(G1341), .ZN(n589) );
  NAND2_X1 U651 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U652 ( .A(n591), .B(KEYINPUT83), .ZN(n602) );
  NAND2_X1 U653 ( .A1(n783), .A2(G81), .ZN(n592) );
  XNOR2_X1 U654 ( .A(KEYINPUT12), .B(n592), .ZN(n595) );
  NAND2_X1 U655 ( .A1(G68), .A2(n518), .ZN(n593) );
  XOR2_X1 U656 ( .A(KEYINPUT71), .B(n593), .Z(n594) );
  NAND2_X1 U657 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U658 ( .A(n596), .B(KEYINPUT13), .ZN(n598) );
  NAND2_X1 U659 ( .A1(G43), .A2(n786), .ZN(n597) );
  NAND2_X1 U660 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U661 ( .A1(n787), .A2(G56), .ZN(n599) );
  XOR2_X1 U662 ( .A(KEYINPUT14), .B(n599), .Z(n600) );
  NOR2_X2 U663 ( .A1(n601), .A2(n600), .ZN(n971) );
  NAND2_X1 U664 ( .A1(n602), .A2(n971), .ZN(n603) );
  XNOR2_X1 U665 ( .A(KEYINPUT64), .B(n603), .ZN(n618) );
  NAND2_X1 U666 ( .A1(n786), .A2(G54), .ZN(n605) );
  NAND2_X1 U667 ( .A1(G66), .A2(n787), .ZN(n604) );
  NAND2_X1 U668 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U669 ( .A1(G92), .A2(n783), .ZN(n607) );
  NAND2_X1 U670 ( .A1(G79), .A2(n518), .ZN(n606) );
  NAND2_X1 U671 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U672 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U673 ( .A(n610), .B(KEYINPUT15), .ZN(n983) );
  XNOR2_X1 U674 ( .A(n612), .B(n611), .ZN(n617) );
  NAND2_X1 U675 ( .A1(G1348), .A2(n656), .ZN(n614) );
  INV_X1 U676 ( .A(n656), .ZN(n639) );
  NAND2_X1 U677 ( .A1(n639), .A2(G2067), .ZN(n613) );
  NAND2_X1 U678 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U679 ( .A(KEYINPUT85), .B(n615), .Z(n616) );
  NAND2_X1 U680 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U681 ( .A1(n618), .A2(n983), .ZN(n619) );
  NAND2_X1 U682 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U683 ( .A(n621), .B(KEYINPUT86), .ZN(n632) );
  NAND2_X1 U684 ( .A1(n639), .A2(G2072), .ZN(n622) );
  XNOR2_X1 U685 ( .A(n622), .B(KEYINPUT27), .ZN(n624) );
  AND2_X1 U686 ( .A1(G1956), .A2(n656), .ZN(n623) );
  NOR2_X1 U687 ( .A1(n624), .A2(n623), .ZN(n633) );
  NAND2_X1 U688 ( .A1(n786), .A2(G53), .ZN(n626) );
  NAND2_X1 U689 ( .A1(G65), .A2(n787), .ZN(n625) );
  NAND2_X1 U690 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U691 ( .A1(G91), .A2(n783), .ZN(n628) );
  NAND2_X1 U692 ( .A1(G78), .A2(n518), .ZN(n627) );
  NAND2_X1 U693 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U694 ( .A1(n630), .A2(n629), .ZN(n972) );
  NAND2_X1 U695 ( .A1(n633), .A2(n972), .ZN(n631) );
  NAND2_X1 U696 ( .A1(n632), .A2(n631), .ZN(n636) );
  NOR2_X1 U697 ( .A1(n633), .A2(n972), .ZN(n634) );
  XOR2_X1 U698 ( .A(n634), .B(KEYINPUT28), .Z(n635) );
  NAND2_X1 U699 ( .A1(n636), .A2(n635), .ZN(n638) );
  NOR2_X1 U700 ( .A1(n639), .A2(G1961), .ZN(n640) );
  XNOR2_X1 U701 ( .A(n640), .B(KEYINPUT80), .ZN(n642) );
  XOR2_X1 U702 ( .A(G2078), .B(KEYINPUT25), .Z(n954) );
  NOR2_X1 U703 ( .A1(n656), .A2(n954), .ZN(n641) );
  NOR2_X1 U704 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U705 ( .A(KEYINPUT81), .B(n643), .ZN(n649) );
  NAND2_X1 U706 ( .A1(n649), .A2(G171), .ZN(n644) );
  NAND2_X1 U707 ( .A1(n645), .A2(n644), .ZN(n655) );
  NAND2_X1 U708 ( .A1(G8), .A2(n656), .ZN(n741) );
  NOR2_X1 U709 ( .A1(G1966), .A2(n741), .ZN(n670) );
  NOR2_X1 U710 ( .A1(G2084), .A2(n656), .ZN(n667) );
  NOR2_X1 U711 ( .A1(n670), .A2(n667), .ZN(n646) );
  NAND2_X1 U712 ( .A1(G8), .A2(n646), .ZN(n647) );
  XNOR2_X1 U713 ( .A(KEYINPUT30), .B(n647), .ZN(n648) );
  NOR2_X1 U714 ( .A1(G168), .A2(n648), .ZN(n651) );
  NOR2_X1 U715 ( .A1(n649), .A2(G171), .ZN(n650) );
  NOR2_X1 U716 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U717 ( .A(n652), .B(KEYINPUT87), .ZN(n653) );
  XNOR2_X1 U718 ( .A(n653), .B(KEYINPUT31), .ZN(n654) );
  NAND2_X1 U719 ( .A1(n655), .A2(n654), .ZN(n668) );
  NAND2_X1 U720 ( .A1(n668), .A2(G286), .ZN(n663) );
  NOR2_X1 U721 ( .A1(G2090), .A2(n656), .ZN(n657) );
  XNOR2_X1 U722 ( .A(n657), .B(KEYINPUT88), .ZN(n659) );
  NOR2_X1 U723 ( .A1(n741), .A2(G1971), .ZN(n658) );
  NOR2_X1 U724 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U725 ( .A(KEYINPUT89), .B(n660), .Z(n661) );
  NAND2_X1 U726 ( .A1(n661), .A2(G303), .ZN(n662) );
  NAND2_X1 U727 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U728 ( .A(n664), .B(KEYINPUT90), .ZN(n665) );
  NAND2_X1 U729 ( .A1(n665), .A2(G8), .ZN(n666) );
  XNOR2_X1 U730 ( .A(n666), .B(KEYINPUT32), .ZN(n674) );
  NAND2_X1 U731 ( .A1(G8), .A2(n667), .ZN(n672) );
  INV_X1 U732 ( .A(n668), .ZN(n669) );
  NOR2_X1 U733 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U734 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U735 ( .A1(G1976), .A2(G288), .ZN(n974) );
  NOR2_X1 U736 ( .A1(G1971), .A2(G303), .ZN(n675) );
  NOR2_X1 U737 ( .A1(n974), .A2(n675), .ZN(n676) );
  XOR2_X1 U738 ( .A(KEYINPUT91), .B(n676), .Z(n677) );
  NAND2_X1 U739 ( .A1(n737), .A2(n677), .ZN(n678) );
  XNOR2_X1 U740 ( .A(n678), .B(KEYINPUT92), .ZN(n719) );
  NAND2_X1 U741 ( .A1(G1976), .A2(G288), .ZN(n977) );
  INV_X1 U742 ( .A(n977), .ZN(n679) );
  NOR2_X1 U743 ( .A1(n741), .A2(n679), .ZN(n682) );
  NAND2_X1 U744 ( .A1(n974), .A2(KEYINPUT33), .ZN(n680) );
  NOR2_X1 U745 ( .A1(n680), .A2(n741), .ZN(n743) );
  INV_X1 U746 ( .A(n743), .ZN(n681) );
  AND2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U748 ( .A(G1981), .B(G305), .Z(n967) );
  AND2_X1 U749 ( .A1(n683), .A2(n967), .ZN(n717) );
  NOR2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n730) );
  XNOR2_X1 U751 ( .A(KEYINPUT78), .B(n730), .ZN(n703) );
  NAND2_X1 U752 ( .A1(G95), .A2(n578), .ZN(n687) );
  NAND2_X1 U753 ( .A1(G119), .A2(n876), .ZN(n686) );
  NAND2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n690) );
  NAND2_X1 U755 ( .A1(G107), .A2(n875), .ZN(n688) );
  XNOR2_X1 U756 ( .A(KEYINPUT77), .B(n688), .ZN(n689) );
  NOR2_X1 U757 ( .A1(n690), .A2(n689), .ZN(n693) );
  NAND2_X1 U758 ( .A1(n691), .A2(G131), .ZN(n692) );
  NAND2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n886) );
  NAND2_X1 U760 ( .A1(G1991), .A2(n886), .ZN(n702) );
  NAND2_X1 U761 ( .A1(G141), .A2(n691), .ZN(n695) );
  NAND2_X1 U762 ( .A1(G129), .A2(n876), .ZN(n694) );
  NAND2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n698) );
  NAND2_X1 U764 ( .A1(n578), .A2(G105), .ZN(n696) );
  XOR2_X1 U765 ( .A(KEYINPUT38), .B(n696), .Z(n697) );
  NOR2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n700) );
  NAND2_X1 U767 ( .A1(n875), .A2(G117), .ZN(n699) );
  NAND2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n859) );
  NAND2_X1 U769 ( .A1(G1996), .A2(n859), .ZN(n701) );
  NAND2_X1 U770 ( .A1(n702), .A2(n701), .ZN(n916) );
  NAND2_X1 U771 ( .A1(n703), .A2(n916), .ZN(n722) );
  NAND2_X1 U772 ( .A1(G104), .A2(n578), .ZN(n705) );
  NAND2_X1 U773 ( .A1(G140), .A2(n691), .ZN(n704) );
  NAND2_X1 U774 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U775 ( .A(KEYINPUT34), .B(n706), .ZN(n711) );
  NAND2_X1 U776 ( .A1(G116), .A2(n875), .ZN(n708) );
  NAND2_X1 U777 ( .A1(G128), .A2(n876), .ZN(n707) );
  NAND2_X1 U778 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U779 ( .A(KEYINPUT35), .B(n709), .Z(n710) );
  NOR2_X1 U780 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U781 ( .A(KEYINPUT36), .B(n712), .ZN(n872) );
  XNOR2_X1 U782 ( .A(G2067), .B(KEYINPUT37), .ZN(n728) );
  NOR2_X1 U783 ( .A1(n872), .A2(n728), .ZN(n929) );
  NAND2_X1 U784 ( .A1(n730), .A2(n929), .ZN(n727) );
  NAND2_X1 U785 ( .A1(n722), .A2(n727), .ZN(n713) );
  XNOR2_X1 U786 ( .A(n713), .B(KEYINPUT79), .ZN(n715) );
  XNOR2_X1 U787 ( .A(G1986), .B(G290), .ZN(n976) );
  NAND2_X1 U788 ( .A1(n730), .A2(n976), .ZN(n714) );
  NAND2_X1 U789 ( .A1(n715), .A2(n714), .ZN(n750) );
  INV_X1 U790 ( .A(n750), .ZN(n716) );
  AND2_X1 U791 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U792 ( .A1(n719), .A2(n718), .ZN(n734) );
  NOR2_X1 U793 ( .A1(G1986), .A2(G290), .ZN(n720) );
  NOR2_X1 U794 ( .A1(G1991), .A2(n886), .ZN(n918) );
  NOR2_X1 U795 ( .A1(n720), .A2(n918), .ZN(n721) );
  XNOR2_X1 U796 ( .A(n721), .B(KEYINPUT93), .ZN(n723) );
  NAND2_X1 U797 ( .A1(n723), .A2(n722), .ZN(n724) );
  OR2_X1 U798 ( .A1(n859), .A2(G1996), .ZN(n934) );
  NAND2_X1 U799 ( .A1(n724), .A2(n934), .ZN(n725) );
  XOR2_X1 U800 ( .A(KEYINPUT39), .B(n725), .Z(n726) );
  NAND2_X1 U801 ( .A1(n727), .A2(n726), .ZN(n729) );
  NAND2_X1 U802 ( .A1(n872), .A2(n728), .ZN(n927) );
  NAND2_X1 U803 ( .A1(n729), .A2(n927), .ZN(n731) );
  NAND2_X1 U804 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U805 ( .A(KEYINPUT94), .B(n732), .ZN(n733) );
  NAND2_X1 U806 ( .A1(n734), .A2(n733), .ZN(n753) );
  NOR2_X1 U807 ( .A1(G2090), .A2(G303), .ZN(n735) );
  NAND2_X1 U808 ( .A1(G8), .A2(n735), .ZN(n736) );
  NAND2_X1 U809 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U810 ( .A1(n738), .A2(n741), .ZN(n749) );
  NOR2_X1 U811 ( .A1(G1981), .A2(G305), .ZN(n739) );
  XOR2_X1 U812 ( .A(n739), .B(KEYINPUT24), .Z(n740) );
  OR2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n747) );
  INV_X1 U814 ( .A(n967), .ZN(n745) );
  INV_X1 U815 ( .A(KEYINPUT33), .ZN(n742) );
  OR2_X1 U816 ( .A1(n743), .A2(n742), .ZN(n744) );
  OR2_X1 U817 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U818 ( .A1(n747), .A2(n746), .ZN(n748) );
  AND2_X1 U819 ( .A1(n749), .A2(n748), .ZN(n751) );
  NOR2_X1 U820 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U821 ( .A1(n753), .A2(n752), .ZN(n755) );
  XNOR2_X1 U822 ( .A(n755), .B(n754), .ZN(G329) );
  AND2_X1 U823 ( .A1(n757), .A2(n756), .ZN(G160) );
  INV_X1 U824 ( .A(G57), .ZN(G237) );
  INV_X1 U825 ( .A(G132), .ZN(G219) );
  AND2_X1 U826 ( .A1(G138), .A2(n691), .ZN(n759) );
  NOR2_X1 U827 ( .A1(n759), .A2(n758), .ZN(G164) );
  NAND2_X1 U828 ( .A1(G94), .A2(G452), .ZN(n760) );
  XNOR2_X1 U829 ( .A(n760), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U830 ( .A1(G7), .A2(G661), .ZN(n761) );
  XNOR2_X1 U831 ( .A(n761), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U832 ( .A(G223), .ZN(n820) );
  NAND2_X1 U833 ( .A1(n820), .A2(G567), .ZN(n762) );
  XOR2_X1 U834 ( .A(KEYINPUT11), .B(n762), .Z(G234) );
  NAND2_X1 U835 ( .A1(n971), .A2(G860), .ZN(G153) );
  INV_X1 U836 ( .A(G171), .ZN(G301) );
  NAND2_X1 U837 ( .A1(G301), .A2(G868), .ZN(n764) );
  INV_X1 U838 ( .A(G868), .ZN(n804) );
  NAND2_X1 U839 ( .A1(n983), .A2(n804), .ZN(n763) );
  NAND2_X1 U840 ( .A1(n764), .A2(n763), .ZN(G284) );
  INV_X1 U841 ( .A(n972), .ZN(G299) );
  NOR2_X1 U842 ( .A1(G286), .A2(n804), .ZN(n766) );
  NOR2_X1 U843 ( .A1(G868), .A2(G299), .ZN(n765) );
  NOR2_X1 U844 ( .A1(n766), .A2(n765), .ZN(G297) );
  INV_X1 U845 ( .A(G860), .ZN(n767) );
  NAND2_X1 U846 ( .A1(n767), .A2(G559), .ZN(n768) );
  INV_X1 U847 ( .A(n983), .ZN(n792) );
  NAND2_X1 U848 ( .A1(n768), .A2(n792), .ZN(n769) );
  XNOR2_X1 U849 ( .A(n769), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U850 ( .A1(n792), .A2(G868), .ZN(n770) );
  NOR2_X1 U851 ( .A1(G559), .A2(n770), .ZN(n772) );
  AND2_X1 U852 ( .A1(n804), .A2(n971), .ZN(n771) );
  NOR2_X1 U853 ( .A1(n772), .A2(n771), .ZN(G282) );
  NAND2_X1 U854 ( .A1(G123), .A2(n876), .ZN(n773) );
  XNOR2_X1 U855 ( .A(n773), .B(KEYINPUT18), .ZN(n776) );
  NAND2_X1 U856 ( .A1(G135), .A2(n691), .ZN(n774) );
  XNOR2_X1 U857 ( .A(n774), .B(KEYINPUT72), .ZN(n775) );
  NAND2_X1 U858 ( .A1(n776), .A2(n775), .ZN(n780) );
  NAND2_X1 U859 ( .A1(G99), .A2(n578), .ZN(n778) );
  NAND2_X1 U860 ( .A1(G111), .A2(n875), .ZN(n777) );
  NAND2_X1 U861 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U862 ( .A1(n780), .A2(n779), .ZN(n917) );
  XNOR2_X1 U863 ( .A(n917), .B(G2096), .ZN(n782) );
  INV_X1 U864 ( .A(G2100), .ZN(n781) );
  NAND2_X1 U865 ( .A1(n782), .A2(n781), .ZN(G156) );
  NAND2_X1 U866 ( .A1(G93), .A2(n783), .ZN(n785) );
  NAND2_X1 U867 ( .A1(G80), .A2(n518), .ZN(n784) );
  NAND2_X1 U868 ( .A1(n785), .A2(n784), .ZN(n791) );
  NAND2_X1 U869 ( .A1(n786), .A2(G55), .ZN(n789) );
  NAND2_X1 U870 ( .A1(G67), .A2(n787), .ZN(n788) );
  NAND2_X1 U871 ( .A1(n789), .A2(n788), .ZN(n790) );
  OR2_X1 U872 ( .A1(n791), .A2(n790), .ZN(n803) );
  NAND2_X1 U873 ( .A1(n792), .A2(G559), .ZN(n801) );
  XOR2_X1 U874 ( .A(n971), .B(n801), .Z(n793) );
  NOR2_X1 U875 ( .A1(G860), .A2(n793), .ZN(n794) );
  XOR2_X1 U876 ( .A(n803), .B(n794), .Z(G145) );
  INV_X1 U877 ( .A(G303), .ZN(G166) );
  XOR2_X1 U878 ( .A(n803), .B(G290), .Z(n799) );
  XNOR2_X1 U879 ( .A(n972), .B(G166), .ZN(n797) );
  XOR2_X1 U880 ( .A(KEYINPUT19), .B(G305), .Z(n795) );
  XNOR2_X1 U881 ( .A(G288), .B(n795), .ZN(n796) );
  XNOR2_X1 U882 ( .A(n797), .B(n796), .ZN(n798) );
  XNOR2_X1 U883 ( .A(n799), .B(n798), .ZN(n800) );
  XNOR2_X1 U884 ( .A(n971), .B(n800), .ZN(n892) );
  XNOR2_X1 U885 ( .A(n801), .B(n892), .ZN(n802) );
  NAND2_X1 U886 ( .A1(n802), .A2(G868), .ZN(n806) );
  NAND2_X1 U887 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U888 ( .A1(n806), .A2(n805), .ZN(G295) );
  NAND2_X1 U889 ( .A1(G2078), .A2(G2084), .ZN(n807) );
  XOR2_X1 U890 ( .A(KEYINPUT20), .B(n807), .Z(n808) );
  NAND2_X1 U891 ( .A1(G2090), .A2(n808), .ZN(n810) );
  XNOR2_X1 U892 ( .A(KEYINPUT21), .B(KEYINPUT76), .ZN(n809) );
  XNOR2_X1 U893 ( .A(n810), .B(n809), .ZN(n811) );
  NAND2_X1 U894 ( .A1(G2072), .A2(n811), .ZN(G158) );
  XNOR2_X1 U895 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U896 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NOR2_X1 U897 ( .A1(G220), .A2(G219), .ZN(n812) );
  XOR2_X1 U898 ( .A(KEYINPUT22), .B(n812), .Z(n813) );
  NOR2_X1 U899 ( .A1(G218), .A2(n813), .ZN(n814) );
  NAND2_X1 U900 ( .A1(G96), .A2(n814), .ZN(n826) );
  NAND2_X1 U901 ( .A1(n826), .A2(G2106), .ZN(n818) );
  NAND2_X1 U902 ( .A1(G69), .A2(G120), .ZN(n815) );
  NOR2_X1 U903 ( .A1(G237), .A2(n815), .ZN(n816) );
  NAND2_X1 U904 ( .A1(G108), .A2(n816), .ZN(n827) );
  NAND2_X1 U905 ( .A1(n827), .A2(G567), .ZN(n817) );
  NAND2_X1 U906 ( .A1(n818), .A2(n817), .ZN(n828) );
  NAND2_X1 U907 ( .A1(G483), .A2(G661), .ZN(n819) );
  NOR2_X1 U908 ( .A1(n828), .A2(n819), .ZN(n825) );
  NAND2_X1 U909 ( .A1(n825), .A2(G36), .ZN(G176) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n820), .ZN(G217) );
  NAND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n821) );
  XOR2_X1 U912 ( .A(KEYINPUT100), .B(n821), .Z(n822) );
  NAND2_X1 U913 ( .A1(n822), .A2(G661), .ZN(n823) );
  XOR2_X1 U914 ( .A(KEYINPUT101), .B(n823), .Z(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n825), .A2(n824), .ZN(G188) );
  INV_X1 U918 ( .A(G120), .ZN(G236) );
  INV_X1 U919 ( .A(G96), .ZN(G221) );
  INV_X1 U920 ( .A(G69), .ZN(G235) );
  NOR2_X1 U921 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U922 ( .A(G325), .ZN(G261) );
  INV_X1 U923 ( .A(n828), .ZN(G319) );
  XNOR2_X1 U924 ( .A(G1981), .B(KEYINPUT41), .ZN(n838) );
  XOR2_X1 U925 ( .A(G1986), .B(G1971), .Z(n830) );
  XNOR2_X1 U926 ( .A(G1966), .B(G1961), .ZN(n829) );
  XNOR2_X1 U927 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U928 ( .A(G1991), .B(G1976), .Z(n832) );
  XNOR2_X1 U929 ( .A(G1956), .B(G1996), .ZN(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U931 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U932 ( .A(KEYINPUT104), .B(G2474), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U934 ( .A(n838), .B(n837), .ZN(G229) );
  XOR2_X1 U935 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n840) );
  XNOR2_X1 U936 ( .A(G2678), .B(KEYINPUT43), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U938 ( .A(KEYINPUT42), .B(G2090), .Z(n842) );
  XNOR2_X1 U939 ( .A(G2072), .B(G2067), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U941 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U942 ( .A(G2096), .B(G2100), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n848) );
  XOR2_X1 U944 ( .A(G2078), .B(G2084), .Z(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(G227) );
  NAND2_X1 U946 ( .A1(G124), .A2(n876), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n849), .B(KEYINPUT44), .ZN(n851) );
  NAND2_X1 U948 ( .A1(n875), .A2(G112), .ZN(n850) );
  NAND2_X1 U949 ( .A1(n851), .A2(n850), .ZN(n855) );
  NAND2_X1 U950 ( .A1(G100), .A2(n578), .ZN(n853) );
  NAND2_X1 U951 ( .A1(G136), .A2(n691), .ZN(n852) );
  NAND2_X1 U952 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U953 ( .A1(n855), .A2(n854), .ZN(G162) );
  XOR2_X1 U954 ( .A(KEYINPUT48), .B(KEYINPUT110), .Z(n857) );
  XNOR2_X1 U955 ( .A(KEYINPUT46), .B(KEYINPUT109), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U957 ( .A(n858), .B(G162), .Z(n861) );
  XOR2_X1 U958 ( .A(G160), .B(n859), .Z(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U960 ( .A(n917), .B(n862), .ZN(n874) );
  NAND2_X1 U961 ( .A1(n578), .A2(G103), .ZN(n863) );
  XNOR2_X1 U962 ( .A(KEYINPUT107), .B(n863), .ZN(n871) );
  NAND2_X1 U963 ( .A1(G115), .A2(n875), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G127), .A2(n876), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n866), .B(KEYINPUT47), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n867), .B(KEYINPUT108), .ZN(n869) );
  NAND2_X1 U968 ( .A1(n691), .A2(G139), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U970 ( .A1(n871), .A2(n870), .ZN(n922) );
  XNOR2_X1 U971 ( .A(n872), .B(n922), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(n890) );
  NAND2_X1 U973 ( .A1(G118), .A2(n875), .ZN(n878) );
  NAND2_X1 U974 ( .A1(G130), .A2(n876), .ZN(n877) );
  NAND2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n885) );
  XNOR2_X1 U976 ( .A(KEYINPUT45), .B(KEYINPUT106), .ZN(n883) );
  NAND2_X1 U977 ( .A1(n691), .A2(G142), .ZN(n881) );
  NAND2_X1 U978 ( .A1(n578), .A2(G106), .ZN(n879) );
  XOR2_X1 U979 ( .A(KEYINPUT105), .B(n879), .Z(n880) );
  NAND2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U981 ( .A(n883), .B(n882), .Z(n884) );
  NOR2_X1 U982 ( .A1(n885), .A2(n884), .ZN(n887) );
  XNOR2_X1 U983 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U984 ( .A(G164), .B(n888), .ZN(n889) );
  XNOR2_X1 U985 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U986 ( .A1(G37), .A2(n891), .ZN(G395) );
  XNOR2_X1 U987 ( .A(G286), .B(n983), .ZN(n893) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n894), .B(G171), .ZN(n895) );
  NOR2_X1 U990 ( .A1(G37), .A2(n895), .ZN(G397) );
  XOR2_X1 U991 ( .A(KEYINPUT96), .B(G2443), .Z(n897) );
  XNOR2_X1 U992 ( .A(G1341), .B(G1348), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n907) );
  XOR2_X1 U994 ( .A(G2427), .B(G2435), .Z(n899) );
  XNOR2_X1 U995 ( .A(G2430), .B(G2438), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n903) );
  XOR2_X1 U997 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n901) );
  XNOR2_X1 U998 ( .A(G2446), .B(G2454), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1000 ( .A(n903), .B(n902), .Z(n905) );
  XNOR2_X1 U1001 ( .A(G2451), .B(KEYINPUT97), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n908) );
  NAND2_X1 U1004 ( .A1(n908), .A2(G14), .ZN(n914) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n914), .ZN(n911) );
  NOR2_X1 U1006 ( .A1(G229), .A2(G227), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  INV_X1 U1013 ( .A(n914), .ZN(G401) );
  XOR2_X1 U1014 ( .A(G160), .B(G2084), .Z(n915) );
  NOR2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1017 ( .A(KEYINPUT111), .B(n919), .Z(n920) );
  NAND2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n933) );
  XOR2_X1 U1019 ( .A(G2072), .B(n922), .Z(n924) );
  XOR2_X1 U1020 ( .A(G164), .B(G2078), .Z(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(KEYINPUT112), .B(n925), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(n926), .B(KEYINPUT50), .ZN(n931) );
  INV_X1 U1024 ( .A(n927), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n938) );
  XNOR2_X1 U1028 ( .A(G2090), .B(G162), .ZN(n935) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1030 ( .A(n936), .B(KEYINPUT51), .ZN(n937) );
  NAND2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(n939), .B(KEYINPUT52), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(KEYINPUT113), .B(n940), .ZN(n941) );
  INV_X1 U1034 ( .A(KEYINPUT55), .ZN(n963) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n963), .ZN(n942) );
  NAND2_X1 U1036 ( .A1(n942), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1037 ( .A(KEYINPUT54), .B(KEYINPUT115), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(n943), .B(G34), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(G2084), .B(n944), .ZN(n961) );
  XNOR2_X1 U1040 ( .A(G2090), .B(G35), .ZN(n959) );
  XNOR2_X1 U1041 ( .A(G2072), .B(G33), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(G1991), .B(G25), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n953) );
  XNOR2_X1 U1044 ( .A(G32), .B(n947), .ZN(n948) );
  NAND2_X1 U1045 ( .A1(n948), .A2(G28), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(KEYINPUT114), .B(G2067), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(G26), .B(n949), .ZN(n950) );
  NOR2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(G27), .B(n954), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(KEYINPUT53), .B(n957), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(n963), .B(n962), .ZN(n965) );
  INV_X1 U1056 ( .A(G29), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1058 ( .A1(G11), .A2(n966), .ZN(n1028) );
  XNOR2_X1 U1059 ( .A(G16), .B(KEYINPUT56), .ZN(n994) );
  XNOR2_X1 U1060 ( .A(G1966), .B(G168), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(n969), .B(KEYINPUT57), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(KEYINPUT116), .B(n970), .ZN(n992) );
  XOR2_X1 U1064 ( .A(n971), .B(G1341), .Z(n990) );
  XNOR2_X1 U1065 ( .A(G1961), .B(G171), .ZN(n982) );
  XNOR2_X1 U1066 ( .A(n972), .B(G1956), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(n973), .B(KEYINPUT117), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(KEYINPUT118), .B(n974), .ZN(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n978) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n987) );
  XOR2_X1 U1073 ( .A(n983), .B(G1348), .Z(n985) );
  XNOR2_X1 U1074 ( .A(G166), .B(G1971), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(KEYINPUT119), .B(n988), .ZN(n989) );
  NOR2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n1026) );
  INV_X1 U1081 ( .A(G16), .ZN(n1024) );
  XOR2_X1 U1082 ( .A(G1961), .B(KEYINPUT120), .Z(n995) );
  XNOR2_X1 U1083 ( .A(G5), .B(n995), .ZN(n1020) );
  XOR2_X1 U1084 ( .A(G1976), .B(KEYINPUT125), .Z(n996) );
  XNOR2_X1 U1085 ( .A(G23), .B(n996), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G22), .B(G1971), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1088 ( .A(KEYINPUT126), .B(n999), .Z(n1001) );
  XNOR2_X1 U1089 ( .A(G1986), .B(G24), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(KEYINPUT58), .B(n1002), .ZN(n1015) );
  XNOR2_X1 U1092 ( .A(KEYINPUT59), .B(G1348), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(n1003), .B(G4), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(G1956), .B(G20), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(G1341), .B(G19), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(G1981), .B(G6), .ZN(n1004) );
  NOR2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1098 ( .A(KEYINPUT121), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n1011) );
  XNOR2_X1 U1102 ( .A(n1011), .B(KEYINPUT60), .ZN(n1012) );
  XNOR2_X1 U1103 ( .A(n1013), .B(n1012), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT124), .B(G1966), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(G21), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1109 ( .A(n1021), .B(KEYINPUT127), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

