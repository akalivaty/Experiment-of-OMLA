//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1275, new_n1276, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT1), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n209), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT0), .Z(new_n219));
  AND3_X1   g0019(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n220));
  AOI21_X1  g0020(.A(KEYINPUT65), .B1(G1), .B2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n201), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n216), .B(new_n219), .C1(new_n224), .C2(new_n227), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G58), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  AOI21_X1  g0045(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT68), .B(G1698), .ZN(new_n248));
  AND2_X1   g0048(.A1(new_n248), .A2(G222), .ZN(new_n249));
  INV_X1    g0049(.A(G223), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n247), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI221_X1 g0052(.A(new_n246), .B1(G77), .B2(new_n247), .C1(new_n249), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n255), .A2(G274), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(G226), .A2(new_n259), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n253), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G179), .ZN(new_n266));
  XOR2_X1   g0066(.A(new_n266), .B(KEYINPUT73), .Z(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT8), .B(G58), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT70), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G58), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(KEYINPUT70), .A3(KEYINPUT8), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n223), .A2(G33), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n269), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT69), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n280), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n222), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n223), .A2(G1), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n288), .B(KEYINPUT71), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n287), .A2(G50), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n286), .A2(new_n202), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n290), .A2(KEYINPUT72), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT72), .B1(new_n290), .B2(new_n291), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n284), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G169), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n265), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n267), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G20), .A2(G77), .ZN(new_n299));
  INV_X1    g0099(.A(new_n268), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT15), .B(G87), .ZN(new_n301));
  OAI221_X1 g0101(.A(new_n299), .B1(new_n270), .B2(new_n300), .C1(new_n276), .C2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G77), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n302), .A2(new_n283), .B1(new_n303), .B2(new_n286), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n287), .A2(G77), .A3(new_n289), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n263), .A2(new_n255), .A3(G274), .ZN(new_n307));
  INV_X1    g0107(.A(G244), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(new_n258), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT3), .ZN(new_n310));
  INV_X1    g0110(.A(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n251), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G238), .ZN(new_n315));
  INV_X1    g0115(.A(G107), .ZN(new_n316));
  INV_X1    g0116(.A(G232), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n251), .A2(KEYINPUT68), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT68), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G1698), .ZN(new_n320));
  AND2_X1   g0120(.A1(KEYINPUT3), .A2(G33), .ZN(new_n321));
  NOR2_X1   g0121(.A1(KEYINPUT3), .A2(G33), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n318), .B(new_n320), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  OAI221_X1 g0123(.A(new_n315), .B1(new_n316), .B2(new_n247), .C1(new_n317), .C2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n309), .B1(new_n324), .B2(new_n246), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n306), .B1(new_n325), .B2(G190), .ZN(new_n326));
  INV_X1    g0126(.A(G200), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n326), .B1(new_n327), .B2(new_n325), .ZN(new_n328));
  INV_X1    g0128(.A(G179), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n330), .B(new_n306), .C1(G169), .C2(new_n325), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n298), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(KEYINPUT9), .B(new_n284), .C1(new_n292), .C2(new_n293), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n253), .A2(G190), .A3(new_n264), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n335), .A2(KEYINPUT74), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n335), .A2(KEYINPUT74), .B1(new_n265), .B2(G200), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT9), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n294), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n338), .A2(KEYINPUT75), .A3(KEYINPUT10), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n342));
  OR2_X1    g0142(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n343));
  INV_X1    g0143(.A(new_n340), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n342), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G68), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n268), .A2(G50), .B1(G20), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n303), .B2(new_n276), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n283), .A2(new_n351), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n352), .A2(KEYINPUT11), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n286), .A2(new_n349), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT12), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n352), .A2(KEYINPUT11), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n287), .A2(G68), .A3(new_n289), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n353), .A2(new_n355), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT14), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n321), .A2(new_n322), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n318), .A2(new_n320), .A3(G226), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G232), .A2(G1698), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G97), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n246), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT13), .ZN(new_n367));
  AOI22_X1  g0167(.A1(G238), .A2(new_n259), .B1(new_n260), .B2(new_n263), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n367), .B1(new_n366), .B2(new_n368), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n359), .B(G169), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n371), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n369), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n372), .B1(new_n374), .B2(new_n329), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n359), .B1(new_n374), .B2(G169), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n358), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n370), .A2(new_n371), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n358), .B1(new_n378), .B2(G190), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT76), .ZN(new_n380));
  OAI21_X1  g0180(.A(G200), .B1(new_n370), .B2(new_n371), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n380), .B1(new_n379), .B2(new_n381), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n377), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AND3_X1   g0185(.A1(new_n289), .A2(new_n274), .A3(new_n272), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(new_n287), .B1(new_n275), .B2(new_n286), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n312), .A2(new_n223), .A3(new_n313), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT77), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n312), .A2(KEYINPUT7), .A3(new_n223), .A4(new_n313), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n392), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT77), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(G68), .A3(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n273), .A2(new_n349), .ZN(new_n397));
  OAI21_X1  g0197(.A(G20), .B1(new_n397), .B2(new_n201), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n268), .A2(G159), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT16), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT7), .B1(new_n360), .B2(new_n223), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n403), .B2(new_n394), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(KEYINPUT16), .A3(new_n401), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n283), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n387), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  OAI211_X1 g0207(.A(G226), .B(G1698), .C1(new_n321), .C2(new_n322), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G87), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n408), .B(new_n409), .C1(new_n323), .C2(new_n250), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n246), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n307), .B1(new_n317), .B2(new_n258), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n411), .A2(new_n413), .A3(G179), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n295), .B1(new_n411), .B2(new_n413), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n407), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT18), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n386), .A2(new_n287), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n275), .A2(new_n286), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n396), .A2(new_n401), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT16), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n283), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n390), .A2(new_n392), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n400), .B1(new_n426), .B2(G68), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n425), .B1(new_n427), .B2(KEYINPUT16), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n421), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n412), .B1(new_n246), .B2(new_n410), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT79), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT78), .B(G190), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n411), .A2(new_n413), .A3(new_n432), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n434), .B(KEYINPUT79), .C1(G200), .C2(new_n430), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n429), .A2(KEYINPUT17), .A3(new_n433), .A4(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n434), .A2(KEYINPUT79), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n430), .A2(G200), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n433), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n437), .B1(new_n440), .B2(new_n407), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT18), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n407), .A2(new_n416), .A3(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n418), .A2(new_n436), .A3(new_n441), .A4(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n333), .A2(new_n348), .A3(new_n385), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n286), .A2(new_n316), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n448), .B(KEYINPUT25), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n256), .A2(G33), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n282), .A2(new_n222), .A3(new_n285), .A4(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(new_n316), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n247), .A2(new_n223), .A3(G87), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT22), .ZN(new_n456));
  AOI21_X1  g0256(.A(G20), .B1(new_n312), .B2(new_n313), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT22), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n458), .A3(G87), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G116), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G20), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT23), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n223), .B2(G107), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n316), .A2(KEYINPUT23), .A3(G20), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT24), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT24), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n460), .A2(new_n469), .A3(new_n466), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n454), .B1(new_n471), .B2(new_n283), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT90), .ZN(new_n473));
  INV_X1    g0273(.A(G250), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n323), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g0275(.A1(KEYINPUT88), .A2(G294), .ZN(new_n476));
  NOR2_X1   g0276(.A1(KEYINPUT88), .A2(G294), .ZN(new_n477));
  OAI21_X1  g0277(.A(G33), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G257), .A2(G1698), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n478), .B1(new_n360), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(KEYINPUT89), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n248), .A2(new_n247), .A3(G250), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT89), .ZN(new_n483));
  INV_X1    g0283(.A(new_n479), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n247), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n482), .A2(new_n483), .A3(new_n478), .A4(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n481), .A2(new_n246), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n255), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n256), .A2(G45), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT5), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(G41), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT81), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n492), .B1(new_n261), .B2(KEYINPUT5), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n488), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT81), .B1(new_n490), .B2(G41), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(new_n491), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n262), .A2(G1), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n495), .B2(KEYINPUT81), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(G264), .A2(new_n497), .B1(new_n502), .B2(new_n260), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n295), .B1(new_n487), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n497), .A2(G264), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(new_n260), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n486), .A2(new_n246), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n481), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n473), .A2(new_n504), .B1(new_n509), .B2(G179), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT90), .B1(new_n509), .B2(new_n295), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n472), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n466), .ZN(new_n513));
  AOI211_X1 g0313(.A(KEYINPUT24), .B(new_n513), .C1(new_n456), .C2(new_n459), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n469), .B1(new_n460), .B2(new_n466), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n283), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(G190), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n486), .A2(new_n246), .ZN(new_n518));
  XNOR2_X1  g0318(.A(KEYINPUT88), .B(G294), .ZN(new_n519));
  AOI22_X1  g0319(.A1(G33), .A2(new_n519), .B1(new_n247), .B2(new_n484), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n483), .B1(new_n520), .B2(new_n482), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n503), .B(new_n517), .C1(new_n518), .C2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(G200), .B1(new_n487), .B2(new_n503), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n516), .B(new_n453), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n512), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n285), .A2(G116), .ZN(new_n528));
  INV_X1    g0328(.A(new_n451), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(G116), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n223), .A2(G116), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n282), .B2(new_n222), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G283), .ZN(new_n533));
  INV_X1    g0333(.A(G97), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n223), .C1(G33), .C2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT87), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n311), .A2(G97), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n538), .A2(KEYINPUT87), .A3(new_n223), .A4(new_n533), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT20), .B1(new_n532), .B2(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n532), .A2(KEYINPUT20), .A3(new_n540), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n530), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n432), .ZN(new_n544));
  OAI211_X1 g0344(.A(G270), .B(new_n255), .C1(new_n499), .C2(new_n501), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n506), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G303), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT86), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT86), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G303), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n314), .A2(G264), .B1(new_n551), .B2(new_n360), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT85), .ZN(new_n553));
  INV_X1    g0353(.A(G257), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n323), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n248), .A2(new_n247), .A3(KEYINPUT85), .A4(G257), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n552), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n546), .B1(new_n246), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n543), .B1(new_n544), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n327), .B2(new_n558), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(new_n246), .ZN(new_n561));
  AOI22_X1  g0361(.A1(G270), .A2(new_n497), .B1(new_n502), .B2(new_n260), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n543), .A2(new_n563), .A3(KEYINPUT21), .A4(G169), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n543), .A2(new_n558), .A3(G179), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n543), .A2(new_n563), .A3(G169), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT21), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n560), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n248), .A2(new_n247), .A3(KEYINPUT4), .A4(G244), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n314), .A2(G250), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n572), .A3(new_n533), .ZN(new_n573));
  INV_X1    g0373(.A(new_n323), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT4), .B1(new_n574), .B2(G244), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n246), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(G257), .A2(new_n497), .B1(new_n502), .B2(new_n260), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n295), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n329), .A3(new_n577), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n300), .A2(new_n303), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT6), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n583), .A2(new_n534), .A3(G107), .ZN(new_n584));
  XNOR2_X1  g0384(.A(G97), .B(G107), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n584), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(KEYINPUT80), .B(new_n582), .C1(new_n586), .C2(new_n223), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT80), .ZN(new_n588));
  AND2_X1   g0388(.A1(G97), .A2(G107), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n583), .B1(new_n589), .B2(new_n205), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n316), .A2(KEYINPUT6), .A3(G97), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n223), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n588), .B1(new_n592), .B2(new_n581), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n393), .A2(G107), .A3(new_n395), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n425), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n286), .A2(new_n534), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n451), .B2(new_n534), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n579), .B(new_n580), .C1(new_n596), .C2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n578), .A2(G200), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n595), .A2(new_n593), .A3(new_n587), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n598), .B1(new_n601), .B2(new_n283), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n576), .A2(G190), .A3(new_n577), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT84), .ZN(new_n606));
  OAI211_X1 g0406(.A(G244), .B(G1698), .C1(new_n321), .C2(new_n322), .ZN(new_n607));
  INV_X1    g0407(.A(G238), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n461), .B(new_n607), .C1(new_n323), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n246), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n255), .A2(G274), .A3(new_n500), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n255), .A2(G250), .A3(new_n489), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  AND4_X1   g0414(.A1(new_n606), .A2(new_n610), .A3(G190), .A4(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n613), .B1(new_n609), .B2(new_n246), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n606), .B1(new_n616), .B2(G190), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n610), .A2(new_n614), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G200), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT19), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT82), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT82), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT19), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n364), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT83), .B1(new_n625), .B2(G20), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n206), .A2(G87), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT83), .ZN(new_n629));
  XNOR2_X1  g0429(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n629), .B(new_n223), .C1(new_n630), .C2(new_n364), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n626), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n457), .A2(G68), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n630), .B1(new_n534), .B2(new_n276), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n425), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n301), .A2(new_n286), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(G87), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n451), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n636), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n618), .A2(new_n620), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n301), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n529), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n633), .A2(new_n634), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n622), .A2(new_n624), .ZN(new_n646));
  AOI21_X1  g0446(.A(G20), .B1(new_n646), .B2(new_n365), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n627), .B1(new_n647), .B2(new_n629), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n645), .B1(new_n648), .B2(new_n626), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n637), .B(new_n644), .C1(new_n649), .C2(new_n425), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n616), .A2(new_n329), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n650), .B(new_n651), .C1(G169), .C2(new_n616), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n642), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n605), .A2(new_n653), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n447), .A2(new_n527), .A3(new_n570), .A4(new_n654), .ZN(G372));
  AND3_X1   g0455(.A1(new_n341), .A2(new_n346), .A3(KEYINPUT95), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT95), .B1(new_n341), .B2(new_n346), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n382), .A2(new_n383), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n377), .B1(new_n659), .B2(new_n331), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(new_n441), .A3(new_n436), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n418), .A2(new_n443), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n658), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(new_n298), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT26), .B1(new_n653), .B2(new_n599), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n613), .A2(KEYINPUT91), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT91), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n611), .A2(new_n612), .A3(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n610), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n295), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n650), .A2(new_n651), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n579), .A2(new_n580), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n602), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT92), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n667), .A2(new_n669), .B1(new_n609), .B2(new_n246), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n677), .B1(new_n678), .B2(new_n327), .ZN(new_n679));
  OAI211_X1 g0479(.A(KEYINPUT92), .B(G200), .C1(new_n670), .C2(new_n671), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n618), .A2(new_n641), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n675), .A2(new_n676), .A3(new_n673), .A4(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n666), .A2(new_n673), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n569), .A2(new_n565), .A3(new_n564), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT93), .B1(new_n512), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n681), .A2(new_n525), .A3(new_n673), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n605), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n516), .A2(new_n453), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n503), .B1(new_n518), .B2(new_n521), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n689), .A2(new_n473), .A3(G169), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n487), .A2(G179), .A3(new_n503), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n504), .A2(new_n473), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n688), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT93), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(new_n566), .A4(new_n569), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n685), .A2(new_n687), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT94), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n685), .A2(new_n687), .A3(KEYINPUT94), .A4(new_n696), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n683), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n665), .B1(new_n446), .B2(new_n701), .ZN(G369));
  INV_X1    g0502(.A(new_n570), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n256), .A2(new_n223), .A3(G13), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G213), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G343), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n543), .A2(new_n709), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n684), .A2(new_n710), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G330), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n709), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n527), .B1(new_n472), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n694), .B2(new_n717), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n512), .A2(new_n717), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n684), .A2(new_n717), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n527), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n720), .A2(new_n721), .A3(new_n724), .ZN(G399));
  INV_X1    g0525(.A(new_n217), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G41), .ZN(new_n727));
  INV_X1    g0527(.A(G116), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n627), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT96), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n727), .A2(new_n256), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n227), .B2(new_n727), .ZN(new_n732));
  XOR2_X1   g0532(.A(new_n732), .B(KEYINPUT28), .Z(new_n733));
  NOR2_X1   g0533(.A1(new_n636), .A2(new_n638), .ZN(new_n734));
  OAI21_X1  g0534(.A(KEYINPUT84), .B1(new_n619), .B2(new_n517), .ZN(new_n735));
  INV_X1    g0535(.A(new_n640), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n616), .A2(new_n606), .A3(G190), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n734), .A2(new_n735), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n680), .A2(new_n679), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n673), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(KEYINPUT26), .B1(new_n740), .B2(new_n599), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n675), .A2(new_n676), .A3(new_n652), .A4(new_n642), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n741), .A2(new_n673), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n694), .A2(new_n569), .A3(new_n566), .ZN(new_n744));
  INV_X1    g0544(.A(new_n686), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n599), .A2(new_n604), .A3(KEYINPUT98), .ZN(new_n746));
  AOI21_X1  g0546(.A(KEYINPUT98), .B1(new_n599), .B2(new_n604), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n744), .B(new_n745), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n709), .B1(new_n743), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT29), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n701), .A2(new_n709), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n751), .B1(new_n752), .B2(new_n750), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n487), .A2(new_n505), .A3(new_n616), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n578), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT97), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(new_n563), .B2(new_n329), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n558), .A2(KEYINPUT97), .A3(G179), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n755), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT30), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n755), .A2(new_n757), .A3(new_n758), .A4(KEYINPUT30), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n558), .A2(G179), .A3(new_n678), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(new_n689), .A3(new_n578), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n709), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT31), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n765), .A2(KEYINPUT31), .A3(new_n709), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n570), .A2(new_n527), .A3(new_n654), .A4(new_n717), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n771), .A2(G330), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n753), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT99), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n733), .B1(new_n776), .B2(G1), .ZN(G364));
  NOR2_X1   g0577(.A1(new_n713), .A2(G330), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT100), .ZN(new_n779));
  INV_X1    g0579(.A(G13), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G45), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n782), .A2(KEYINPUT101), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(KEYINPUT101), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n783), .A2(G1), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n727), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n779), .B(new_n787), .C1(new_n715), .C2(new_n714), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n222), .B1(G20), .B2(new_n295), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT103), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n217), .A2(new_n247), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT102), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n796), .A2(G355), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n726), .A2(new_n247), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(G45), .B2(new_n226), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n244), .A2(new_n262), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n799), .A2(new_n800), .B1(G116), .B2(new_n217), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n794), .B1(new_n797), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n786), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n223), .A2(G179), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n804), .A2(new_n517), .A3(new_n327), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G159), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT32), .ZN(new_n808));
  NAND2_X1  g0608(.A1(G20), .A2(G179), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT104), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n810), .A2(new_n544), .A3(G200), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n810), .A2(new_n517), .A3(G200), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n202), .A2(new_n811), .B1(new_n812), .B2(new_n349), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n517), .A2(G179), .A3(G200), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n223), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n247), .B1(new_n815), .B2(new_n534), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n804), .A2(new_n517), .A3(G200), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(G107), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n804), .A2(G190), .A3(G200), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n639), .B2(new_n820), .ZN(new_n821));
  NOR4_X1   g0621(.A1(new_n808), .A2(new_n813), .A3(new_n816), .A4(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT105), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n810), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(G200), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n810), .A2(new_n823), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(new_n544), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n825), .A2(new_n517), .A3(new_n826), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n822), .B1(new_n273), .B2(new_n827), .C1(new_n303), .C2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n828), .ZN(new_n830));
  INV_X1    g0630(.A(new_n827), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n830), .A2(G311), .B1(new_n831), .B2(G322), .ZN(new_n832));
  INV_X1    g0632(.A(new_n815), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n833), .A2(new_n519), .B1(new_n806), .B2(G329), .ZN(new_n834));
  INV_X1    g0634(.A(G283), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n835), .B2(new_n817), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n360), .B1(new_n820), .B2(new_n547), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n836), .B1(KEYINPUT106), .B2(new_n837), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n837), .A2(KEYINPUT106), .ZN(new_n839));
  INV_X1    g0639(.A(new_n811), .ZN(new_n840));
  INV_X1    g0640(.A(new_n812), .ZN(new_n841));
  XNOR2_X1  g0641(.A(KEYINPUT33), .B(G317), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G326), .A2(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n832), .A2(new_n838), .A3(new_n839), .A4(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT107), .B1(new_n829), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n789), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n829), .A2(new_n844), .A3(KEYINPUT107), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n803), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n792), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n849), .B1(new_n713), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n788), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G396));
  NAND2_X1  g0653(.A1(new_n306), .A2(new_n709), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n328), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n331), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n331), .A2(new_n709), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n332), .A2(new_n709), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n752), .A2(new_n859), .B1(new_n701), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n786), .B1(new_n862), .B2(new_n773), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n773), .B2(new_n862), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n789), .A2(new_n790), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n787), .B1(new_n303), .B2(new_n865), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n639), .A2(new_n817), .B1(new_n820), .B2(new_n316), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n247), .B1(new_n806), .B2(G311), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n534), .B2(new_n815), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n867), .B(new_n869), .C1(G283), .C2(new_n841), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n547), .B2(new_n811), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(G116), .B2(new_n830), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n831), .A2(G294), .ZN(new_n873));
  AOI22_X1  g0673(.A1(G137), .A2(new_n840), .B1(new_n841), .B2(G150), .ZN(new_n874));
  INV_X1    g0674(.A(G159), .ZN(new_n875));
  INV_X1    g0675(.A(G143), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n874), .B1(new_n828), .B2(new_n875), .C1(new_n876), .C2(new_n827), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT34), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n360), .B1(new_n806), .B2(G132), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n349), .B2(new_n817), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n815), .A2(new_n273), .B1(new_n820), .B2(new_n202), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n872), .A2(new_n873), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  OAI221_X1 g0683(.A(new_n866), .B1(new_n883), .B2(new_n846), .C1(new_n791), .C2(new_n859), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n864), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(G384));
  NOR2_X1   g0686(.A1(new_n781), .A2(new_n256), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT110), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n857), .B1(new_n701), .B2(new_n861), .ZN(new_n889));
  INV_X1    g0689(.A(new_n358), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(new_n717), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n384), .A2(new_n891), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n377), .B1(new_n890), .B2(new_n717), .C1(new_n382), .C2(new_n383), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT109), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT108), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n429), .B2(new_n707), .ZN(new_n899));
  INV_X1    g0699(.A(new_n707), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n407), .A2(KEYINPUT108), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n440), .A2(new_n407), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n414), .A2(new_n415), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n424), .A2(new_n428), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n905), .B2(new_n387), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT37), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n902), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n428), .B1(KEYINPUT16), .B2(new_n427), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n910), .A2(new_n387), .B1(new_n904), .B2(new_n707), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT37), .B1(new_n903), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n707), .B1(new_n910), .B2(new_n387), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n909), .A2(new_n912), .B1(new_n444), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n897), .B1(new_n914), .B2(KEYINPUT38), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  INV_X1    g0716(.A(new_n911), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n905), .A2(new_n387), .A3(new_n433), .A4(new_n435), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n908), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n417), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n899), .B2(new_n901), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n919), .B1(new_n921), .B2(new_n908), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n444), .A2(new_n913), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n916), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n915), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n897), .B(new_n916), .C1(new_n922), .C2(new_n924), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n896), .A2(new_n929), .B1(new_n662), .B2(new_n707), .ZN(new_n930));
  INV_X1    g0730(.A(new_n377), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n717), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n926), .A2(KEYINPUT39), .A3(new_n927), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n407), .A2(KEYINPUT108), .A3(new_n900), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT108), .B1(new_n407), .B2(new_n900), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n444), .A2(new_n936), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n936), .A2(KEYINPUT37), .A3(new_n920), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n908), .B1(new_n902), .B2(new_n907), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n916), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT39), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n914), .A2(KEYINPUT38), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n932), .B1(new_n933), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n888), .B1(new_n930), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n662), .A2(new_n707), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n889), .A2(new_n895), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n948), .B1(new_n949), .B2(new_n928), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n950), .A2(KEYINPUT110), .A3(new_n945), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n665), .B1(new_n753), .B2(new_n446), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n858), .B1(new_n892), .B2(new_n893), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT40), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n955), .A2(new_n771), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n928), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n955), .A2(new_n771), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n941), .A2(new_n943), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n447), .A2(new_n771), .ZN(new_n963));
  OAI21_X1  g0763(.A(G330), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n963), .B2(new_n962), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n887), .B1(new_n954), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n966), .B2(new_n954), .ZN(new_n968));
  INV_X1    g0768(.A(new_n586), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(KEYINPUT35), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(KEYINPUT35), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n970), .A2(new_n971), .A3(G116), .A4(new_n224), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT36), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n226), .A2(new_n303), .A3(new_n397), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n349), .A2(G50), .ZN(new_n975));
  OAI211_X1 g0775(.A(G1), .B(new_n780), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n968), .A2(new_n973), .A3(new_n976), .ZN(G367));
  NOR2_X1   g0777(.A1(new_n641), .A2(new_n717), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n978), .A2(new_n650), .A3(new_n651), .A4(new_n672), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n740), .B2(new_n978), .ZN(new_n980));
  AOI21_X1  g0780(.A(KEYINPUT43), .B1(new_n980), .B2(KEYINPUT111), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(KEYINPUT111), .B2(new_n980), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n746), .A2(new_n747), .B1(new_n602), .B2(new_n717), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n675), .A2(new_n709), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(new_n724), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT42), .Z(new_n989));
  OAI21_X1  g0789(.A(new_n599), .B1(new_n985), .B2(new_n694), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n989), .B1(new_n717), .B2(new_n990), .ZN(new_n991));
  MUX2_X1   g0791(.A(new_n984), .B(new_n982), .S(new_n991), .Z(new_n992));
  NOR2_X1   g0792(.A1(new_n720), .A2(new_n987), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n992), .B(new_n993), .Z(new_n994));
  INV_X1    g0794(.A(new_n785), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n724), .B1(new_n719), .B2(new_n723), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n716), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n724), .A2(new_n721), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n987), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT44), .Z(new_n1000));
  NOR2_X1   g0800(.A1(new_n987), .A2(new_n998), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(new_n720), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n775), .B1(new_n997), .B2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n727), .B(KEYINPUT41), .Z(new_n1006));
  OAI21_X1  g0806(.A(new_n995), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n994), .A2(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n798), .A2(new_n236), .B1(new_n726), .B2(new_n643), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n787), .B1(new_n794), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(G317), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n360), .B1(new_n805), .B2(new_n1011), .C1(new_n534), .C2(new_n817), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(G107), .B2(new_n833), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G311), .A2(new_n840), .B1(new_n841), .B2(new_n519), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n820), .A2(new_n728), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT46), .Z(new_n1016));
  AND3_X1   g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n551), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1017), .B1(new_n835), .B2(new_n828), .C1(new_n1018), .C2(new_n827), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n830), .A2(G50), .B1(new_n831), .B2(G150), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n247), .B1(new_n817), .B2(new_n303), .C1(new_n815), .C2(new_n349), .ZN(new_n1021));
  INV_X1    g0821(.A(G137), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n805), .A2(new_n1022), .B1(new_n820), .B2(new_n273), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1021), .B1(KEYINPUT112), .B2(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n1023), .A2(KEYINPUT112), .B1(new_n812), .B2(new_n875), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G143), .B2(new_n840), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1020), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1019), .A2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT47), .Z(new_n1029));
  OAI221_X1 g0829(.A(new_n1010), .B1(new_n850), .B2(new_n980), .C1(new_n1029), .C2(new_n846), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1008), .A2(new_n1030), .ZN(G387));
  NAND2_X1  g0831(.A1(new_n997), .A2(new_n785), .ZN(new_n1032));
  XOR2_X1   g0832(.A(KEYINPUT115), .B(G322), .Z(new_n1033));
  AOI22_X1  g0833(.A1(new_n840), .A2(new_n1033), .B1(new_n841), .B2(G311), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n828), .B2(new_n1018), .C1(new_n1011), .C2(new_n827), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n820), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n833), .A2(G283), .B1(new_n1039), .B2(new_n519), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT116), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1042), .A2(KEYINPUT49), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(KEYINPUT49), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n817), .A2(new_n728), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n247), .B(new_n1045), .C1(G326), .C2(new_n806), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n812), .A2(new_n275), .ZN(new_n1048));
  INV_X1    g0848(.A(G150), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n247), .B1(new_n805), .B2(new_n1049), .C1(new_n534), .C2(new_n817), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n820), .A2(new_n303), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n815), .A2(new_n301), .ZN(new_n1052));
  OR3_X1    g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1048), .B(new_n1053), .C1(G159), .C2(new_n840), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n202), .B2(new_n827), .C1(new_n349), .C2(new_n828), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n846), .B1(new_n1047), .B2(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n796), .A2(new_n730), .B1(new_n316), .B2(new_n726), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n270), .A2(G50), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT114), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT50), .Z(new_n1060));
  AOI211_X1 g0860(.A(G45), .B(new_n730), .C1(G68), .C2(G77), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1060), .B1(new_n1061), .B2(KEYINPUT113), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(KEYINPUT113), .B2(new_n1061), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n233), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n798), .B1(new_n1064), .B2(new_n262), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1057), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n787), .B1(new_n1066), .B2(new_n794), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n719), .B2(new_n850), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n776), .A2(new_n997), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n727), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n776), .A2(new_n997), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1032), .B1(new_n1056), .B2(new_n1068), .C1(new_n1070), .C2(new_n1071), .ZN(G393));
  NAND3_X1  g0872(.A1(new_n776), .A2(new_n997), .A3(new_n1004), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1004), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1069), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1073), .A2(new_n727), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n794), .B1(new_n534), .B2(new_n217), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n241), .A2(new_n798), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n786), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n987), .A2(new_n792), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n827), .A2(new_n875), .B1(new_n1049), .B2(new_n811), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT51), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n828), .A2(new_n270), .B1(new_n202), .B2(new_n812), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1084), .A2(KEYINPUT117), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(KEYINPUT117), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n247), .B1(new_n805), .B2(new_n876), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n815), .A2(new_n303), .B1(new_n820), .B2(new_n349), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(G87), .C2(new_n818), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1082), .A2(new_n1085), .A3(new_n1086), .A4(new_n1089), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1090), .A2(KEYINPUT118), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n831), .A2(G311), .B1(G317), .B2(new_n840), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT52), .Z(new_n1093));
  AOI22_X1  g0893(.A1(new_n833), .A2(G116), .B1(new_n1039), .B2(G283), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n247), .B1(new_n806), .B2(new_n1033), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n819), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n551), .B2(new_n841), .ZN(new_n1097));
  INV_X1    g0897(.A(G294), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1093), .B(new_n1097), .C1(new_n1098), .C2(new_n828), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1090), .A2(KEYINPUT118), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1091), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1079), .B(new_n1080), .C1(new_n789), .C2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n1004), .B2(new_n785), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1076), .A2(new_n1103), .ZN(G390));
  NAND3_X1  g0904(.A1(new_n772), .A2(new_n859), .A3(new_n895), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT119), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n744), .A2(new_n745), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n746), .A2(new_n747), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n741), .A2(new_n673), .A3(new_n742), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n717), .B(new_n856), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n894), .B1(new_n1112), .B2(new_n857), .ZN(new_n1113));
  OAI21_X1  g0913(.A(KEYINPUT37), .B1(new_n936), .B2(new_n920), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n909), .ZN(new_n1115));
  AOI21_X1  g0915(.A(KEYINPUT38), .B1(new_n1115), .B2(new_n937), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n909), .A2(new_n912), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1117), .A2(KEYINPUT38), .A3(new_n923), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n932), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1107), .B1(new_n1113), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n932), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n941), .B2(new_n943), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n857), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n749), .B2(new_n856), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1122), .B(KEYINPUT119), .C1(new_n894), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n933), .A2(new_n944), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1121), .B1(new_n889), .B2(new_n895), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT120), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1106), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1126), .B(KEYINPUT120), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1131), .B1(new_n1134), .B2(new_n1106), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT121), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n772), .A2(new_n859), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1136), .B1(new_n1137), .B2(new_n894), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1105), .A2(new_n1124), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1137), .A2(new_n1136), .A3(new_n894), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1137), .A2(new_n894), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1105), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1140), .A2(new_n1141), .B1(new_n889), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n772), .A2(new_n447), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n665), .B(new_n1145), .C1(new_n753), .C2(new_n446), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1135), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1133), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n949), .A2(new_n932), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n933), .A2(new_n944), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT120), .B1(new_n1152), .B2(new_n1126), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1106), .B1(new_n1149), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1131), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n1155), .A3(new_n1147), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1148), .A2(new_n727), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1151), .A2(new_n790), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n828), .A2(new_n534), .B1(new_n316), .B2(new_n812), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT122), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n360), .B1(new_n805), .B2(new_n1098), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G87), .B2(new_n1039), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n833), .A2(G77), .B1(new_n818), .B2(G68), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(new_n835), .C2(new_n811), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G116), .B2(new_n831), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1161), .A2(new_n1162), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(G125), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n247), .B1(new_n805), .B2(new_n1169), .C1(new_n202), .C2(new_n817), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1039), .A2(G150), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT53), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(G159), .C2(new_n833), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n831), .A2(G132), .ZN(new_n1174));
  XOR2_X1   g0974(.A(KEYINPUT54), .B(G143), .Z(new_n1175));
  NAND2_X1  g0975(.A1(new_n830), .A2(new_n1175), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G128), .A2(new_n840), .B1(new_n841), .B2(G137), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1173), .A2(new_n1174), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n846), .B1(new_n1168), .B2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n787), .B(new_n1179), .C1(new_n275), .C2(new_n865), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1135), .A2(new_n785), .B1(new_n1158), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1157), .A2(new_n1181), .ZN(G378));
  OAI21_X1  g0982(.A(G330), .B1(new_n958), .B2(new_n961), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n294), .A2(new_n900), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT95), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n347), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n341), .A2(new_n346), .A3(KEYINPUT95), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1186), .B1(new_n1190), .B2(new_n297), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n297), .B(new_n1186), .C1(new_n656), .C2(new_n657), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1185), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n294), .B(new_n900), .C1(new_n658), .C2(new_n298), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1195), .A2(new_n1192), .A3(new_n1184), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1183), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1199), .B(G330), .C1(new_n961), .C2(new_n958), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n947), .B2(new_n951), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n896), .A2(new_n929), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1203), .A2(new_n946), .A3(new_n888), .A4(new_n948), .ZN(new_n1204));
  OAI21_X1  g1004(.A(KEYINPUT110), .B1(new_n950), .B2(new_n945), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1204), .A2(new_n1205), .A3(new_n1200), .A4(new_n1198), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1202), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1146), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n1156), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(KEYINPUT125), .B1(new_n1209), .B2(KEYINPUT57), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n727), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1209), .B2(KEYINPUT57), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT125), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT57), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1146), .B1(new_n1135), .B2(new_n1147), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1213), .B(new_n1214), .C1(new_n1215), .C2(new_n1207), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1210), .A2(new_n1212), .A3(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1207), .A2(new_n995), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1197), .A2(new_n790), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n865), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n786), .B1(G50), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n360), .A2(new_n261), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1222), .B(new_n1051), .C1(G283), .C2(new_n806), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n273), .B2(new_n817), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT123), .Z(new_n1225));
  OAI22_X1  g1025(.A1(new_n812), .A2(new_n534), .B1(new_n349), .B2(new_n815), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G116), .B2(new_n840), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n830), .A2(new_n643), .B1(new_n831), .B2(G107), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1225), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT58), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n831), .A2(G128), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n833), .A2(G150), .B1(new_n1039), .B2(new_n1175), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n1169), .B2(new_n811), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G132), .B2(new_n841), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1232), .B(new_n1235), .C1(new_n1022), .C2(new_n828), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n818), .A2(G159), .ZN(new_n1240));
  AOI211_X1 g1040(.A(G33), .B(G41), .C1(new_n806), .C2(G124), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1222), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1231), .A2(new_n1242), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1221), .B1(new_n1245), .B2(new_n789), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1218), .B1(new_n1219), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1217), .A2(new_n1247), .ZN(G375));
  OAI22_X1  g1048(.A1(new_n1098), .A2(new_n811), .B1(new_n812), .B2(new_n728), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n830), .B2(G107), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT126), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n805), .A2(new_n547), .B1(new_n820), .B2(new_n534), .ZN(new_n1252));
  XOR2_X1   g1052(.A(new_n1252), .B(KEYINPUT127), .Z(new_n1253));
  AOI211_X1 g1053(.A(new_n247), .B(new_n1052), .C1(G77), .C2(new_n818), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(new_n827), .C2(new_n835), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1251), .A2(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n827), .A2(new_n1022), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n817), .A2(new_n273), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n360), .B(new_n1258), .C1(G128), .C2(new_n806), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n840), .A2(G132), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n841), .A2(new_n1175), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n833), .A2(G50), .B1(new_n1039), .B2(G159), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1257), .B(new_n1263), .C1(G150), .C2(new_n830), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n789), .B1(new_n1256), .B2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1265), .B(new_n786), .C1(G68), .C2(new_n1220), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(new_n894), .B2(new_n790), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1144), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1267), .B1(new_n1268), .B2(new_n785), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1147), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1006), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1268), .A2(new_n1208), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1269), .B1(new_n1272), .B2(new_n1273), .ZN(G381));
  OR2_X1    g1074(.A1(G381), .A2(G384), .ZN(new_n1275));
  OR4_X1    g1075(.A1(G396), .A2(G390), .A3(new_n1275), .A4(G393), .ZN(new_n1276));
  OR4_X1    g1076(.A1(G387), .A2(new_n1276), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1077(.A(G378), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n708), .A2(G213), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G407), .B(G213), .C1(G375), .C2(new_n1281), .ZN(G409));
  NAND3_X1  g1082(.A1(new_n1217), .A2(G378), .A3(new_n1247), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1209), .A2(new_n1271), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1247), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1278), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1279), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1144), .A2(KEYINPUT60), .A3(new_n1146), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1289), .A2(new_n727), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1270), .A2(KEYINPUT60), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1290), .B1(new_n1291), .B2(new_n1273), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(G384), .A3(new_n1269), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G384), .B1(new_n1292), .B2(new_n1269), .ZN(new_n1295));
  OAI211_X1 g1095(.A(G2897), .B(new_n1280), .C1(new_n1294), .C2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1295), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1280), .A2(G2897), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n1293), .A3(new_n1298), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1296), .A2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT61), .B1(new_n1288), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT63), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1302), .B1(new_n1288), .B2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(G387), .A2(new_n1076), .A3(new_n1103), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(G393), .B(new_n852), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1008), .A2(new_n1030), .A3(G390), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1307), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1280), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(KEYINPUT63), .A3(new_n1303), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1301), .A2(new_n1305), .A3(new_n1311), .A4(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT62), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1312), .A2(new_n1315), .A3(new_n1303), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT61), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1296), .A2(new_n1299), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1317), .B1(new_n1312), .B2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1315), .B1(new_n1312), .B2(new_n1303), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(new_n1316), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1314), .B1(new_n1321), .B2(new_n1311), .ZN(G405));
  NAND2_X1  g1122(.A1(G375), .A2(new_n1278), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1283), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1303), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1323), .A2(new_n1304), .A3(new_n1283), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  OR2_X1    g1127(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1327), .B(new_n1328), .ZN(G402));
endmodule


