//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n612, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n457), .A2(KEYINPUT67), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(G567), .B2(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(KEYINPUT67), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n465), .B(KEYINPUT69), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n464), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g045(.A(G137), .B(new_n464), .C1(new_n467), .C2(new_n468), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n464), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n467), .A2(new_n468), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT70), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(new_n482), .A3(new_n464), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n479), .A2(new_n464), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n478), .B(new_n486), .C1(G124), .C2(new_n487), .ZN(G162));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n467), .B2(new_n468), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n495), .B(new_n498), .C1(new_n468), .C2(new_n467), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n493), .B1(new_n497), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G62), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n501), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(G651), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(G651), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(new_n515), .B1(new_n512), .B2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n504), .A2(new_n506), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(G88), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n516), .A2(G50), .A3(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n510), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(G166));
  NAND2_X1  g096(.A1(G63), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n513), .A2(new_n515), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n512), .A2(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(new_n517), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT73), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n516), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n528), .A2(new_n531), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n514), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n533), .A2(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n516), .A2(new_n517), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G90), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  NAND2_X1  g120(.A1(new_n533), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n542), .A2(G81), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n514), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n541), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n516), .A2(KEYINPUT74), .A3(new_n517), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n558), .A2(G91), .A3(new_n559), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n523), .A2(G53), .A3(G543), .A4(new_n524), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n516), .A2(new_n563), .A3(G53), .A4(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n517), .A2(G65), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT75), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n560), .A2(new_n565), .A3(new_n569), .ZN(G299));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n520), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n510), .A2(new_n518), .A3(new_n519), .A4(KEYINPUT76), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(G303));
  NAND3_X1  g149(.A1(new_n558), .A2(G87), .A3(new_n559), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n516), .A2(G49), .A3(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n578), .ZN(G288));
  NAND3_X1  g154(.A1(new_n558), .A2(G86), .A3(new_n559), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n516), .A2(G48), .A3(G543), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(new_n504), .B2(new_n506), .ZN(new_n584));
  AND2_X1   g159(.A1(G73), .A2(G543), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n582), .B(G651), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n584), .B2(new_n585), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT77), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n580), .A2(new_n581), .A3(new_n586), .A4(new_n588), .ZN(G305));
  XNOR2_X1  g164(.A(KEYINPUT78), .B(G85), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n542), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n533), .A2(G47), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n514), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n558), .A2(new_n559), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(G92), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n597), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n517), .A2(G66), .ZN(new_n603));
  INV_X1    g178(.A(G79), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n502), .ZN(new_n605));
  AOI22_X1  g180(.A1(G54), .A2(new_n533), .B1(new_n605), .B2(G651), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n596), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n596), .B1(new_n607), .B2(G868), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT79), .ZN(new_n611));
  INV_X1    g186(.A(G299), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(G868), .B2(new_n612), .ZN(G297));
  OAI21_X1  g188(.A(new_n611), .B1(G868), .B2(new_n612), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n607), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n607), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n485), .A2(G135), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  INV_X1    g197(.A(G111), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G2105), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(new_n487), .B2(G123), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT80), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n481), .A2(new_n472), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n628), .A2(new_n633), .ZN(G156));
  INV_X1    g209(.A(G14), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2438), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2430), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(KEYINPUT14), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT82), .Z(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n637), .B2(new_n639), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT83), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n643), .B(KEYINPUT83), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(new_n646), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n651), .B(new_n652), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  AND3_X1   g229(.A1(new_n648), .A2(new_n650), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n654), .B1(new_n648), .B2(new_n650), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n635), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n658), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(new_n655), .B2(new_n656), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n659), .A2(new_n661), .ZN(G401));
  INV_X1    g237(.A(KEYINPUT18), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n663), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(new_n632), .ZN(new_n670));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n666), .B2(KEYINPUT18), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(G2096), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  OR3_X1    g256(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(new_n681), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n677), .A2(new_n680), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n682), .B(new_n683), .C1(new_n684), .C2(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n684), .B2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(G229));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G35), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G162), .B2(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT29), .B(G2090), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G2084), .ZN(new_n702));
  INV_X1    g277(.A(G34), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n703), .A2(KEYINPUT24), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(KEYINPUT24), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n697), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G160), .B2(new_n697), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT94), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n701), .B1(new_n702), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n697), .A2(G32), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n485), .A2(G141), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT95), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n472), .A2(G105), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT26), .ZN(new_n715));
  AOI211_X1 g290(.A(new_n713), .B(new_n715), .C1(G129), .C2(new_n487), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n710), .B1(new_n717), .B2(new_n697), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT27), .B(G1996), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT31), .B(G11), .Z(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT98), .B(G28), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(KEYINPUT30), .ZN(new_n723));
  AOI21_X1  g298(.A(G29), .B1(new_n722), .B2(KEYINPUT30), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n721), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(G164), .A2(G29), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G27), .B2(G29), .ZN(new_n727));
  INV_X1    g302(.A(G2078), .ZN(new_n728));
  OAI221_X1 g303(.A(new_n725), .B1(new_n626), .B2(new_n697), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n697), .A2(G26), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT28), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n487), .A2(G128), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n464), .A2(G116), .ZN(new_n733));
  OAI21_X1  g308(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n734));
  INV_X1    g309(.A(G140), .ZN(new_n735));
  OAI221_X1 g310(.A(new_n732), .B1(new_n733), .B2(new_n734), .C1(new_n484), .C2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n731), .B1(new_n736), .B2(G29), .ZN(new_n737));
  INV_X1    g312(.A(G2067), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n729), .B(new_n739), .C1(new_n728), .C2(new_n727), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n709), .A2(new_n720), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(G16), .A2(G19), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n551), .B2(G16), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT90), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(G1341), .Z(new_n745));
  INV_X1    g320(.A(G16), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G4), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n607), .B2(new_n746), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G1348), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(G1348), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n746), .A2(G20), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT100), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT23), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n612), .B2(new_n746), .ZN(new_n754));
  INV_X1    g329(.A(G1956), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n745), .A2(new_n749), .A3(new_n750), .A4(new_n756), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n481), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(new_n464), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT91), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT25), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n485), .B2(G139), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT92), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n760), .A2(KEYINPUT92), .A3(new_n763), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n697), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n697), .B2(G33), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT93), .B(G2072), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G168), .A2(new_n746), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n746), .B2(G21), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT97), .B(G1966), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT99), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n773), .A2(new_n774), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n746), .A2(G5), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G171), .B2(new_n746), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1961), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n708), .A2(new_n702), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n777), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n771), .A2(new_n776), .A3(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n718), .A2(new_n719), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT96), .ZN(new_n785));
  NOR4_X1   g360(.A1(new_n741), .A2(new_n757), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n746), .A2(G22), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G166), .B2(new_n746), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1971), .ZN(new_n789));
  MUX2_X1   g364(.A(G6), .B(G305), .S(G16), .Z(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT32), .B(G1981), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n791), .B2(new_n790), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G23), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT88), .ZN(new_n795));
  AND3_X1   g370(.A1(new_n575), .A2(new_n795), .A3(new_n578), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n795), .B1(new_n575), .B2(new_n578), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n794), .B1(new_n798), .B2(G16), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT33), .B(G1976), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  OR3_X1    g376(.A1(new_n793), .A2(new_n801), .A3(KEYINPUT34), .ZN(new_n802));
  NOR2_X1   g377(.A1(G16), .A2(G24), .ZN(new_n803));
  INV_X1    g378(.A(G290), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G16), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1986), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n697), .A2(G25), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT86), .B1(G95), .B2(G2105), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(KEYINPUT86), .A2(G95), .A3(G2105), .ZN(new_n810));
  OAI221_X1 g385(.A(G2104), .B1(G107), .B2(new_n464), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT87), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n487), .A2(G119), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n485), .A2(G131), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n807), .B1(new_n817), .B2(new_n697), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT35), .B(G1991), .Z(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n818), .B(new_n820), .ZN(new_n821));
  AOI211_X1 g396(.A(new_n806), .B(new_n821), .C1(KEYINPUT89), .C2(KEYINPUT36), .ZN(new_n822));
  OAI21_X1  g397(.A(KEYINPUT34), .B1(new_n793), .B2(new_n801), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n802), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n786), .A2(new_n826), .A3(new_n827), .ZN(G150));
  INV_X1    g403(.A(G150), .ZN(G311));
  INV_X1    g404(.A(G55), .ZN(new_n830));
  INV_X1    g405(.A(G93), .ZN(new_n831));
  OAI22_X1  g406(.A1(new_n830), .A2(new_n532), .B1(new_n541), .B2(new_n831), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(new_n514), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n832), .A2(new_n834), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT101), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n837), .A2(new_n550), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n551), .A2(KEYINPUT101), .A3(new_n838), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n607), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n846));
  AOI21_X1  g421(.A(G860), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n846), .B2(new_n845), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n835), .A2(G860), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT37), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT102), .Z(G145));
  XNOR2_X1  g427(.A(new_n626), .B(G160), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G162), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n764), .A2(KEYINPUT103), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n736), .B(G164), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n717), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n717), .A2(new_n856), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n855), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n764), .A2(new_n765), .A3(KEYINPUT103), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n857), .A2(new_n767), .A3(new_n858), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n817), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n630), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n485), .A2(G142), .ZN(new_n866));
  INV_X1    g441(.A(G118), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT104), .B1(new_n867), .B2(G2105), .ZN(new_n868));
  INV_X1    g443(.A(G2104), .ZN(new_n869));
  NOR2_X1   g444(.A1(G106), .A2(G2105), .ZN(new_n870));
  NOR3_X1   g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n867), .A2(KEYINPUT104), .A3(G2105), .ZN(new_n872));
  AOI22_X1  g447(.A1(G130), .A2(new_n487), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n866), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n630), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n817), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n865), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n875), .B1(new_n865), .B2(new_n877), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n854), .B1(new_n863), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n883));
  NOR3_X1   g458(.A1(new_n879), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n865), .A2(new_n877), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n874), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT105), .B1(new_n886), .B2(new_n878), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n860), .B(new_n862), .C1(new_n884), .C2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(G37), .B1(new_n882), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n881), .A2(KEYINPUT105), .ZN(new_n890));
  INV_X1    g465(.A(new_n887), .ZN(new_n891));
  INV_X1    g466(.A(new_n862), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n890), .B(new_n891), .C1(new_n892), .C2(new_n859), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n888), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT106), .B1(new_n894), .B2(new_n854), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n896));
  INV_X1    g471(.A(new_n854), .ZN(new_n897));
  AOI211_X1 g472(.A(new_n896), .B(new_n897), .C1(new_n893), .C2(new_n888), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n889), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g475(.A(new_n617), .B(new_n842), .Z(new_n901));
  NAND2_X1  g476(.A1(new_n602), .A2(new_n606), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(G299), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n602), .A2(new_n612), .A3(new_n606), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n602), .A2(new_n612), .A3(new_n606), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n612), .B1(new_n602), .B2(new_n606), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n901), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n909), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(new_n901), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n798), .A2(new_n804), .ZN(new_n916));
  NAND2_X1  g491(.A1(G288), .A2(KEYINPUT88), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n575), .A2(new_n795), .A3(new_n578), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(G290), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n920), .A3(KEYINPUT108), .ZN(new_n921));
  XNOR2_X1  g496(.A(G305), .B(G166), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n916), .A2(new_n920), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n924), .A2(KEYINPUT108), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n921), .A2(new_n922), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n912), .B(new_n928), .C1(new_n913), .C2(new_n901), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n915), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n927), .B1(new_n915), .B2(new_n929), .ZN(new_n931));
  OAI21_X1  g506(.A(G868), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n838), .A2(G868), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(G295));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n933), .ZN(G331));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n936));
  NAND2_X1  g511(.A1(G301), .A2(KEYINPUT109), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n539), .A2(new_n540), .A3(new_n543), .A4(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(G286), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(G171), .A2(G168), .A3(new_n938), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n842), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n840), .A2(new_n940), .A3(new_n941), .A4(new_n841), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n909), .B(new_n943), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(new_n944), .ZN(new_n949));
  INV_X1    g524(.A(new_n910), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n903), .A2(new_n905), .A3(new_n950), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n949), .B(new_n951), .C1(new_n909), .C2(KEYINPUT41), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n925), .A2(new_n926), .ZN(new_n954));
  INV_X1    g529(.A(new_n923), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n911), .ZN(new_n959));
  AND4_X1   g534(.A1(new_n903), .A2(new_n943), .A3(new_n905), .A4(new_n944), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(new_n927), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G37), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n957), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n936), .B1(new_n964), .B2(KEYINPUT43), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n960), .B1(new_n958), .B2(new_n911), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT43), .B1(new_n966), .B2(new_n927), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n956), .B1(new_n966), .B2(KEYINPUT111), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n969));
  AOI211_X1 g544(.A(new_n969), .B(new_n960), .C1(new_n911), .C2(new_n958), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n963), .B(new_n967), .C1(new_n968), .C2(new_n970), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n965), .A2(KEYINPUT112), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT112), .B1(new_n965), .B2(new_n971), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n963), .B(new_n962), .C1(new_n968), .C2(new_n970), .ZN(new_n974));
  AOI21_X1  g549(.A(G37), .B1(new_n953), .B2(new_n956), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n974), .A2(KEYINPUT43), .B1(new_n967), .B2(new_n975), .ZN(new_n976));
  OAI22_X1  g551(.A1(new_n972), .A2(new_n973), .B1(KEYINPUT44), .B2(new_n976), .ZN(G397));
  INV_X1    g552(.A(G1996), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n717), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n736), .B(G2067), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  INV_X1    g557(.A(new_n499), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n498), .B1(new_n481), .B2(new_n495), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n982), .B1(new_n985), .B2(new_n493), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n987));
  INV_X1    g562(.A(G40), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n470), .A2(new_n474), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT113), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(G1996), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n981), .A2(new_n991), .B1(new_n717), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n817), .B(new_n820), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n994), .A2(KEYINPUT114), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(KEYINPUT114), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(new_n991), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n990), .ZN(new_n999));
  XNOR2_X1  g574(.A(G290), .B(G1986), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT123), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n982), .B(new_n1004), .C1(new_n985), .C2(new_n493), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n497), .A2(new_n499), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n489), .A2(new_n492), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1384), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1005), .B(KEYINPUT116), .C1(new_n1006), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n1011), .A3(new_n1004), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n466), .A2(new_n469), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G2105), .ZN(new_n1015));
  INV_X1    g590(.A(new_n474), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(G40), .A3(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(G2084), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n987), .B1(G164), .B2(G1384), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT45), .B(new_n982), .C1(new_n985), .C2(new_n493), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n989), .A3(new_n1020), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1013), .A2(new_n1018), .B1(new_n774), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1002), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(KEYINPUT117), .B(G8), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G286), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1021), .A2(new_n774), .ZN(new_n1028));
  NOR4_X1   g603(.A1(G164), .A2(KEYINPUT116), .A3(G1384), .A4(new_n1003), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n986), .A2(KEYINPUT50), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1011), .B1(new_n1009), .B2(new_n1004), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1018), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1028), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(KEYINPUT123), .A3(G8), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1024), .A2(new_n1027), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT51), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT124), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT51), .B1(G286), .B2(new_n1026), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI211_X1 g615(.A(new_n1038), .B(new_n1040), .C1(new_n1034), .C2(new_n1026), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1028), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1033), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1026), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT124), .B1(new_n1044), .B2(new_n1039), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1037), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT62), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G1976), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n796), .A2(new_n797), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n989), .A2(new_n1009), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n1026), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT52), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1053), .ZN(new_n1055));
  INV_X1    g630(.A(new_n581), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(G1981), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n580), .A2(new_n1057), .A3(new_n586), .A4(new_n588), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n516), .A2(G86), .A3(new_n517), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n588), .A2(new_n581), .A3(new_n586), .A4(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G1981), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n1061), .A3(KEYINPUT49), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1063));
  XOR2_X1   g638(.A(KEYINPUT118), .B(KEYINPUT49), .Z(new_n1064));
  OAI211_X1 g639(.A(new_n1055), .B(new_n1062), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT52), .B1(G288), .B2(new_n1050), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1055), .B(new_n1066), .C1(new_n919), .C2(new_n1050), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1054), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT126), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n572), .A2(G8), .A3(new_n573), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n572), .A2(KEYINPUT55), .A3(G8), .A4(new_n573), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1971), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1021), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G2090), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n989), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1078), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1074), .B(G8), .C1(new_n1076), .C2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n989), .B1(new_n1009), .B2(new_n1004), .ZN(new_n1081));
  NOR3_X1   g656(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1083), .A2(new_n1077), .B1(new_n1021), .B2(new_n1075), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1072), .B(new_n1073), .C1(new_n1084), .C2(new_n1025), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1068), .A2(new_n1069), .A3(new_n1080), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1080), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1054), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT126), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1048), .B1(new_n1037), .B2(new_n1046), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1017), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n1094), .A2(G1961), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1021), .B2(G2078), .ZN(new_n1097));
  OR3_X1    g672(.A1(new_n1021), .A2(new_n1096), .A3(G2078), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1099), .A2(G171), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1049), .A2(new_n1090), .A3(new_n1093), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1044), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G168), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT63), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1085), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1080), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1068), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1108), .A2(new_n1023), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1102), .B(G168), .C1(new_n1109), .C2(new_n1074), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT63), .B1(new_n1110), .B2(new_n1088), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1053), .B(KEYINPUT119), .ZN(new_n1112));
  AND4_X1   g687(.A1(new_n1050), .A2(new_n1065), .A3(new_n575), .A4(new_n578), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1058), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1107), .A2(new_n1111), .A3(new_n1115), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT58), .B(G1341), .Z(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n986), .B2(new_n1017), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1019), .A2(new_n978), .A3(new_n1020), .A4(new_n989), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1052), .A2(KEYINPUT120), .A3(new_n1117), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n551), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT59), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1126), .A3(new_n551), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT57), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n560), .A2(new_n565), .A3(new_n1130), .A4(new_n569), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n755), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT56), .B(G2072), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1019), .A2(new_n989), .A3(new_n1020), .A4(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1134), .A2(new_n1129), .A3(new_n1131), .A4(new_n1136), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT121), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1137), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1142), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1134), .A2(new_n1136), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1138), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1128), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1128), .A2(new_n1144), .A3(KEYINPUT122), .A4(new_n1147), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1052), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n738), .ZN(new_n1153));
  OAI211_X1 g728(.A(KEYINPUT60), .B(new_n1153), .C1(new_n1094), .C2(G1348), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(new_n607), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1094), .B2(G1348), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT60), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1150), .A2(new_n1151), .A3(new_n1159), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1156), .A2(new_n607), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1142), .B1(new_n1161), .B2(new_n1146), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(G301), .B(KEYINPUT54), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1095), .A2(new_n1164), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1165));
  AOI211_X1 g740(.A(new_n1096), .B(G2078), .C1(new_n1017), .C2(KEYINPUT125), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n1017), .A2(KEYINPUT125), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1166), .A2(new_n1019), .A3(new_n1020), .A4(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1168), .B(new_n1097), .C1(new_n1094), .C2(G1961), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1165), .B1(new_n1170), .B2(new_n1164), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1086), .A2(new_n1089), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1091), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1116), .B1(new_n1163), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1101), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI211_X1 g751(.A(KEYINPUT127), .B(new_n1116), .C1(new_n1163), .C2(new_n1173), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1001), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n717), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n991), .B1(new_n1179), .B2(new_n980), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n992), .B(KEYINPUT46), .Z(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT47), .Z(new_n1183));
  INV_X1    g758(.A(new_n991), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n993), .A2(new_n819), .A3(new_n817), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n736), .A2(G2067), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n998), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n990), .A2(G290), .A3(G1986), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT48), .Z(new_n1190));
  AOI211_X1 g765(.A(new_n1183), .B(new_n1187), .C1(new_n1188), .C2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1178), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g767(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n975), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g770(.A1(new_n462), .A2(G227), .ZN(new_n1197));
  OAI21_X1  g771(.A(new_n1197), .B1(new_n694), .B2(new_n695), .ZN(new_n1198));
  AOI21_X1  g772(.A(new_n1198), .B1(new_n659), .B2(new_n661), .ZN(new_n1199));
  AND3_X1   g773(.A1(new_n1196), .A2(new_n899), .A3(new_n1199), .ZN(G308));
  NAND3_X1  g774(.A1(new_n1196), .A2(new_n899), .A3(new_n1199), .ZN(G225));
endmodule


