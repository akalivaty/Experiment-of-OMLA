// Benchmark "locked_c1908" written by ABC on Sat Dec 16 10:46:19 2023

module locked_c1908 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110,
    G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146,
    G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478,
    G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104,
    G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140,
    G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472,
    G475, G478, G898, G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n123, new_n124, new_n125, new_n126, new_n127, new_n128, new_n129,
    new_n130, new_n131, new_n132, new_n133, new_n134, new_n135, new_n136,
    new_n137, new_n138, new_n139, new_n140, new_n141, new_n142, new_n143,
    new_n144, new_n145, new_n146, new_n147, new_n148, new_n149, new_n150,
    new_n151, new_n152, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191, new_n192,
    new_n193, new_n194, new_n195, new_n196, new_n197, new_n198, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n324, new_n325,
    new_n326, new_n327, new_n328, new_n329, new_n330, new_n331, new_n332,
    new_n333, new_n334, new_n335, new_n336, new_n337, new_n338, new_n339,
    new_n340, new_n341, new_n342, new_n343, new_n344, new_n345, new_n346,
    new_n347, new_n348, new_n349, new_n350, new_n351, new_n352, new_n353,
    new_n354, new_n355, new_n356, new_n357, new_n358, new_n359, new_n360,
    new_n361, new_n362, new_n363, new_n364, new_n365, new_n366, new_n367,
    new_n368, new_n369, new_n370, new_n371, new_n372, new_n373, new_n374,
    new_n375, new_n376, new_n377, new_n378, new_n379, new_n380, new_n381,
    new_n382, new_n383, new_n384, new_n385, new_n386, new_n387, new_n388,
    new_n389, new_n390, new_n391, new_n392, new_n393, new_n394, new_n395,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423,
    new_n424, new_n425, new_n426, new_n427, new_n428, new_n429, new_n430,
    new_n431, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n449, new_n450, new_n451, new_n452, new_n454,
    new_n455, new_n456, new_n457, new_n458, new_n459, new_n460, new_n461,
    new_n462, new_n463, new_n465, new_n466, new_n467, new_n468, new_n469,
    new_n470, new_n471, new_n473, new_n474, new_n475, new_n476, new_n477,
    new_n478, new_n479, new_n480, new_n481, new_n482, new_n483, new_n484,
    new_n485, new_n487, new_n488, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n497, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n508, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n525, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707;
  INV_X1    g000(.A(G134), .ZN(new_n123));
  OAI21_X1  g001(.A(KEYINPUT11), .B1(new_n123), .B2(G137), .ZN(new_n124));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n125));
  INV_X1    g003(.A(G137), .ZN(new_n126));
  NAND3_X1  g004(.A1(new_n125), .A2(new_n126), .A3(G134), .ZN(new_n127));
  NAND2_X1  g005(.A1(new_n124), .A2(new_n127), .ZN(new_n128));
  INV_X1    g006(.A(G131), .ZN(new_n129));
  NAND2_X1  g007(.A1(new_n123), .A2(G137), .ZN(new_n130));
  AND3_X1   g008(.A1(new_n128), .A2(new_n129), .A3(new_n130), .ZN(new_n131));
  AOI21_X1  g009(.A(new_n129), .B1(new_n128), .B2(new_n130), .ZN(new_n132));
  INV_X1    g010(.A(G146), .ZN(new_n133));
  NAND2_X1  g011(.A1(new_n133), .A2(G143), .ZN(new_n134));
  INV_X1    g012(.A(G143), .ZN(new_n135));
  NAND2_X1  g013(.A1(new_n135), .A2(G146), .ZN(new_n136));
  INV_X1    g014(.A(G128), .ZN(new_n137));
  NAND3_X1  g015(.A1(new_n134), .A2(new_n136), .A3(new_n137), .ZN(new_n138));
  AOI21_X1  g016(.A(new_n137), .B1(new_n134), .B2(new_n136), .ZN(new_n139));
  OAI21_X1  g017(.A(new_n138), .B1(new_n139), .B2(KEYINPUT0), .ZN(new_n140));
  XNOR2_X1  g018(.A(G143), .B(G146), .ZN(new_n141));
  INV_X1    g019(.A(KEYINPUT0), .ZN(new_n142));
  NOR3_X1   g020(.A1(new_n141), .A2(new_n142), .A3(new_n137), .ZN(new_n143));
  OAI22_X1  g021(.A1(new_n131), .A2(new_n132), .B1(new_n140), .B2(new_n143), .ZN(new_n144));
  INV_X1    g022(.A(G119), .ZN(new_n145));
  NAND2_X1  g023(.A1(new_n145), .A2(G116), .ZN(new_n146));
  INV_X1    g024(.A(G116), .ZN(new_n147));
  NAND2_X1  g025(.A1(new_n147), .A2(G119), .ZN(new_n148));
  NAND2_X1  g026(.A1(new_n146), .A2(new_n148), .ZN(new_n149));
  XNOR2_X1  g027(.A(KEYINPUT2), .B(G113), .ZN(new_n150));
  XNOR2_X1  g028(.A(new_n149), .B(new_n150), .ZN(new_n151));
  INV_X1    g029(.A(new_n151), .ZN(new_n152));
  NAND3_X1  g030(.A1(new_n128), .A2(new_n129), .A3(new_n130), .ZN(new_n153));
  NAND2_X1  g031(.A1(new_n134), .A2(new_n136), .ZN(new_n154));
  NAND2_X1  g032(.A1(new_n134), .A2(KEYINPUT1), .ZN(new_n155));
  NAND3_X1  g033(.A1(new_n154), .A2(new_n155), .A3(G128), .ZN(new_n156));
  OAI211_X1 g034(.A(new_n134), .B(new_n136), .C1(KEYINPUT1), .C2(new_n137), .ZN(new_n157));
  NAND2_X1  g035(.A1(new_n126), .A2(G134), .ZN(new_n158));
  NAND2_X1  g036(.A1(new_n158), .A2(new_n130), .ZN(new_n159));
  NAND2_X1  g037(.A1(new_n159), .A2(G131), .ZN(new_n160));
  NAND4_X1  g038(.A1(new_n153), .A2(new_n156), .A3(new_n157), .A4(new_n160), .ZN(new_n161));
  NAND3_X1  g039(.A1(new_n144), .A2(new_n152), .A3(new_n161), .ZN(new_n162));
  INV_X1    g040(.A(new_n162), .ZN(new_n163));
  AOI21_X1  g041(.A(new_n152), .B1(new_n144), .B2(new_n161), .ZN(new_n164));
  OAI21_X1  g042(.A(KEYINPUT28), .B1(new_n163), .B2(new_n164), .ZN(new_n165));
  XNOR2_X1  g043(.A(KEYINPUT26), .B(G101), .ZN(new_n166));
  XNOR2_X1  g044(.A(new_n166), .B(KEYINPUT27), .ZN(new_n167));
  NOR2_X1   g045(.A1(G237), .A2(G953), .ZN(new_n168));
  NAND2_X1  g046(.A1(new_n168), .A2(G210), .ZN(new_n169));
  XNOR2_X1  g047(.A(new_n167), .B(new_n169), .ZN(new_n170));
  INV_X1    g048(.A(KEYINPUT28), .ZN(new_n171));
  NAND2_X1  g049(.A1(new_n162), .A2(new_n171), .ZN(new_n172));
  NAND3_X1  g050(.A1(new_n165), .A2(new_n170), .A3(new_n172), .ZN(new_n173));
  NAND2_X1  g051(.A1(new_n173), .A2(KEYINPUT29), .ZN(new_n174));
  INV_X1    g052(.A(KEYINPUT29), .ZN(new_n175));
  NAND4_X1  g053(.A1(new_n165), .A2(new_n175), .A3(new_n170), .A4(new_n172), .ZN(new_n176));
  INV_X1    g054(.A(KEYINPUT30), .ZN(new_n177));
  AND3_X1   g055(.A1(new_n144), .A2(new_n177), .A3(new_n161), .ZN(new_n178));
  AOI21_X1  g056(.A(new_n177), .B1(new_n144), .B2(new_n161), .ZN(new_n179));
  OAI21_X1  g057(.A(new_n151), .B1(new_n178), .B2(new_n179), .ZN(new_n180));
  NAND2_X1  g058(.A1(new_n180), .A2(new_n162), .ZN(new_n181));
  INV_X1    g059(.A(new_n170), .ZN(new_n182));
  NAND2_X1  g060(.A1(new_n181), .A2(new_n182), .ZN(new_n183));
  AND3_X1   g061(.A1(new_n174), .A2(new_n176), .A3(new_n183), .ZN(new_n184));
  OAI21_X1  g062(.A(G472), .B1(new_n184), .B2(G902), .ZN(new_n185));
  INV_X1    g063(.A(KEYINPUT32), .ZN(new_n186));
  NAND4_X1  g064(.A1(new_n180), .A2(KEYINPUT31), .A3(new_n170), .A4(new_n162), .ZN(new_n187));
  INV_X1    g065(.A(G902), .ZN(new_n188));
  NAND2_X1  g066(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  AND3_X1   g067(.A1(new_n134), .A2(new_n136), .A3(new_n137), .ZN(new_n190));
  NAND2_X1  g068(.A1(new_n154), .A2(G128), .ZN(new_n191));
  AOI21_X1  g069(.A(new_n190), .B1(new_n191), .B2(new_n142), .ZN(new_n192));
  NAND2_X1  g070(.A1(new_n139), .A2(KEYINPUT0), .ZN(new_n193));
  AOI21_X1  g071(.A(new_n125), .B1(G134), .B2(new_n126), .ZN(new_n194));
  NOR3_X1   g072(.A1(new_n123), .A2(KEYINPUT11), .A3(G137), .ZN(new_n195));
  OAI21_X1  g073(.A(new_n130), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g074(.A1(new_n196), .A2(G131), .ZN(new_n197));
  AOI22_X1  g075(.A1(new_n192), .A2(new_n193), .B1(new_n197), .B2(new_n153), .ZN(new_n198));
  INV_X1    g076(.A(new_n161), .ZN(new_n199));
  OAI21_X1  g077(.A(new_n151), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  AOI21_X1  g078(.A(new_n171), .B1(new_n200), .B2(new_n162), .ZN(new_n201));
  INV_X1    g079(.A(new_n172), .ZN(new_n202));
  OAI21_X1  g080(.A(new_n182), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  OAI21_X1  g081(.A(KEYINPUT30), .B1(new_n198), .B2(new_n199), .ZN(new_n204));
  NAND3_X1  g082(.A1(new_n144), .A2(new_n177), .A3(new_n161), .ZN(new_n205));
  NAND2_X1  g083(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g084(.A(new_n163), .B1(new_n206), .B2(new_n151), .ZN(new_n207));
  AOI21_X1  g085(.A(KEYINPUT31), .B1(new_n207), .B2(new_n170), .ZN(new_n208));
  AOI21_X1  g086(.A(new_n189), .B1(new_n203), .B2(new_n208), .ZN(new_n209));
  INV_X1    g087(.A(G472), .ZN(new_n210));
  AOI21_X1  g088(.A(new_n186), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g089(.A(new_n189), .ZN(new_n212));
  INV_X1    g090(.A(KEYINPUT31), .ZN(new_n213));
  NAND3_X1  g091(.A1(new_n180), .A2(new_n170), .A3(new_n162), .ZN(new_n214));
  NAND3_X1  g092(.A1(new_n203), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND4_X1  g093(.A1(new_n212), .A2(new_n215), .A3(new_n186), .A4(new_n210), .ZN(new_n216));
  INV_X1    g094(.A(new_n216), .ZN(new_n217));
  OAI21_X1  g095(.A(new_n185), .B1(new_n211), .B2(new_n217), .ZN(new_n218));
  INV_X1    g096(.A(G217), .ZN(new_n219));
  AOI21_X1  g097(.A(new_n219), .B1(G234), .B2(new_n188), .ZN(new_n220));
  INV_X1    g098(.A(G125), .ZN(new_n221));
  NAND2_X1  g099(.A1(new_n221), .A2(G140), .ZN(new_n222));
  INV_X1    g100(.A(KEYINPUT16), .ZN(new_n223));
  INV_X1    g101(.A(G140), .ZN(new_n224));
  AOI21_X1  g102(.A(new_n223), .B1(G125), .B2(new_n224), .ZN(new_n225));
  NOR3_X1   g103(.A1(new_n221), .A2(KEYINPUT16), .A3(G140), .ZN(new_n226));
  OAI21_X1  g104(.A(new_n222), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g105(.A1(new_n227), .A2(G146), .ZN(new_n228));
  OAI211_X1 g106(.A(new_n133), .B(new_n222), .C1(new_n225), .C2(new_n226), .ZN(new_n229));
  NAND2_X1  g107(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g108(.A(KEYINPUT23), .ZN(new_n231));
  OAI21_X1  g109(.A(new_n231), .B1(new_n145), .B2(G128), .ZN(new_n232));
  NAND3_X1  g110(.A1(new_n137), .A2(KEYINPUT23), .A3(G119), .ZN(new_n233));
  OAI211_X1 g111(.A(new_n232), .B(new_n233), .C1(G119), .C2(new_n137), .ZN(new_n234));
  XOR2_X1   g112(.A(KEYINPUT24), .B(G110), .Z(new_n235));
  XNOR2_X1  g113(.A(G119), .B(G128), .ZN(new_n236));
  AOI22_X1  g114(.A1(new_n234), .A2(G110), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g115(.A1(new_n230), .A2(new_n237), .ZN(new_n238));
  OAI22_X1  g116(.A1(new_n234), .A2(G110), .B1(new_n235), .B2(new_n236), .ZN(new_n239));
  NAND2_X1  g117(.A1(new_n224), .A2(G125), .ZN(new_n240));
  NAND3_X1  g118(.A1(new_n222), .A2(new_n240), .A3(new_n133), .ZN(new_n241));
  NAND3_X1  g119(.A1(new_n239), .A2(new_n228), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g120(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  INV_X1    g121(.A(G953), .ZN(new_n244));
  NAND3_X1  g122(.A1(new_n244), .A2(G221), .A3(G234), .ZN(new_n245));
  XNOR2_X1  g123(.A(new_n245), .B(KEYINPUT22), .ZN(new_n246));
  XNOR2_X1  g124(.A(new_n246), .B(G137), .ZN(new_n247));
  INV_X1    g125(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g126(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g127(.A1(new_n247), .A2(new_n238), .A3(new_n242), .ZN(new_n250));
  NAND3_X1  g128(.A1(new_n249), .A2(new_n188), .A3(new_n250), .ZN(new_n251));
  INV_X1    g129(.A(KEYINPUT25), .ZN(new_n252));
  AND2_X1   g130(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g131(.A1(new_n251), .A2(new_n252), .ZN(new_n254));
  OAI21_X1  g132(.A(new_n220), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OR2_X1    g133(.A1(new_n251), .A2(new_n220), .ZN(new_n256));
  NAND2_X1  g134(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g135(.A(new_n257), .ZN(new_n258));
  INV_X1    g136(.A(G469), .ZN(new_n259));
  INV_X1    g137(.A(G104), .ZN(new_n260));
  NAND2_X1  g138(.A1(new_n260), .A2(G107), .ZN(new_n261));
  INV_X1    g139(.A(G107), .ZN(new_n262));
  NAND3_X1  g140(.A1(new_n262), .A2(KEYINPUT3), .A3(G104), .ZN(new_n263));
  INV_X1    g141(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g142(.A(KEYINPUT3), .B1(new_n262), .B2(G104), .ZN(new_n265));
  OAI21_X1  g143(.A(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g144(.A1(new_n266), .A2(KEYINPUT4), .A3(G101), .ZN(new_n267));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n268));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n269));
  OAI21_X1  g147(.A(new_n269), .B1(new_n260), .B2(G107), .ZN(new_n270));
  AOI22_X1  g148(.A1(new_n270), .A2(new_n263), .B1(new_n260), .B2(G107), .ZN(new_n271));
  INV_X1    g149(.A(G101), .ZN(new_n272));
  OAI21_X1  g150(.A(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI211_X1 g151(.A(new_n272), .B(new_n261), .C1(new_n264), .C2(new_n265), .ZN(new_n274));
  NAND3_X1  g152(.A1(new_n267), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g153(.A(new_n142), .B1(new_n141), .B2(new_n137), .ZN(new_n276));
  NAND3_X1  g154(.A1(new_n193), .A2(new_n276), .A3(new_n138), .ZN(new_n277));
  NAND2_X1  g155(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g156(.A1(new_n131), .A2(new_n132), .ZN(new_n279));
  NAND2_X1  g157(.A1(new_n262), .A2(G104), .ZN(new_n280));
  AOI21_X1  g158(.A(new_n272), .B1(new_n280), .B2(new_n261), .ZN(new_n281));
  AOI21_X1  g159(.A(new_n281), .B1(new_n271), .B2(new_n272), .ZN(new_n282));
  NAND4_X1  g160(.A1(new_n282), .A2(KEYINPUT10), .A3(new_n157), .A4(new_n156), .ZN(new_n283));
  INV_X1    g161(.A(KEYINPUT10), .ZN(new_n284));
  INV_X1    g162(.A(new_n281), .ZN(new_n285));
  NAND2_X1  g163(.A1(new_n274), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g164(.A1(new_n156), .A2(new_n157), .ZN(new_n287));
  OAI21_X1  g165(.A(new_n284), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND4_X1  g166(.A1(new_n278), .A2(new_n279), .A3(new_n283), .A4(new_n288), .ZN(new_n289));
  INV_X1    g167(.A(new_n279), .ZN(new_n290));
  NOR2_X1   g168(.A1(new_n286), .A2(new_n287), .ZN(new_n291));
  AOI22_X1  g169(.A1(new_n274), .A2(new_n285), .B1(new_n156), .B2(new_n157), .ZN(new_n292));
  OAI21_X1  g170(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g171(.A1(new_n293), .A2(KEYINPUT12), .ZN(new_n294));
  XNOR2_X1  g172(.A(G110), .B(G140), .ZN(new_n295));
  INV_X1    g173(.A(G227), .ZN(new_n296));
  NOR2_X1   g174(.A1(new_n296), .A2(G953), .ZN(new_n297));
  XNOR2_X1  g175(.A(new_n295), .B(new_n297), .ZN(new_n298));
  INV_X1    g176(.A(new_n298), .ZN(new_n299));
  INV_X1    g177(.A(KEYINPUT12), .ZN(new_n300));
  OAI211_X1 g178(.A(new_n290), .B(new_n300), .C1(new_n291), .C2(new_n292), .ZN(new_n301));
  AND4_X1   g179(.A1(new_n289), .A2(new_n294), .A3(new_n299), .A4(new_n301), .ZN(new_n302));
  AND2_X1   g180(.A1(new_n275), .A2(new_n277), .ZN(new_n303));
  NAND2_X1  g181(.A1(new_n288), .A2(new_n283), .ZN(new_n304));
  OAI21_X1  g182(.A(new_n290), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g183(.A(new_n299), .B1(new_n305), .B2(new_n289), .ZN(new_n306));
  OAI211_X1 g184(.A(new_n259), .B(new_n188), .C1(new_n302), .C2(new_n306), .ZN(new_n307));
  NOR2_X1   g185(.A1(new_n259), .A2(new_n188), .ZN(new_n308));
  INV_X1    g186(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g187(.A1(new_n294), .A2(new_n289), .A3(new_n301), .ZN(new_n310));
  NAND2_X1  g188(.A1(new_n310), .A2(new_n298), .ZN(new_n311));
  NAND3_X1  g189(.A1(new_n305), .A2(new_n289), .A3(new_n299), .ZN(new_n312));
  NAND3_X1  g190(.A1(new_n311), .A2(G469), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g191(.A1(new_n307), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g192(.A(KEYINPUT9), .B(G234), .ZN(new_n315));
  OAI21_X1  g193(.A(G221), .B1(new_n315), .B2(G902), .ZN(new_n316));
  NAND2_X1  g194(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g195(.A(G214), .B1(G237), .B2(G902), .ZN(new_n318));
  NAND2_X1  g196(.A1(new_n277), .A2(G125), .ZN(new_n319));
  NAND3_X1  g197(.A1(new_n156), .A2(new_n221), .A3(new_n157), .ZN(new_n320));
  NAND2_X1  g198(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g199(.A(G224), .ZN(new_n322));
  NOR2_X1   g200(.A1(new_n322), .A2(G953), .ZN(new_n323));
  XOR2_X1   g201(.A(new_n321), .B(new_n323), .Z(new_n324));
  NAND2_X1  g202(.A1(new_n275), .A2(new_n151), .ZN(new_n325));
  INV_X1    g203(.A(KEYINPUT5), .ZN(new_n326));
  OAI21_X1  g204(.A(new_n326), .B1(new_n147), .B2(G119), .ZN(new_n327));
  NAND3_X1  g205(.A1(new_n145), .A2(KEYINPUT5), .A3(G116), .ZN(new_n328));
  NAND3_X1  g206(.A1(new_n327), .A2(new_n148), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g207(.A1(new_n329), .A2(G113), .ZN(new_n330));
  OAI21_X1  g208(.A(new_n330), .B1(new_n150), .B2(new_n149), .ZN(new_n331));
  OR2_X1    g209(.A1(new_n331), .A2(new_n286), .ZN(new_n332));
  XNOR2_X1  g210(.A(G110), .B(G122), .ZN(new_n333));
  NAND3_X1  g211(.A1(new_n325), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g212(.A(new_n333), .B1(new_n325), .B2(new_n332), .ZN(new_n335));
  OAI21_X1  g213(.A(new_n334), .B1(new_n335), .B2(KEYINPUT6), .ZN(new_n336));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n337));
  AOI211_X1 g215(.A(new_n337), .B(new_n333), .C1(new_n325), .C2(new_n332), .ZN(new_n338));
  OAI21_X1  g216(.A(new_n324), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g217(.A(G210), .B1(G237), .B2(G902), .ZN(new_n340));
  OAI21_X1  g218(.A(KEYINPUT7), .B1(new_n322), .B2(G953), .ZN(new_n341));
  NAND2_X1  g219(.A1(new_n321), .A2(new_n341), .ZN(new_n342));
  INV_X1    g220(.A(new_n341), .ZN(new_n343));
  NAND3_X1  g221(.A1(new_n319), .A2(new_n320), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g222(.A(new_n331), .B(new_n286), .ZN(new_n345));
  XNOR2_X1  g223(.A(new_n333), .B(KEYINPUT8), .ZN(new_n346));
  AOI22_X1  g224(.A1(new_n342), .A2(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g225(.A(G902), .B1(new_n347), .B2(new_n334), .ZN(new_n348));
  AND3_X1   g226(.A1(new_n339), .A2(new_n340), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g227(.A(new_n340), .B1(new_n339), .B2(new_n348), .ZN(new_n350));
  OAI21_X1  g228(.A(new_n318), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g229(.A1(new_n317), .A2(new_n351), .ZN(new_n352));
  INV_X1    g230(.A(G478), .ZN(new_n353));
  OR2_X1    g231(.A1(new_n353), .A2(KEYINPUT15), .ZN(new_n354));
  NAND2_X1  g232(.A1(new_n135), .A2(G128), .ZN(new_n355));
  NAND2_X1  g233(.A1(new_n137), .A2(G143), .ZN(new_n356));
  NAND2_X1  g234(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g235(.A(KEYINPUT13), .ZN(new_n358));
  NAND2_X1  g236(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g237(.A1(new_n357), .A2(new_n359), .A3(G134), .ZN(new_n360));
  OAI211_X1 g238(.A(new_n355), .B(new_n356), .C1(new_n358), .C2(new_n123), .ZN(new_n361));
  INV_X1    g239(.A(G122), .ZN(new_n362));
  NAND2_X1  g240(.A1(new_n362), .A2(G116), .ZN(new_n363));
  NAND2_X1  g241(.A1(new_n147), .A2(G122), .ZN(new_n364));
  NAND2_X1  g242(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g243(.A1(new_n365), .A2(G107), .ZN(new_n366));
  AOI21_X1  g244(.A(new_n262), .B1(new_n363), .B2(new_n364), .ZN(new_n367));
  OAI211_X1 g245(.A(new_n360), .B(new_n361), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g246(.A1(new_n363), .A2(KEYINPUT14), .ZN(new_n369));
  NAND3_X1  g247(.A1(new_n365), .A2(new_n369), .A3(G107), .ZN(new_n370));
  OAI211_X1 g248(.A(new_n363), .B(new_n364), .C1(KEYINPUT14), .C2(new_n262), .ZN(new_n371));
  NOR2_X1   g249(.A1(new_n357), .A2(G134), .ZN(new_n372));
  AOI21_X1  g250(.A(new_n123), .B1(new_n355), .B2(new_n356), .ZN(new_n373));
  OAI211_X1 g251(.A(new_n370), .B(new_n371), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g252(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  NOR3_X1   g253(.A1(new_n315), .A2(new_n219), .A3(G953), .ZN(new_n376));
  INV_X1    g254(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g255(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g256(.A(new_n376), .B1(new_n368), .B2(new_n374), .ZN(new_n379));
  OR2_X1    g257(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g258(.A(new_n354), .B1(new_n380), .B2(new_n188), .ZN(new_n381));
  OAI211_X1 g259(.A(new_n188), .B(new_n354), .C1(new_n378), .C2(new_n379), .ZN(new_n382));
  INV_X1    g260(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g261(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g262(.A1(new_n168), .A2(G143), .A3(G214), .ZN(new_n385));
  INV_X1    g263(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g264(.A(G143), .B1(new_n168), .B2(G214), .ZN(new_n387));
  OAI21_X1  g265(.A(G131), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g266(.A1(new_n168), .A2(G214), .ZN(new_n389));
  NAND2_X1  g267(.A1(new_n389), .A2(new_n135), .ZN(new_n390));
  NAND3_X1  g268(.A1(new_n390), .A2(new_n129), .A3(new_n385), .ZN(new_n391));
  INV_X1    g269(.A(KEYINPUT17), .ZN(new_n392));
  NAND3_X1  g270(.A1(new_n388), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  OAI211_X1 g271(.A(KEYINPUT17), .B(G131), .C1(new_n386), .C2(new_n387), .ZN(new_n394));
  NAND4_X1  g272(.A1(new_n393), .A2(new_n228), .A3(new_n229), .A4(new_n394), .ZN(new_n395));
  XNOR2_X1  g273(.A(G113), .B(G122), .ZN(new_n396));
  XNOR2_X1  g274(.A(new_n396), .B(new_n260), .ZN(new_n397));
  OAI211_X1 g275(.A(KEYINPUT18), .B(G131), .C1(new_n386), .C2(new_n387), .ZN(new_n398));
  NAND2_X1  g276(.A1(new_n222), .A2(new_n240), .ZN(new_n399));
  NAND2_X1  g277(.A1(new_n399), .A2(G146), .ZN(new_n400));
  NAND2_X1  g278(.A1(new_n400), .A2(new_n241), .ZN(new_n401));
  NAND2_X1  g279(.A1(KEYINPUT18), .A2(G131), .ZN(new_n402));
  NAND3_X1  g280(.A1(new_n390), .A2(new_n385), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g281(.A1(new_n398), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g282(.A1(new_n395), .A2(new_n397), .A3(new_n404), .ZN(new_n405));
  INV_X1    g283(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g284(.A(new_n397), .B1(new_n395), .B2(new_n404), .ZN(new_n407));
  OAI21_X1  g285(.A(new_n188), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g286(.A1(new_n408), .A2(G475), .ZN(new_n409));
  INV_X1    g287(.A(KEYINPUT20), .ZN(new_n410));
  NAND2_X1  g288(.A1(new_n388), .A2(new_n391), .ZN(new_n411));
  AND3_X1   g289(.A1(new_n222), .A2(new_n240), .A3(KEYINPUT19), .ZN(new_n412));
  AOI21_X1  g290(.A(KEYINPUT19), .B1(new_n222), .B2(new_n240), .ZN(new_n413));
  OAI21_X1  g291(.A(new_n133), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g292(.A1(new_n411), .A2(new_n414), .A3(new_n228), .ZN(new_n415));
  AND2_X1   g293(.A1(new_n415), .A2(new_n404), .ZN(new_n416));
  OAI21_X1  g294(.A(new_n405), .B1(new_n416), .B2(new_n397), .ZN(new_n417));
  NOR2_X1   g295(.A1(G475), .A2(G902), .ZN(new_n418));
  AOI21_X1  g296(.A(new_n410), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g297(.A1(new_n417), .A2(new_n410), .A3(new_n418), .ZN(new_n420));
  INV_X1    g298(.A(new_n420), .ZN(new_n421));
  OAI211_X1 g299(.A(new_n384), .B(new_n409), .C1(new_n419), .C2(new_n421), .ZN(new_n422));
  INV_X1    g300(.A(G952), .ZN(new_n423));
  AOI211_X1 g301(.A(G953), .B(new_n423), .C1(G234), .C2(G237), .ZN(new_n424));
  OR2_X1    g302(.A1(KEYINPUT21), .A2(G898), .ZN(new_n425));
  NAND2_X1  g303(.A1(KEYINPUT21), .A2(G898), .ZN(new_n426));
  AOI21_X1  g304(.A(new_n244), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g305(.A(new_n188), .B1(G234), .B2(G237), .ZN(new_n428));
  AOI21_X1  g306(.A(new_n424), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g307(.A1(new_n422), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g308(.A1(new_n218), .A2(new_n258), .A3(new_n352), .A4(new_n430), .ZN(new_n431));
  XNOR2_X1  g309(.A(new_n431), .B(G101), .ZN(G3));
  AND3_X1   g310(.A1(new_n212), .A2(new_n210), .A3(new_n215), .ZN(new_n433));
  AOI21_X1  g311(.A(new_n210), .B1(new_n212), .B2(new_n215), .ZN(new_n434));
  NOR3_X1   g312(.A1(new_n433), .A2(new_n434), .A3(new_n257), .ZN(new_n435));
  NAND2_X1  g313(.A1(new_n417), .A2(new_n418), .ZN(new_n436));
  NAND2_X1  g314(.A1(new_n436), .A2(KEYINPUT20), .ZN(new_n437));
  NAND2_X1  g315(.A1(new_n437), .A2(new_n420), .ZN(new_n438));
  AND2_X1   g316(.A1(new_n438), .A2(new_n409), .ZN(new_n439));
  NOR2_X1   g317(.A1(new_n353), .A2(new_n188), .ZN(new_n440));
  INV_X1    g318(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g319(.A1(new_n380), .A2(new_n353), .A3(new_n188), .ZN(new_n442));
  XNOR2_X1  g320(.A(new_n380), .B(KEYINPUT33), .ZN(new_n443));
  OAI211_X1 g321(.A(new_n441), .B(new_n442), .C1(new_n443), .C2(new_n353), .ZN(new_n444));
  NOR3_X1   g322(.A1(new_n439), .A2(new_n429), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g323(.A1(new_n352), .A2(new_n435), .A3(new_n445), .ZN(new_n446));
  XOR2_X1   g324(.A(KEYINPUT34), .B(G104), .Z(new_n447));
  XNOR2_X1  g325(.A(new_n446), .B(new_n447), .ZN(G6));
  OAI211_X1 g326(.A(new_n438), .B(new_n409), .C1(new_n383), .C2(new_n381), .ZN(new_n449));
  NOR2_X1   g327(.A1(new_n449), .A2(new_n429), .ZN(new_n450));
  NAND3_X1  g328(.A1(new_n352), .A2(new_n435), .A3(new_n450), .ZN(new_n451));
  XOR2_X1   g329(.A(KEYINPUT35), .B(G107), .Z(new_n452));
  XNOR2_X1  g330(.A(new_n451), .B(new_n452), .ZN(G9));
  NAND2_X1  g331(.A1(new_n212), .A2(new_n215), .ZN(new_n454));
  NAND2_X1  g332(.A1(new_n454), .A2(G472), .ZN(new_n455));
  NAND3_X1  g333(.A1(new_n212), .A2(new_n210), .A3(new_n215), .ZN(new_n456));
  NOR2_X1   g334(.A1(new_n248), .A2(KEYINPUT36), .ZN(new_n457));
  XNOR2_X1  g335(.A(new_n457), .B(new_n243), .ZN(new_n458));
  OAI211_X1 g336(.A(new_n458), .B(new_n188), .C1(new_n219), .C2(G234), .ZN(new_n459));
  NAND2_X1  g337(.A1(new_n255), .A2(new_n459), .ZN(new_n460));
  AND3_X1   g338(.A1(new_n455), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g339(.A1(new_n461), .A2(new_n352), .A3(new_n430), .ZN(new_n462));
  XOR2_X1   g340(.A(KEYINPUT37), .B(G110), .Z(new_n463));
  XNOR2_X1  g341(.A(new_n462), .B(new_n463), .ZN(G12));
  INV_X1    g342(.A(new_n424), .ZN(new_n465));
  INV_X1    g343(.A(G900), .ZN(new_n466));
  NAND3_X1  g344(.A1(new_n428), .A2(new_n466), .A3(G953), .ZN(new_n467));
  NAND2_X1  g345(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g346(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g347(.A1(new_n449), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g348(.A1(new_n218), .A2(new_n352), .A3(new_n460), .A4(new_n470), .ZN(new_n471));
  XNOR2_X1  g349(.A(new_n471), .B(G128), .ZN(G30));
  XNOR2_X1  g350(.A(new_n468), .B(KEYINPUT39), .ZN(new_n473));
  NAND3_X1  g351(.A1(new_n314), .A2(new_n316), .A3(new_n473), .ZN(new_n474));
  XOR2_X1   g352(.A(new_n474), .B(KEYINPUT40), .Z(new_n475));
  AOI21_X1  g353(.A(new_n170), .B1(new_n200), .B2(new_n162), .ZN(new_n476));
  AOI21_X1  g354(.A(new_n476), .B1(new_n207), .B2(new_n170), .ZN(new_n477));
  OAI21_X1  g355(.A(G472), .B1(new_n477), .B2(G902), .ZN(new_n478));
  OAI21_X1  g356(.A(new_n478), .B1(new_n211), .B2(new_n217), .ZN(new_n479));
  NOR2_X1   g357(.A1(new_n349), .A2(new_n350), .ZN(new_n480));
  XNOR2_X1  g358(.A(new_n480), .B(KEYINPUT38), .ZN(new_n481));
  INV_X1    g359(.A(new_n481), .ZN(new_n482));
  INV_X1    g360(.A(new_n318), .ZN(new_n483));
  NOR4_X1   g361(.A1(new_n439), .A2(new_n460), .A3(new_n384), .A4(new_n483), .ZN(new_n484));
  NAND4_X1  g362(.A1(new_n475), .A2(new_n479), .A3(new_n482), .A4(new_n484), .ZN(new_n485));
  XNOR2_X1  g363(.A(new_n485), .B(G143), .ZN(G45));
  NOR3_X1   g364(.A1(new_n439), .A2(new_n444), .A3(new_n469), .ZN(new_n487));
  NAND4_X1  g365(.A1(new_n218), .A2(new_n352), .A3(new_n460), .A4(new_n487), .ZN(new_n488));
  XNOR2_X1  g366(.A(new_n488), .B(G146), .ZN(G48));
  OAI21_X1  g367(.A(new_n188), .B1(new_n302), .B2(new_n306), .ZN(new_n490));
  NAND2_X1  g368(.A1(new_n490), .A2(G469), .ZN(new_n491));
  NAND3_X1  g369(.A1(new_n491), .A2(new_n316), .A3(new_n307), .ZN(new_n492));
  NOR2_X1   g370(.A1(new_n351), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g371(.A1(new_n218), .A2(new_n258), .A3(new_n445), .A4(new_n493), .ZN(new_n494));
  XNOR2_X1  g372(.A(KEYINPUT41), .B(G113), .ZN(new_n495));
  XNOR2_X1  g373(.A(new_n494), .B(new_n495), .ZN(G15));
  NAND4_X1  g374(.A1(new_n218), .A2(new_n258), .A3(new_n450), .A4(new_n493), .ZN(new_n497));
  XNOR2_X1  g375(.A(new_n497), .B(G116), .ZN(G18));
  NAND4_X1  g376(.A1(new_n218), .A2(new_n430), .A3(new_n460), .A4(new_n493), .ZN(new_n499));
  XNOR2_X1  g377(.A(new_n499), .B(G119), .ZN(G21));
  AOI21_X1  g378(.A(new_n384), .B1(new_n438), .B2(new_n409), .ZN(new_n501));
  OAI211_X1 g379(.A(new_n501), .B(new_n318), .C1(new_n350), .C2(new_n349), .ZN(new_n502));
  INV_X1    g380(.A(new_n502), .ZN(new_n503));
  INV_X1    g381(.A(new_n429), .ZN(new_n504));
  INV_X1    g382(.A(new_n492), .ZN(new_n505));
  NAND4_X1  g383(.A1(new_n503), .A2(new_n435), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  XNOR2_X1  g384(.A(new_n506), .B(G122), .ZN(G24));
  NAND3_X1  g385(.A1(new_n461), .A2(new_n493), .A3(new_n487), .ZN(new_n508));
  XNOR2_X1  g386(.A(new_n508), .B(G125), .ZN(G27));
  NAND2_X1  g387(.A1(new_n339), .A2(new_n348), .ZN(new_n510));
  INV_X1    g388(.A(new_n340), .ZN(new_n511));
  NAND2_X1  g389(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g390(.A1(new_n339), .A2(new_n340), .A3(new_n348), .ZN(new_n513));
  NAND3_X1  g391(.A1(new_n512), .A2(new_n318), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g392(.A1(new_n317), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g393(.A1(new_n218), .A2(new_n258), .A3(new_n515), .A4(new_n487), .ZN(new_n516));
  INV_X1    g394(.A(KEYINPUT42), .ZN(new_n517));
  NAND2_X1  g395(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g396(.A1(new_n456), .A2(KEYINPUT32), .ZN(new_n519));
  NAND2_X1  g397(.A1(new_n519), .A2(new_n216), .ZN(new_n520));
  AOI21_X1  g398(.A(new_n257), .B1(new_n520), .B2(new_n185), .ZN(new_n521));
  NAND4_X1  g399(.A1(new_n521), .A2(KEYINPUT42), .A3(new_n487), .A4(new_n515), .ZN(new_n522));
  NAND2_X1  g400(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g401(.A(new_n523), .B(G131), .ZN(G33));
  AND4_X1   g402(.A1(new_n218), .A2(new_n258), .A3(new_n470), .A4(new_n515), .ZN(new_n525));
  XNOR2_X1  g403(.A(new_n525), .B(new_n123), .ZN(G36));
  INV_X1    g404(.A(new_n444), .ZN(new_n527));
  INV_X1    g405(.A(KEYINPUT43), .ZN(new_n528));
  NAND3_X1  g406(.A1(new_n527), .A2(new_n439), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g407(.A1(new_n438), .A2(new_n409), .ZN(new_n530));
  OAI21_X1  g408(.A(KEYINPUT43), .B1(new_n444), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g409(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g410(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g411(.A1(new_n455), .A2(new_n456), .ZN(new_n534));
  NAND4_X1  g412(.A1(new_n533), .A2(KEYINPUT44), .A3(new_n534), .A4(new_n460), .ZN(new_n535));
  INV_X1    g413(.A(new_n514), .ZN(new_n536));
  INV_X1    g414(.A(KEYINPUT44), .ZN(new_n537));
  NAND2_X1  g415(.A1(new_n534), .A2(new_n460), .ZN(new_n538));
  OAI21_X1  g416(.A(new_n537), .B1(new_n538), .B2(new_n532), .ZN(new_n539));
  AND3_X1   g417(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  INV_X1    g418(.A(new_n316), .ZN(new_n541));
  INV_X1    g419(.A(new_n307), .ZN(new_n542));
  NAND2_X1  g420(.A1(new_n311), .A2(new_n312), .ZN(new_n543));
  NAND2_X1  g421(.A1(new_n543), .A2(KEYINPUT45), .ZN(new_n544));
  INV_X1    g422(.A(KEYINPUT45), .ZN(new_n545));
  NAND3_X1  g423(.A1(new_n311), .A2(new_n545), .A3(new_n312), .ZN(new_n546));
  NAND3_X1  g424(.A1(new_n544), .A2(new_n188), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g425(.A1(new_n547), .A2(G469), .ZN(new_n548));
  AOI21_X1  g426(.A(new_n542), .B1(new_n548), .B2(KEYINPUT46), .ZN(new_n549));
  INV_X1    g427(.A(KEYINPUT46), .ZN(new_n550));
  NAND3_X1  g428(.A1(new_n547), .A2(new_n550), .A3(G469), .ZN(new_n551));
  AOI21_X1  g429(.A(new_n541), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  AND2_X1   g430(.A1(new_n552), .A2(new_n473), .ZN(new_n553));
  NAND2_X1  g431(.A1(new_n540), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g432(.A(new_n554), .B(G137), .ZN(G39));
  XNOR2_X1  g433(.A(new_n552), .B(KEYINPUT47), .ZN(new_n556));
  NAND3_X1  g434(.A1(new_n487), .A2(new_n257), .A3(new_n536), .ZN(new_n557));
  NOR2_X1   g435(.A1(new_n557), .A2(new_n218), .ZN(new_n558));
  NAND2_X1  g436(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g437(.A(new_n559), .B(G140), .ZN(G42));
  INV_X1    g438(.A(KEYINPUT53), .ZN(new_n561));
  NAND3_X1  g439(.A1(new_n314), .A2(new_n316), .A3(new_n468), .ZN(new_n562));
  NOR2_X1   g440(.A1(new_n562), .A2(new_n460), .ZN(new_n563));
  NAND3_X1  g441(.A1(new_n479), .A2(new_n503), .A3(new_n563), .ZN(new_n564));
  NAND4_X1  g442(.A1(new_n471), .A2(new_n488), .A3(new_n508), .A4(new_n564), .ZN(new_n565));
  XNOR2_X1  g443(.A(new_n565), .B(KEYINPUT52), .ZN(new_n566));
  AOI21_X1  g444(.A(new_n525), .B1(new_n518), .B2(new_n522), .ZN(new_n567));
  AND4_X1   g445(.A1(new_n431), .A2(new_n494), .A3(new_n497), .A4(new_n446), .ZN(new_n568));
  AND4_X1   g446(.A1(new_n451), .A2(new_n499), .A3(new_n462), .A4(new_n506), .ZN(new_n569));
  NOR3_X1   g447(.A1(new_n562), .A2(new_n514), .A3(new_n422), .ZN(new_n570));
  NAND3_X1  g448(.A1(new_n570), .A2(new_n218), .A3(new_n460), .ZN(new_n571));
  NAND3_X1  g449(.A1(new_n461), .A2(new_n515), .A3(new_n487), .ZN(new_n572));
  AND2_X1   g450(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g451(.A1(new_n567), .A2(new_n568), .A3(new_n569), .A4(new_n573), .ZN(new_n574));
  OAI21_X1  g452(.A(new_n561), .B1(new_n566), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g453(.A1(new_n471), .A2(new_n508), .ZN(new_n576));
  NAND4_X1  g454(.A1(new_n576), .A2(KEYINPUT52), .A3(new_n488), .A4(new_n564), .ZN(new_n577));
  INV_X1    g455(.A(KEYINPUT52), .ZN(new_n578));
  NAND2_X1  g456(.A1(new_n565), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g457(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g458(.A(new_n525), .ZN(new_n581));
  AND3_X1   g459(.A1(new_n523), .A2(new_n581), .A3(new_n573), .ZN(new_n582));
  NAND4_X1  g460(.A1(new_n431), .A2(new_n494), .A3(new_n497), .A4(new_n446), .ZN(new_n583));
  NAND4_X1  g461(.A1(new_n499), .A2(new_n506), .A3(new_n451), .A4(new_n462), .ZN(new_n584));
  NOR2_X1   g462(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g463(.A1(new_n580), .A2(new_n582), .A3(KEYINPUT53), .A4(new_n585), .ZN(new_n586));
  AND3_X1   g464(.A1(new_n575), .A2(KEYINPUT54), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g465(.A(KEYINPUT54), .B1(new_n575), .B2(new_n586), .ZN(new_n588));
  NOR2_X1   g466(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g467(.A(new_n479), .ZN(new_n590));
  NOR2_X1   g468(.A1(new_n514), .A2(new_n492), .ZN(new_n591));
  NAND4_X1  g469(.A1(new_n590), .A2(new_n258), .A3(new_n424), .A4(new_n591), .ZN(new_n592));
  OR3_X1    g470(.A1(new_n592), .A2(new_n530), .A3(new_n527), .ZN(new_n593));
  NOR2_X1   g471(.A1(new_n532), .A2(new_n465), .ZN(new_n594));
  NAND3_X1  g472(.A1(new_n594), .A2(new_n461), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g473(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g474(.A1(new_n594), .A2(new_n435), .A3(new_n505), .ZN(new_n597));
  INV_X1    g475(.A(KEYINPUT50), .ZN(new_n598));
  NAND2_X1  g476(.A1(new_n481), .A2(new_n483), .ZN(new_n599));
  OR3_X1    g477(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g478(.A(new_n598), .B1(new_n597), .B2(new_n599), .ZN(new_n601));
  AOI21_X1  g479(.A(new_n596), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g480(.A1(new_n491), .A2(new_n307), .ZN(new_n603));
  INV_X1    g481(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g482(.A(new_n556), .B1(new_n541), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g483(.A1(new_n594), .A2(new_n435), .A3(new_n536), .ZN(new_n606));
  OAI211_X1 g484(.A(new_n602), .B(KEYINPUT51), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  INV_X1    g485(.A(KEYINPUT51), .ZN(new_n608));
  NOR2_X1   g486(.A1(new_n605), .A2(new_n606), .ZN(new_n609));
  NAND2_X1  g487(.A1(new_n600), .A2(new_n601), .ZN(new_n610));
  NAND3_X1  g488(.A1(new_n610), .A2(new_n595), .A3(new_n593), .ZN(new_n611));
  OAI21_X1  g489(.A(new_n608), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g490(.A1(new_n439), .A2(new_n444), .ZN(new_n613));
  INV_X1    g491(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g492(.A1(new_n592), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g493(.A1(new_n594), .A2(new_n521), .A3(new_n591), .ZN(new_n616));
  INV_X1    g494(.A(KEYINPUT48), .ZN(new_n617));
  OAI22_X1  g495(.A1(new_n597), .A2(new_n351), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI211_X1 g496(.A(new_n615), .B(new_n618), .C1(new_n617), .C2(new_n616), .ZN(new_n619));
  NAND3_X1  g497(.A1(new_n607), .A2(new_n612), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g498(.A(G952), .B1(new_n589), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g499(.A(new_n603), .B(KEYINPUT49), .ZN(new_n622));
  NAND2_X1  g500(.A1(new_n527), .A2(new_n439), .ZN(new_n623));
  NAND3_X1  g501(.A1(new_n258), .A2(new_n318), .A3(new_n316), .ZN(new_n624));
  NOR4_X1   g502(.A1(new_n482), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  AOI21_X1  g503(.A(G953), .B1(new_n625), .B2(new_n590), .ZN(new_n626));
  NAND2_X1  g504(.A1(new_n621), .A2(new_n626), .ZN(G75));
  NAND2_X1  g505(.A1(new_n575), .A2(new_n586), .ZN(new_n628));
  NOR2_X1   g506(.A1(new_n340), .A2(new_n188), .ZN(new_n629));
  AOI21_X1  g507(.A(KEYINPUT56), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g508(.A1(new_n336), .A2(new_n338), .ZN(new_n631));
  XNOR2_X1  g509(.A(new_n631), .B(new_n324), .ZN(new_n632));
  XOR2_X1   g510(.A(new_n632), .B(KEYINPUT55), .Z(new_n633));
  INV_X1    g511(.A(new_n633), .ZN(new_n634));
  AND2_X1   g512(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g513(.A1(new_n630), .A2(new_n634), .ZN(new_n636));
  NOR2_X1   g514(.A1(new_n244), .A2(G952), .ZN(new_n637));
  NOR3_X1   g515(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(G51));
  INV_X1    g516(.A(KEYINPUT54), .ZN(new_n639));
  NAND2_X1  g517(.A1(new_n628), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g518(.A1(new_n575), .A2(new_n586), .A3(KEYINPUT54), .ZN(new_n641));
  XNOR2_X1  g519(.A(new_n308), .B(KEYINPUT57), .ZN(new_n642));
  NAND3_X1  g520(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  OR2_X1    g521(.A1(new_n302), .A2(new_n306), .ZN(new_n644));
  NAND2_X1  g522(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g523(.A(new_n309), .B1(new_n544), .B2(new_n546), .ZN(new_n646));
  NAND2_X1  g524(.A1(new_n628), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g525(.A(new_n637), .B1(new_n645), .B2(new_n647), .ZN(G54));
  AND3_X1   g526(.A1(KEYINPUT58), .A2(G475), .A3(G902), .ZN(new_n649));
  AND3_X1   g527(.A1(new_n628), .A2(new_n417), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g528(.A(new_n417), .B1(new_n628), .B2(new_n649), .ZN(new_n651));
  NOR3_X1   g529(.A1(new_n650), .A2(new_n651), .A3(new_n637), .ZN(G60));
  XOR2_X1   g530(.A(new_n440), .B(KEYINPUT59), .Z(new_n653));
  AOI21_X1  g531(.A(new_n443), .B1(new_n589), .B2(new_n653), .ZN(new_n654));
  NAND4_X1  g532(.A1(new_n640), .A2(new_n443), .A3(new_n641), .A4(new_n653), .ZN(new_n655));
  INV_X1    g533(.A(new_n637), .ZN(new_n656));
  NAND2_X1  g534(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g535(.A1(new_n654), .A2(new_n657), .ZN(G63));
  INV_X1    g536(.A(KEYINPUT61), .ZN(new_n659));
  NAND2_X1  g537(.A1(G217), .A2(G902), .ZN(new_n660));
  XOR2_X1   g538(.A(new_n660), .B(KEYINPUT60), .Z(new_n661));
  INV_X1    g539(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g540(.A(new_n662), .B1(new_n575), .B2(new_n586), .ZN(new_n663));
  NAND2_X1  g541(.A1(new_n663), .A2(new_n458), .ZN(new_n664));
  INV_X1    g542(.A(new_n664), .ZN(new_n665));
  AND2_X1   g543(.A1(new_n249), .A2(new_n250), .ZN(new_n666));
  OAI21_X1  g544(.A(new_n656), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g545(.A(new_n659), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  OR2_X1    g546(.A1(new_n663), .A2(new_n666), .ZN(new_n669));
  NAND4_X1  g547(.A1(new_n669), .A2(KEYINPUT61), .A3(new_n656), .A4(new_n664), .ZN(new_n670));
  NAND2_X1  g548(.A1(new_n668), .A2(new_n670), .ZN(G66));
  AOI21_X1  g549(.A(new_n427), .B1(new_n322), .B2(G953), .ZN(new_n672));
  OAI21_X1  g550(.A(new_n672), .B1(new_n585), .B2(G953), .ZN(new_n673));
  OAI21_X1  g551(.A(new_n631), .B1(G898), .B2(new_n244), .ZN(new_n674));
  XNOR2_X1  g552(.A(new_n673), .B(new_n674), .ZN(G69));
  NAND2_X1  g553(.A1(new_n559), .A2(new_n554), .ZN(new_n676));
  NAND3_X1  g554(.A1(new_n553), .A2(new_n521), .A3(new_n503), .ZN(new_n677));
  NAND4_X1  g555(.A1(new_n677), .A2(new_n488), .A3(new_n576), .A4(new_n567), .ZN(new_n678));
  NOR2_X1   g556(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g557(.A1(new_n679), .A2(G953), .ZN(new_n680));
  OR2_X1    g558(.A1(new_n412), .A2(new_n413), .ZN(new_n681));
  XNOR2_X1  g559(.A(new_n206), .B(new_n681), .ZN(new_n682));
  OAI21_X1  g560(.A(new_n682), .B1(G900), .B2(new_n244), .ZN(new_n683));
  NOR2_X1   g561(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  AOI22_X1  g562(.A1(new_n556), .A2(new_n558), .B1(new_n540), .B2(new_n553), .ZN(new_n685));
  NAND3_X1  g563(.A1(new_n485), .A2(new_n576), .A3(new_n488), .ZN(new_n686));
  NAND2_X1  g564(.A1(new_n686), .A2(KEYINPUT62), .ZN(new_n687));
  INV_X1    g565(.A(KEYINPUT62), .ZN(new_n688));
  NAND4_X1  g566(.A1(new_n485), .A2(new_n576), .A3(new_n688), .A4(new_n488), .ZN(new_n689));
  AOI21_X1  g567(.A(new_n474), .B1(new_n614), .B2(new_n449), .ZN(new_n690));
  NAND3_X1  g568(.A1(new_n690), .A2(new_n521), .A3(new_n536), .ZN(new_n691));
  AND4_X1   g569(.A1(new_n685), .A2(new_n687), .A3(new_n689), .A4(new_n691), .ZN(new_n692));
  OR2_X1    g570(.A1(new_n682), .A2(G953), .ZN(new_n693));
  NOR2_X1   g571(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g572(.A(G953), .B1(new_n296), .B2(new_n466), .ZN(new_n695));
  OR3_X1    g573(.A1(new_n684), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g574(.A(new_n695), .B1(new_n684), .B2(new_n694), .ZN(new_n697));
  NAND2_X1  g575(.A1(new_n696), .A2(new_n697), .ZN(G72));
  NAND2_X1  g576(.A1(G472), .A2(G902), .ZN(new_n699));
  XNOR2_X1  g577(.A(new_n699), .B(KEYINPUT63), .ZN(new_n700));
  INV_X1    g578(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g579(.A1(new_n628), .A2(new_n207), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g580(.A(new_n700), .B1(new_n692), .B2(new_n585), .ZN(new_n703));
  OAI211_X1 g581(.A(new_n170), .B(new_n702), .C1(new_n703), .C2(new_n207), .ZN(new_n704));
  NAND3_X1  g582(.A1(new_n628), .A2(new_n181), .A3(new_n701), .ZN(new_n705));
  AOI21_X1  g583(.A(new_n700), .B1(new_n679), .B2(new_n585), .ZN(new_n706));
  OAI211_X1 g584(.A(new_n705), .B(new_n182), .C1(new_n181), .C2(new_n706), .ZN(new_n707));
  AOI21_X1  g585(.A(new_n637), .B1(new_n704), .B2(new_n707), .ZN(G57));
endmodule


