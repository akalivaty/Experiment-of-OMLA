//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XOR2_X1   g020(.A(KEYINPUT64), .B(KEYINPUT1), .Z(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT65), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n463), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT66), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT66), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI211_X1 g049(.A(new_n469), .B(new_n471), .C1(G2105), .C2(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n463), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n482), .B1(G136), .B2(new_n484), .ZN(G162));
  NAND2_X1  g060(.A1(G126), .A2(G2105), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(new_n476), .B2(new_n477), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n463), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT67), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n494));
  INV_X1    g069(.A(new_n486), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n464), .B2(new_n465), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(KEYINPUT68), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(new_n463), .C1(new_n465), .C2(new_n464), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n476), .A2(new_n477), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n502), .A2(new_n503), .A3(new_n463), .A4(new_n499), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n491), .A2(new_n497), .B1(new_n501), .B2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT69), .A3(G543), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n509), .A2(new_n511), .B1(KEYINPUT5), .B2(new_n508), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n512), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n506), .A2(new_n513), .B1(new_n514), .B2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND2_X1  g095(.A1(new_n517), .A2(KEYINPUT70), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n515), .A2(new_n522), .A3(new_n516), .ZN(new_n523));
  AND3_X1   g098(.A1(new_n521), .A2(G543), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT71), .B(G51), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT72), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n517), .A2(G89), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n512), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n526), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(G168));
  AOI21_X1  g109(.A(new_n508), .B1(new_n517), .B2(KEYINPUT70), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(new_n523), .ZN(new_n536));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n512), .A2(new_n517), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n536), .A2(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n506), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n509), .A2(new_n511), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  XNOR2_X1  g125(.A(KEYINPUT73), .B(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n524), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n547), .A2(new_n518), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G81), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n550), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(KEYINPUT74), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(KEYINPUT74), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  AOI22_X1  g138(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G91), .ZN(new_n565));
  OAI22_X1  g140(.A1(new_n564), .A2(new_n506), .B1(new_n565), .B2(new_n538), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  AND2_X1   g142(.A1(KEYINPUT75), .A2(G53), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n535), .A2(new_n523), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n535), .A2(new_n572), .A3(new_n523), .A4(new_n568), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n571), .B1(new_n570), .B2(new_n573), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n567), .B1(new_n574), .B2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n533), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n526), .A2(new_n529), .A3(KEYINPUT77), .A4(new_n532), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G286));
  NAND4_X1  g157(.A1(new_n521), .A2(G49), .A3(G543), .A4(new_n523), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n512), .A2(G87), .A3(new_n517), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  AOI22_X1  g161(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n506), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n512), .A2(G86), .ZN(new_n589));
  NAND2_X1  g164(.A1(G48), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n518), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n506), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(KEYINPUT78), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(KEYINPUT78), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n524), .A2(G47), .B1(new_n553), .B2(G85), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G290));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NOR2_X1   g175(.A1(G301), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n553), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n538), .B2(new_n604), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n524), .A2(G54), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n506), .B2(new_n608), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(KEYINPUT79), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n606), .A2(new_n609), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT79), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n601), .B1(new_n615), .B2(new_n600), .ZN(G284));
  AOI21_X1  g191(.A(new_n601), .B1(new_n615), .B2(new_n600), .ZN(G321));
  MUX2_X1   g192(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g193(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n615), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n556), .A2(new_n557), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(new_n600), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n615), .A2(new_n620), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n615), .A2(KEYINPUT80), .A3(new_n620), .ZN(new_n627));
  AND2_X1   g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n623), .B1(new_n628), .B2(new_n600), .ZN(G323));
  XNOR2_X1  g204(.A(KEYINPUT81), .B(KEYINPUT11), .ZN(new_n630));
  XNOR2_X1  g205(.A(G323), .B(new_n630), .ZN(G282));
  NAND2_X1  g206(.A1(new_n502), .A2(new_n467), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT12), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT12), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n502), .A2(new_n634), .A3(new_n467), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT82), .Z(new_n640));
  AOI22_X1  g215(.A1(new_n484), .A2(G135), .B1(new_n478), .B2(G123), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT83), .ZN(new_n643));
  INV_X1    g218(.A(G111), .ZN(new_n644));
  AOI22_X1  g219(.A1(new_n642), .A2(new_n643), .B1(new_n644), .B2(G2105), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n643), .B2(new_n642), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(G2096), .Z(new_n648));
  OAI211_X1 g223(.A(new_n640), .B(new_n648), .C1(new_n638), .C2(new_n637), .ZN(G156));
  INV_X1    g224(.A(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n655), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(G14), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n661), .ZN(G401));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n666), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT84), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2100), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT18), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n667), .A2(new_n668), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2096), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n672), .B(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n687));
  INV_X1    g262(.A(new_n684), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n682), .A2(new_n683), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n686), .B(new_n687), .C1(new_n681), .C2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n693), .B(new_n694), .Z(new_n695));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n693), .B(new_n694), .ZN(new_n699));
  INV_X1    g274(.A(new_n696), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AND3_X1   g276(.A1(new_n697), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n698), .B1(new_n697), .B2(new_n701), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(G229));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NOR2_X1   g280(.A1(G168), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n705), .B2(G21), .ZN(new_n707));
  INV_X1    g282(.A(G1966), .ZN(new_n708));
  INV_X1    g283(.A(G2084), .ZN(new_n709));
  NAND2_X1  g284(.A1(G160), .A2(G29), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT87), .B(G29), .Z(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT24), .B(G34), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT94), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n707), .A2(new_n708), .B1(new_n709), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(G5), .A2(G16), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT98), .Z(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G171), .B2(G16), .ZN(new_n720));
  OAI221_X1 g295(.A(new_n716), .B1(G1961), .B2(new_n720), .C1(new_n709), .C2(new_n715), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT31), .B(G11), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT97), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT30), .B(G28), .Z(new_n724));
  OAI221_X1 g299(.A(new_n723), .B1(G29), .B2(new_n724), .C1(new_n647), .C2(new_n711), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT25), .ZN(new_n726));
  NAND2_X1  g301(.A1(G103), .A2(G2104), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(G2105), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n484), .A2(G139), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n502), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n463), .B2(new_n731), .ZN(new_n732));
  MUX2_X1   g307(.A(G33), .B(new_n732), .S(G29), .Z(new_n733));
  AOI21_X1  g308(.A(new_n725), .B1(new_n733), .B2(G2072), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n720), .A2(G1961), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n734), .B(new_n735), .C1(G2072), .C2(new_n733), .ZN(new_n736));
  INV_X1    g311(.A(new_n711), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(G27), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G164), .B2(new_n737), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(G2078), .Z(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n707), .B2(new_n708), .ZN(new_n741));
  NOR3_X1   g316(.A1(new_n721), .A2(new_n736), .A3(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT95), .B(KEYINPUT26), .Z(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n467), .A2(G105), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n484), .A2(G141), .B1(new_n478), .B2(G129), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT96), .ZN(new_n749));
  MUX2_X1   g324(.A(G32), .B(new_n749), .S(G29), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT27), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1996), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n742), .A2(new_n752), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(KEYINPUT99), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n705), .A2(G22), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G166), .B2(new_n705), .ZN(new_n756));
  INV_X1    g331(.A(G1971), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G6), .A2(G16), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n592), .B2(G16), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT32), .B(G1981), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n705), .A2(G23), .ZN(new_n763));
  AND3_X1   g338(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n705), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT33), .B(G1976), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n758), .A2(new_n762), .A3(new_n767), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(KEYINPUT34), .ZN(new_n769));
  NAND2_X1  g344(.A1(G290), .A2(G16), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n705), .A2(G24), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(KEYINPUT88), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(KEYINPUT88), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(G1986), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n737), .A2(G25), .ZN(new_n776));
  OR2_X1    g351(.A1(G95), .A2(G2105), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n777), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n778));
  INV_X1    g353(.A(G131), .ZN(new_n779));
  INV_X1    g354(.A(new_n478), .ZN(new_n780));
  INV_X1    g355(.A(G119), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n778), .B1(new_n483), .B2(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n776), .B1(new_n783), .B2(new_n737), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT35), .B(G1991), .Z(new_n785));
  XOR2_X1   g360(.A(new_n784), .B(new_n785), .Z(new_n786));
  NOR2_X1   g361(.A1(new_n775), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n768), .A2(KEYINPUT34), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n774), .A2(G1986), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n769), .A2(new_n787), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT36), .ZN(new_n791));
  INV_X1    g366(.A(G19), .ZN(new_n792));
  OR3_X1    g367(.A1(new_n792), .A2(KEYINPUT90), .A3(G16), .ZN(new_n793));
  OAI21_X1  g368(.A(KEYINPUT90), .B1(new_n792), .B2(G16), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n793), .B(new_n794), .C1(new_n558), .C2(new_n705), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1341), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n705), .A2(G4), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n615), .B2(new_n705), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT89), .B(G1348), .Z(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n796), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n737), .A2(G35), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G162), .B2(new_n737), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT29), .Z(new_n805));
  INV_X1    g380(.A(G2090), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT100), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n711), .A2(G26), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT28), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n484), .A2(G140), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT91), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n813));
  INV_X1    g388(.A(G116), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G2105), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(KEYINPUT92), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(KEYINPUT92), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n816), .A2(new_n817), .B1(G128), .B2(new_n478), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n812), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n810), .B1(new_n819), .B2(G29), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT93), .B(G2067), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n808), .B(new_n822), .C1(new_n806), .C2(new_n805), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n705), .A2(G20), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT23), .ZN(new_n825));
  INV_X1    g400(.A(G299), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n705), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1956), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n798), .A2(new_n800), .ZN(new_n829));
  NOR4_X1   g404(.A1(new_n802), .A2(new_n823), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n753), .A2(KEYINPUT99), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n754), .A2(new_n791), .A3(new_n830), .A4(new_n831), .ZN(G150));
  INV_X1    g407(.A(G150), .ZN(G311));
  AOI22_X1  g408(.A1(new_n524), .A2(G55), .B1(new_n553), .B2(G93), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(KEYINPUT101), .ZN(new_n836));
  OAI21_X1  g411(.A(G651), .B1(new_n835), .B2(KEYINPUT101), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(KEYINPUT102), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(KEYINPUT102), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n615), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n839), .A2(new_n555), .A3(new_n840), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n556), .A2(new_n557), .A3(new_n838), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n845), .B(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n850));
  INV_X1    g425(.A(G860), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n849), .B2(KEYINPUT39), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n843), .B1(new_n850), .B2(new_n852), .ZN(G145));
  XNOR2_X1  g428(.A(new_n782), .B(new_n636), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n484), .A2(G142), .ZN(new_n855));
  OAI21_X1  g430(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT104), .ZN(new_n857));
  INV_X1    g432(.A(G118), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n856), .A2(new_n857), .B1(new_n858), .B2(G2105), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n857), .B2(new_n856), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n478), .A2(G130), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n855), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n854), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n749), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n819), .B(new_n732), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n501), .A2(new_n504), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n493), .A2(new_n496), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n866), .A2(KEYINPUT103), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT103), .B1(new_n866), .B2(new_n868), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n865), .B(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(G160), .B(new_n647), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(G162), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n864), .A2(new_n872), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n873), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n864), .B(new_n872), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n875), .ZN(new_n880));
  INV_X1    g455(.A(G37), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g458(.A1(new_n628), .A2(new_n848), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n626), .A2(new_n627), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(new_n847), .A3(new_n846), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n610), .A2(G299), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n610), .A2(G299), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(G290), .B(G305), .ZN(new_n894));
  XNOR2_X1  g469(.A(G303), .B(new_n764), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n894), .B(new_n895), .Z(new_n896));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT42), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n897), .A2(KEYINPUT42), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n894), .B(new_n895), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n901), .A2(new_n897), .A3(KEYINPUT42), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n890), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(new_n905), .A3(new_n888), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT41), .B1(new_n889), .B2(new_n890), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT105), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n891), .A2(new_n909), .A3(new_n905), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n884), .A2(new_n886), .A3(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n893), .A2(new_n903), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n903), .B1(new_n893), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n841), .A2(new_n600), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(G295));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n916), .ZN(G331));
  NOR2_X1   g493(.A1(G168), .A2(G171), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n919), .B1(G171), .B2(new_n581), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n848), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n920), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(new_n847), .A3(new_n846), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n908), .A3(new_n910), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(new_n923), .A3(new_n891), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n896), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n881), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n896), .B1(new_n925), .B2(new_n926), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT43), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n921), .A2(new_n923), .A3(new_n931), .A4(new_n891), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n926), .A2(KEYINPUT108), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n921), .A2(new_n923), .B1(new_n906), .B2(new_n907), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n901), .B(new_n932), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n935), .A2(new_n936), .A3(new_n881), .A4(new_n927), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n930), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n929), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n941), .A2(new_n936), .A3(new_n881), .A4(new_n927), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n935), .A2(new_n881), .A3(new_n927), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n942), .B(KEYINPUT44), .C1(new_n943), .C2(new_n936), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n940), .A2(new_n944), .ZN(G397));
  INV_X1    g520(.A(new_n870), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n867), .B1(new_n501), .B2(new_n504), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT103), .ZN(new_n948));
  INV_X1    g523(.A(G1384), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G40), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n953), .B1(new_n474), .B2(G2105), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n466), .A2(new_n468), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT66), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n957), .A3(new_n470), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n952), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G2067), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n819), .B(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n749), .A2(G1996), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n749), .A2(G1996), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n783), .A2(new_n785), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n783), .A2(new_n785), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(G290), .B(G1986), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n959), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n491), .A2(new_n497), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n866), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n951), .A2(G1384), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n958), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n951), .B1(new_n947), .B2(G1384), .ZN(new_n975));
  AOI21_X1  g550(.A(G1966), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n866), .A2(new_n868), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n979), .A3(new_n949), .ZN(new_n980));
  AND4_X1   g555(.A1(new_n709), .A2(new_n954), .A3(new_n957), .A4(new_n470), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n977), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(KEYINPUT120), .B(G8), .C1(new_n976), .C2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n984));
  INV_X1    g559(.A(G8), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(G168), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n471), .A2(new_n469), .ZN(new_n989));
  INV_X1    g564(.A(new_n973), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n989), .B(new_n954), .C1(G164), .C2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT45), .B1(new_n978), .B2(new_n949), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n708), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n977), .A2(new_n980), .A3(new_n981), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n985), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(KEYINPUT120), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT121), .B1(new_n988), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n993), .A2(new_n994), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(G8), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT120), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n986), .B1(new_n995), .B2(KEYINPUT120), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT121), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(G168), .A2(new_n985), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT51), .B1(new_n995), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n997), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT62), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n998), .A2(new_n1005), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT126), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n764), .A2(new_n1012), .A3(G1976), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n989), .A2(new_n978), .A3(new_n949), .A4(new_n954), .ZN(new_n1014));
  INV_X1    g589(.A(G1976), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT111), .B1(G288), .B2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .A4(G8), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT113), .B(G1976), .Z(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(G288), .B2(new_n1019), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n1020), .A2(KEYINPUT114), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(KEYINPUT114), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT49), .ZN(new_n1024));
  OAI21_X1  g599(.A(G1981), .B1(new_n588), .B2(new_n591), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n588), .A2(new_n591), .A3(G1981), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1024), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1027), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(KEYINPUT49), .A3(new_n1025), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1014), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(new_n985), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1017), .A2(new_n1034), .A3(KEYINPUT52), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1034), .B1(new_n1017), .B2(KEYINPUT52), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1023), .B(new_n1033), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT109), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(G166), .B2(new_n985), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT109), .ZN(new_n1042));
  NAND4_X1  g617(.A1(G303), .A2(new_n1042), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n978), .A2(new_n949), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n958), .B1(new_n1045), .B2(KEYINPUT50), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1384), .B1(new_n971), .B2(new_n866), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(new_n979), .ZN(new_n1049));
  NOR4_X1   g624(.A1(G164), .A2(KEYINPUT115), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1046), .B(new_n806), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n869), .A2(new_n870), .A3(new_n990), .ZN(new_n1052));
  INV_X1    g627(.A(new_n958), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n1048), .B2(KEYINPUT45), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n757), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1044), .B1(new_n1056), .B2(G8), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1037), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n972), .A2(new_n949), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n958), .B1(new_n1059), .B2(new_n951), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n946), .A2(new_n948), .A3(new_n973), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1971), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n977), .A2(new_n1053), .A3(new_n980), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(G2090), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1044), .B(G8), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT110), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1055), .B1(G2090), .B2(new_n1063), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1068), .A2(KEYINPUT110), .A3(G8), .A4(new_n1044), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1071), .B1(new_n1072), .B2(G2078), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n991), .A2(new_n992), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1071), .A2(G2078), .ZN(new_n1075));
  XOR2_X1   g650(.A(KEYINPUT123), .B(G1961), .Z(new_n1076));
  AOI22_X1  g651(.A1(new_n1074), .A2(new_n1075), .B1(new_n1063), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(G301), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1058), .A2(new_n1070), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1010), .A2(new_n1011), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT62), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1011), .B1(new_n1010), .B2(new_n1079), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n995), .A2(new_n581), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1068), .A2(G8), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(new_n1044), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT63), .B1(new_n1089), .B2(new_n1037), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1033), .A2(new_n1015), .A3(new_n764), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1032), .B1(new_n1091), .B2(new_n1027), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  OR3_X1    g668(.A1(new_n1057), .A2(KEYINPUT63), .A3(new_n1086), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1037), .B1(new_n1094), .B2(new_n1070), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1097));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n463), .B1(new_n474), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1098), .B2(new_n474), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1100), .A2(new_n989), .A3(G40), .A4(new_n1075), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1052), .A2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1102), .A2(new_n952), .B1(new_n1063), .B2(new_n1076), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1103), .A2(new_n1073), .A3(G301), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1097), .B1(new_n1104), .B2(new_n1078), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(KEYINPUT125), .B(new_n1097), .C1(new_n1104), .C2(new_n1078), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1073), .A2(G301), .A3(new_n1077), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1103), .A2(new_n1073), .ZN(new_n1111));
  OAI211_X1 g686(.A(KEYINPUT54), .B(new_n1110), .C1(new_n1111), .C2(G301), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1112), .A2(new_n1070), .A3(new_n1058), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(new_n1113), .A3(new_n1081), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n570), .A2(new_n573), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1115), .A2(KEYINPUT57), .A3(new_n566), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1046), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1118));
  INV_X1    g693(.A(G1956), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1117), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1063), .A2(new_n799), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1031), .A2(new_n960), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1124), .B1(new_n615), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1117), .A2(new_n1120), .A3(new_n1123), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(KEYINPUT61), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1117), .A2(new_n1120), .A3(new_n1123), .A4(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n1136));
  INV_X1    g711(.A(G1996), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1060), .A2(new_n1137), .A3(new_n1061), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT116), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1140), .B(G1341), .Z(new_n1141));
  AOI22_X1  g716(.A1(new_n1138), .A2(new_n1139), .B1(new_n1014), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1121), .A2(KEYINPUT116), .A3(new_n1137), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1136), .B1(new_n1144), .B2(new_n558), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1136), .ZN(new_n1146));
  AOI211_X1 g721(.A(new_n622), .B(new_n1146), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1135), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT60), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1127), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT119), .B1(new_n611), .B2(new_n614), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n1152), .A2(new_n1153), .B1(new_n1154), .B2(new_n615), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1127), .A2(new_n1149), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1131), .B1(new_n1148), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1096), .B1(new_n1114), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n970), .B1(new_n1085), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(G290), .A2(G1986), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT48), .B1(new_n1161), .B2(new_n959), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1161), .A2(KEYINPUT48), .A3(new_n959), .ZN(new_n1163));
  AOI211_X1 g738(.A(new_n1162), .B(new_n1163), .C1(new_n968), .C2(new_n959), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n959), .B1(new_n962), .B2(new_n749), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n959), .A2(new_n1137), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1166), .A2(KEYINPUT46), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1166), .A2(KEYINPUT46), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1165), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT47), .Z(new_n1170));
  XOR2_X1   g745(.A(new_n966), .B(KEYINPUT127), .Z(new_n1171));
  NAND2_X1  g746(.A1(new_n965), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(G2067), .B2(new_n819), .ZN(new_n1173));
  AOI211_X1 g748(.A(new_n1164), .B(new_n1170), .C1(new_n959), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1160), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g750(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1177));
  OAI211_X1 g751(.A(new_n882), .B(new_n1177), .C1(new_n702), .C2(new_n703), .ZN(new_n1178));
  AOI21_X1  g752(.A(new_n1178), .B1(new_n930), .B2(new_n937), .ZN(G308));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1180));
  NAND2_X1  g754(.A1(new_n1180), .A2(new_n938), .ZN(G225));
endmodule


