//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT5), .ZN(new_n203));
  XOR2_X1   g002(.A(G127gat), .B(G134gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT69), .ZN(new_n205));
  INV_X1    g004(.A(G113gat), .ZN(new_n206));
  INV_X1    g005(.A(G120gat), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT1), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(new_n206), .B2(new_n207), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT70), .B(G120gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n204), .B1(G113gat), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(new_n208), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G141gat), .B(G148gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n217), .B1(G155gat), .B2(G162gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  OAI22_X1  g018(.A1(new_n216), .A2(new_n218), .B1(KEYINPUT77), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G155gat), .B(G162gat), .Z(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n222), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT3), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n215), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT4), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n214), .A2(new_n222), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n228), .B1(new_n214), .B2(new_n222), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n227), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G225gat), .A2(G233gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n203), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT78), .B1(new_n214), .B2(new_n222), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(new_n222), .B2(new_n214), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n215), .A2(new_n225), .A3(KEYINPUT78), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n234), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n231), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n229), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n241), .A2(KEYINPUT5), .A3(new_n233), .A4(new_n227), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n235), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G1gat), .B(G29gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT0), .ZN(new_n245));
  INV_X1    g044(.A(G57gat), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n246), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G85gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n249), .A2(new_n250), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT6), .B1(new_n243), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n243), .A2(new_n254), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n255), .B(new_n256), .Z(new_n257));
  INV_X1    g056(.A(KEYINPUT76), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT75), .ZN(new_n259));
  AND2_X1   g058(.A1(G211gat), .A2(G218gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(G211gat), .A2(G218gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G211gat), .ZN(new_n263));
  INV_X1    g062(.A(G218gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G211gat), .A2(G218gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(KEYINPUT75), .A3(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT74), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n269), .B1(new_n260), .B2(KEYINPUT22), .ZN(new_n270));
  XNOR2_X1  g069(.A(G197gat), .B(G204gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT22), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n266), .A2(KEYINPUT74), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n258), .B1(new_n268), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n273), .ZN(new_n276));
  AND2_X1   g075(.A1(G197gat), .A2(G204gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(G197gat), .A2(G204gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT74), .B1(new_n266), .B2(new_n272), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n276), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n262), .A2(new_n267), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(KEYINPUT76), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n275), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n274), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n288));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(KEYINPUT24), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n290), .B1(G169gat), .B2(G176gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(G169gat), .B2(G176gat), .ZN(new_n293));
  OR2_X1    g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(KEYINPUT24), .A3(new_n289), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n291), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT23), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(KEYINPUT64), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n288), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT65), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n293), .A4(new_n295), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n297), .B(KEYINPUT66), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(new_n292), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n305));
  OR3_X1    g104(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT65), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n307), .B(new_n288), .C1(new_n296), .C2(new_n299), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n305), .B1(new_n302), .B2(new_n304), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n301), .A2(new_n306), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT27), .B(G183gat), .ZN(new_n311));
  INV_X1    g110(.A(G190gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(KEYINPUT28), .A3(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT68), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n311), .A2(new_n312), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(KEYINPUT28), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n303), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT26), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n317), .A2(new_n318), .B1(G169gat), .B2(G176gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(new_n318), .B2(new_n297), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n316), .A2(new_n289), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n310), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT29), .B1(new_n310), .B2(new_n321), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(new_n323), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n287), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n324), .B(new_n286), .C1(new_n323), .C2(new_n326), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G8gat), .B(G36gat), .ZN(new_n332));
  INV_X1    g131(.A(G64gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G92gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n339), .B1(new_n330), .B2(new_n336), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n331), .A2(new_n339), .A3(new_n337), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n257), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT82), .ZN(new_n346));
  INV_X1    g145(.A(G228gat), .ZN(new_n347));
  INV_X1    g146(.A(G233gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT29), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n268), .A2(new_n274), .A3(new_n258), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT76), .B1(new_n281), .B2(new_n282), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n281), .B2(new_n282), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n268), .A2(KEYINPUT79), .A3(new_n274), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n350), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g159(.A(KEYINPUT80), .B(new_n350), .C1(new_n353), .C2(new_n357), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n223), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n225), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT29), .B1(new_n222), .B2(new_n223), .ZN(new_n364));
  OR2_X1    g163(.A1(new_n364), .A2(new_n286), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n349), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n223), .B1(new_n287), .B2(KEYINPUT29), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n225), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(KEYINPUT81), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n364), .A2(new_n286), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n368), .A2(new_n349), .A3(new_n369), .A4(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n346), .B(G22gat), .C1(new_n366), .C2(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(G78gat), .B(G106gat), .Z(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT31), .ZN(new_n377));
  INV_X1    g176(.A(G50gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(G22gat), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n370), .B1(new_n362), .B2(new_n225), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n381), .B(new_n373), .C1(new_n382), .C2(new_n349), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT82), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n355), .A2(new_n356), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT29), .B1(new_n385), .B2(new_n284), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT3), .B1(new_n386), .B2(KEYINPUT80), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n222), .B1(new_n387), .B2(new_n360), .ZN(new_n388));
  OAI22_X1  g187(.A1(new_n388), .A2(new_n370), .B1(new_n347), .B2(new_n348), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n381), .B1(new_n389), .B2(new_n373), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n375), .B(new_n380), .C1(new_n384), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT83), .ZN(new_n392));
  OAI21_X1  g191(.A(G22gat), .B1(new_n366), .B2(new_n374), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(KEYINPUT82), .A3(new_n383), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n394), .A2(new_n395), .A3(new_n375), .A4(new_n380), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n393), .A2(new_n383), .A3(new_n379), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT84), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n398), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n402), .B1(new_n392), .B2(new_n396), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT84), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n345), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n322), .A2(new_n214), .ZN(new_n406));
  AND2_X1   g205(.A1(G227gat), .A2(G233gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n310), .A2(new_n321), .A3(new_n215), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT32), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT71), .B(G71gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(G99gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G15gat), .B(G43gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  NAND3_X1  g215(.A1(new_n410), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n416), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n409), .B(KEYINPUT32), .C1(new_n411), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n406), .A2(new_n408), .ZN(new_n421));
  OAI211_X1 g220(.A(KEYINPUT72), .B(KEYINPUT34), .C1(new_n421), .C2(new_n407), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT34), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n407), .B1(new_n406), .B2(new_n408), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT72), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT73), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n417), .A2(new_n422), .A3(new_n426), .A4(new_n419), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  OR3_X1    g230(.A1(new_n420), .A2(new_n427), .A3(new_n429), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n433), .A2(KEYINPUT36), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(KEYINPUT36), .A3(new_n430), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n202), .B1(new_n405), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n343), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n233), .B1(new_n241), .B2(new_n227), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n234), .B1(new_n237), .B2(new_n238), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT39), .ZN(new_n441));
  OR3_X1    g240(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n254), .A2(KEYINPUT86), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT86), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(new_n252), .B2(new_n253), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n446), .B1(new_n439), .B2(new_n441), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n442), .A2(KEYINPUT40), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n442), .A2(new_n447), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT40), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n232), .A2(new_n234), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n443), .B(new_n445), .C1(new_n454), .C2(KEYINPUT39), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n449), .B(new_n451), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n446), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n243), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n438), .A2(new_n448), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT37), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n328), .A2(new_n462), .A3(new_n329), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n336), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT88), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n466), .B(new_n287), .C1(new_n325), .C2(new_n327), .ZN(new_n467));
  OAI211_X1 g266(.A(KEYINPUT37), .B(new_n467), .C1(new_n330), .C2(new_n466), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT38), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n465), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT89), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n338), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n465), .A2(new_n468), .A3(new_n471), .A4(new_n469), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n331), .A2(new_n462), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT38), .B1(new_n474), .B2(new_n464), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n458), .A2(new_n255), .B1(new_n256), .B2(KEYINPUT6), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n461), .B(new_n399), .C1(new_n472), .C2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT84), .B1(new_n397), .B2(new_n398), .ZN(new_n479));
  AOI211_X1 g278(.A(new_n400), .B(new_n402), .C1(new_n392), .C2(new_n396), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n344), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n434), .A2(new_n435), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(KEYINPUT85), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n437), .A2(new_n478), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n428), .A2(new_n430), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n403), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n345), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT35), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n433), .A2(new_n488), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n489), .A2(new_n403), .A3(new_n438), .ZN(new_n490));
  INV_X1    g289(.A(new_n476), .ZN(new_n491));
  AOI22_X1  g290(.A1(KEYINPUT35), .A2(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n484), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n495));
  INV_X1    g294(.A(G155gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(G127gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(G15gat), .A2(G22gat), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(G15gat), .A2(G22gat), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT92), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G1gat), .ZN(new_n503));
  INV_X1    g302(.A(G15gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n381), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT92), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(new_n499), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n502), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n502), .A2(new_n507), .B1(KEYINPUT16), .B2(new_n503), .ZN(new_n510));
  OAI21_X1  g309(.A(G8gat), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n502), .A2(new_n507), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n503), .A2(KEYINPUT16), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G8gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(new_n515), .A3(new_n508), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(G71gat), .B(G78gat), .Z(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT9), .ZN(new_n520));
  INV_X1    g319(.A(G71gat), .ZN(new_n521));
  INV_X1    g320(.A(G78gat), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(G57gat), .B(G64gat), .Z(new_n524));
  NAND3_X1  g323(.A1(new_n519), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n523), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n518), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n517), .B1(KEYINPUT21), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G231gat), .A2(G233gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(G183gat), .B(G211gat), .Z(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n532), .A2(new_n533), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n498), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n536), .ZN(new_n538));
  INV_X1    g337(.A(new_n498), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n529), .A2(KEYINPUT21), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT96), .B(KEYINPUT97), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n537), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n543), .B1(new_n537), .B2(new_n540), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G162gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT7), .B1(new_n250), .B2(new_n335), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT7), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(G85gat), .A3(G92gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G99gat), .A2(G106gat), .ZN(new_n554));
  AOI22_X1  g353(.A1(KEYINPUT8), .A2(new_n554), .B1(new_n250), .B2(new_n335), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G99gat), .B(G106gat), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT98), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n553), .A2(new_n557), .A3(new_n555), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n553), .A2(KEYINPUT98), .A3(new_n557), .A4(new_n555), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT15), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n378), .A2(G43gat), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n565), .B1(new_n566), .B2(KEYINPUT91), .ZN(new_n567));
  NAND2_X1  g366(.A1(G29gat), .A2(G36gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT14), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(G29gat), .B2(G36gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(G29gat), .A2(G36gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT14), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n567), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n571), .B1(KEYINPUT14), .B2(new_n568), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n571), .A2(KEYINPUT14), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n565), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G43gat), .B(G50gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n573), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n577), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n567), .A2(new_n579), .A3(new_n570), .A4(new_n572), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(KEYINPUT17), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n584), .B1(new_n578), .B2(new_n580), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n549), .B(new_n582), .C1(new_n586), .C2(new_n564), .ZN(new_n587));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT99), .B(G134gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n587), .A2(new_n590), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n548), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  INV_X1    g394(.A(new_n548), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n595), .A2(new_n591), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n546), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G230gat), .A2(G233gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n562), .A2(new_n528), .A3(new_n563), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n559), .A2(new_n525), .A3(new_n527), .A4(new_n561), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT100), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n564), .A2(KEYINPUT10), .A3(new_n529), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n605), .B1(new_n604), .B2(new_n606), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n600), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n601), .A2(new_n603), .ZN(new_n610));
  INV_X1    g409(.A(new_n600), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G120gat), .B(G148gat), .ZN(new_n613));
  INV_X1    g412(.A(G176gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(G204gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n609), .A2(new_n612), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n612), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n611), .B1(new_n604), .B2(new_n606), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n599), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n494), .A2(new_n624), .ZN(new_n625));
  NOR3_X1   g424(.A1(new_n509), .A2(new_n510), .A3(G8gat), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n515), .B1(new_n514), .B2(new_n508), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n583), .B2(new_n585), .ZN(new_n629));
  NAND2_X1  g428(.A1(G229gat), .A2(G233gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n517), .A2(new_n581), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT93), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(KEYINPUT18), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n581), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n628), .A2(KEYINPUT94), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT94), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n517), .B2(new_n581), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n639), .A3(new_n631), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n630), .B(KEYINPUT13), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n634), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n629), .A2(new_n630), .A3(new_n631), .A4(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n635), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n646));
  XNOR2_X1  g445(.A(G113gat), .B(G141gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(G169gat), .B(G197gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT12), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n635), .A2(new_n642), .A3(new_n651), .A4(new_n644), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n653), .A2(KEYINPUT95), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT95), .B1(new_n653), .B2(new_n654), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n625), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n257), .B(KEYINPUT101), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(new_n503), .ZN(G1324gat));
  NOR2_X1   g460(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n662));
  AND2_X1   g461(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n663));
  NOR4_X1   g462(.A1(new_n658), .A2(new_n343), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n625), .A2(new_n657), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n515), .B1(new_n665), .B2(new_n438), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT42), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(KEYINPUT42), .B2(new_n664), .ZN(G1325gat));
  NAND3_X1  g467(.A1(new_n665), .A2(new_n504), .A3(new_n433), .ZN(new_n669));
  OAI21_X1  g468(.A(G15gat), .B1(new_n658), .B2(new_n482), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT102), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n669), .A2(new_n673), .A3(new_n670), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(G1326gat));
  NAND2_X1  g474(.A1(new_n401), .A2(new_n404), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n658), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT43), .B(G22gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  INV_X1    g479(.A(new_n598), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n546), .A2(new_n623), .ZN(new_n682));
  AND4_X1   g481(.A1(new_n657), .A2(new_n494), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(G29gat), .ZN(new_n684));
  INV_X1    g483(.A(new_n659), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT45), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n653), .A2(new_n654), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n598), .A2(KEYINPUT105), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n594), .A2(new_n597), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(KEYINPUT44), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n481), .A2(new_n478), .A3(new_n482), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n481), .A2(KEYINPUT103), .A3(new_n478), .A4(new_n482), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n492), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(KEYINPUT104), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701));
  AOI211_X1 g500(.A(new_n701), .B(new_n492), .C1(new_n697), .C2(new_n698), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n694), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n494), .A2(new_n681), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT44), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n689), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n706), .A2(new_n685), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n687), .B1(new_n684), .B2(new_n707), .ZN(G1328gat));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n709));
  INV_X1    g508(.A(G36gat), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(new_n706), .B2(new_n438), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n683), .A2(new_n712), .A3(new_n710), .A4(new_n438), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n598), .B1(new_n484), .B2(new_n493), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n714), .A2(new_n657), .A3(new_n438), .A4(new_n682), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT46), .B1(new_n715), .B2(G36gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n709), .B1(new_n711), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n689), .ZN(new_n719));
  INV_X1    g518(.A(new_n694), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n697), .A2(new_n698), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n493), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n701), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n699), .A2(KEYINPUT104), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n714), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n438), .B(new_n719), .C1(new_n725), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G36gat), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n713), .A2(new_n716), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(new_n730), .A3(KEYINPUT106), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n718), .A2(new_n731), .ZN(G1329gat));
  INV_X1    g531(.A(KEYINPUT47), .ZN(new_n733));
  INV_X1    g532(.A(G43gat), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n706), .B2(new_n436), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n683), .A2(new_n734), .A3(new_n433), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n733), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  AOI211_X1 g537(.A(new_n482), .B(new_n689), .C1(new_n703), .C2(new_n705), .ZN(new_n739));
  OAI211_X1 g538(.A(KEYINPUT47), .B(new_n736), .C1(new_n739), .C2(new_n734), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(G1330gat));
  NAND3_X1  g540(.A1(new_n683), .A2(new_n378), .A3(new_n676), .ZN(new_n742));
  AOI211_X1 g541(.A(new_n399), .B(new_n689), .C1(new_n703), .C2(new_n705), .ZN(new_n743));
  OAI211_X1 g542(.A(KEYINPUT48), .B(new_n742), .C1(new_n743), .C2(new_n378), .ZN(new_n744));
  INV_X1    g543(.A(new_n742), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n676), .B(new_n719), .C1(new_n725), .C2(new_n727), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(G50gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n744), .B1(KEYINPUT48), .B2(new_n747), .ZN(G1331gat));
  INV_X1    g547(.A(new_n688), .ZN(new_n749));
  INV_X1    g548(.A(new_n623), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n599), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n749), .B(new_n751), .C1(new_n700), .C2(new_n702), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n659), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT107), .B(G57gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1332gat));
  INV_X1    g554(.A(KEYINPUT49), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n333), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n343), .B(KEYINPUT108), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n752), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n756), .A2(new_n333), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n758), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NOR4_X1   g563(.A1(new_n752), .A2(KEYINPUT109), .A3(new_n762), .A4(new_n760), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n757), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n688), .B1(new_n723), .B2(new_n724), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n767), .A2(new_n751), .A3(new_n763), .A4(new_n759), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT109), .ZN(new_n769));
  INV_X1    g568(.A(new_n752), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n770), .A2(new_n758), .A3(new_n763), .A4(new_n759), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n769), .A2(new_n771), .A3(new_n756), .A4(new_n333), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n766), .A2(new_n772), .ZN(G1333gat));
  NAND4_X1  g572(.A1(new_n767), .A2(new_n521), .A3(new_n433), .A4(new_n751), .ZN(new_n774));
  OAI21_X1  g573(.A(G71gat), .B1(new_n752), .B2(new_n482), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1334gat));
  NOR2_X1   g577(.A1(new_n752), .A2(new_n677), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(new_n522), .ZN(G1335gat));
  NOR2_X1   g579(.A1(new_n546), .A2(new_n688), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n681), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n722), .A2(KEYINPUT51), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n699), .B2(new_n782), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n750), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n787), .A2(new_n250), .A3(new_n685), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n781), .A2(new_n623), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n789), .B1(new_n703), .B2(new_n705), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n790), .A2(new_n685), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n788), .B1(new_n791), .B2(new_n250), .ZN(G1336gat));
  AOI21_X1  g591(.A(new_n335), .B1(new_n790), .B2(new_n438), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n760), .A2(G92gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n623), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n722), .A2(new_n796), .A3(new_n783), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT110), .B1(new_n699), .B2(new_n782), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(new_n785), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n797), .A2(new_n798), .A3(new_n800), .A4(new_n785), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n795), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT52), .B1(new_n793), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n787), .A2(new_n794), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807));
  AOI211_X1 g606(.A(new_n760), .B(new_n789), .C1(new_n703), .C2(new_n705), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n806), .B(new_n807), .C1(new_n808), .C2(new_n335), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n805), .A2(new_n809), .ZN(G1337gat));
  INV_X1    g609(.A(G99gat), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n787), .A2(new_n811), .A3(new_n433), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n790), .A2(new_n436), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n813), .B2(new_n811), .ZN(G1338gat));
  INV_X1    g613(.A(G106gat), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n790), .B2(new_n676), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n399), .A2(G106gat), .A3(new_n750), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n802), .B2(new_n803), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT53), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n784), .A2(new_n786), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n817), .ZN(new_n823));
  AOI211_X1 g622(.A(new_n399), .B(new_n789), .C1(new_n703), .C2(new_n705), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n821), .B(new_n823), .C1(new_n824), .C2(new_n815), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n820), .A2(new_n825), .ZN(G1339gat));
  NAND3_X1  g625(.A1(new_n604), .A2(new_n611), .A3(new_n606), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n609), .A2(KEYINPUT54), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n618), .B1(new_n621), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n828), .A2(KEYINPUT55), .A3(new_n830), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n833), .A2(new_n688), .A3(new_n619), .A4(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n640), .A2(new_n641), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n630), .B1(new_n629), .B2(new_n631), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n650), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n654), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n623), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT112), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT112), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n835), .A2(new_n843), .A3(new_n840), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n842), .A2(new_n693), .A3(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n833), .A2(new_n619), .A3(new_n839), .A4(new_n834), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n693), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n546), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n599), .A2(new_n688), .A3(new_n623), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n851), .A2(new_n433), .A3(new_n677), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n659), .A2(new_n759), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n657), .ZN(new_n855));
  OAI21_X1  g654(.A(G113gat), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n851), .A2(new_n685), .A3(new_n486), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n759), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n206), .A3(new_n688), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n859), .ZN(G1340gat));
  OAI21_X1  g659(.A(G120gat), .B1(new_n854), .B2(new_n750), .ZN(new_n861));
  INV_X1    g660(.A(new_n211), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n858), .A2(new_n862), .A3(new_n623), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(G1341gat));
  AOI21_X1  g663(.A(G127gat), .B1(new_n858), .B2(new_n546), .ZN(new_n865));
  INV_X1    g664(.A(G127gat), .ZN(new_n866));
  INV_X1    g665(.A(new_n546), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n854), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT113), .Z(G1342gat));
  OAI21_X1  g669(.A(G134gat), .B1(new_n854), .B2(new_n598), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT114), .ZN(new_n872));
  NOR4_X1   g671(.A1(new_n857), .A2(G134gat), .A3(new_n598), .A4(new_n438), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT56), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(G1343gat));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n877), .B1(new_n831), .B2(new_n832), .ZN(new_n878));
  AOI211_X1 g677(.A(KEYINPUT115), .B(KEYINPUT55), .C1(new_n828), .C2(new_n830), .ZN(new_n879));
  OAI22_X1  g678(.A1(new_n878), .A2(new_n879), .B1(new_n655), .B2(new_n656), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n834), .A2(new_n619), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n840), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n598), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n546), .B1(new_n883), .B2(new_n847), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT57), .B1(new_n884), .B2(new_n849), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n876), .B1(new_n885), .B2(new_n677), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(new_n850), .B2(new_n399), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n624), .A2(new_n749), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n693), .A2(new_n846), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n890), .B1(new_n882), .B2(new_n598), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n889), .B1(new_n891), .B2(new_n546), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n892), .A2(KEYINPUT116), .A3(KEYINPUT57), .A4(new_n676), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n886), .A2(new_n888), .A3(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n436), .A2(new_n659), .A3(new_n759), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n657), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G141gat), .ZN(new_n898));
  OR3_X1    g697(.A1(new_n850), .A2(KEYINPUT118), .A3(new_n659), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT118), .B1(new_n850), .B2(new_n659), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n436), .A2(new_n399), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n899), .A2(new_n900), .A3(new_n760), .A4(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n902), .A2(G141gat), .A3(new_n855), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(KEYINPUT58), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n894), .A2(new_n688), .A3(new_n895), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT117), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n906), .A2(new_n907), .A3(G141gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n906), .B2(G141gat), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n908), .A2(new_n909), .A3(new_n903), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT58), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT119), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n914), .B(new_n905), .C1(new_n910), .C2(new_n911), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1344gat));
  INV_X1    g715(.A(new_n902), .ZN(new_n917));
  INV_X1    g716(.A(G148gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n918), .A3(new_n623), .ZN(new_n919));
  XNOR2_X1  g718(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n851), .A2(KEYINPUT57), .A3(new_n403), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT121), .Z(new_n922));
  OAI21_X1  g721(.A(new_n883), .B1(new_n598), .B2(new_n846), .ZN(new_n923));
  AOI22_X1  g722(.A1(new_n923), .A2(new_n867), .B1(new_n855), .B2(new_n624), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n887), .B1(new_n924), .B2(new_n677), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n750), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n895), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n920), .B1(new_n927), .B2(G148gat), .ZN(new_n928));
  AOI211_X1 g727(.A(KEYINPUT59), .B(new_n918), .C1(new_n896), .C2(new_n623), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n919), .B1(new_n928), .B2(new_n929), .ZN(G1345gat));
  AOI21_X1  g729(.A(G155gat), .B1(new_n917), .B2(new_n546), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n867), .A2(new_n496), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n896), .B2(new_n932), .ZN(G1346gat));
  INV_X1    g732(.A(new_n693), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n896), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n935), .A2(KEYINPUT122), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(KEYINPUT122), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(G162gat), .A3(new_n937), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n438), .A2(G162gat), .A3(new_n598), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n899), .A2(new_n901), .A3(new_n900), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1347gat));
  NOR2_X1   g740(.A1(new_n685), .A2(new_n343), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n852), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(G169gat), .B1(new_n943), .B2(new_n855), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n850), .A2(new_n685), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n486), .A3(new_n759), .ZN(new_n946));
  OR3_X1    g745(.A1(new_n946), .A2(G169gat), .A3(new_n749), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n944), .A2(new_n947), .ZN(G1348gat));
  OAI21_X1  g747(.A(new_n614), .B1(new_n946), .B2(new_n750), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT123), .Z(new_n950));
  NOR3_X1   g749(.A1(new_n943), .A2(new_n614), .A3(new_n750), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(G1349gat));
  OAI21_X1  g751(.A(G183gat), .B1(new_n943), .B2(new_n867), .ZN(new_n953));
  INV_X1    g752(.A(new_n946), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n954), .A2(new_n546), .A3(new_n311), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g756(.A(G190gat), .B1(new_n943), .B2(new_n598), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT61), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n960), .B(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n954), .A2(new_n312), .A3(new_n934), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1351gat));
  XNOR2_X1  g763(.A(KEYINPUT126), .B(G197gat), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n922), .A2(new_n925), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n942), .A2(new_n482), .ZN(new_n967));
  XOR2_X1   g766(.A(new_n967), .B(KEYINPUT127), .Z(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n965), .B1(new_n969), .B2(new_n855), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n945), .A2(new_n759), .A3(new_n901), .ZN(new_n971));
  XOR2_X1   g770(.A(new_n971), .B(KEYINPUT125), .Z(new_n972));
  INV_X1    g771(.A(new_n965), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n972), .A2(new_n688), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n970), .A2(new_n974), .ZN(G1352gat));
  NAND3_X1  g774(.A1(new_n971), .A2(new_n616), .A3(new_n623), .ZN(new_n976));
  XOR2_X1   g775(.A(new_n976), .B(KEYINPUT62), .Z(new_n977));
  AND2_X1   g776(.A1(new_n926), .A2(new_n968), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n977), .B1(new_n978), .B2(new_n616), .ZN(G1353gat));
  NAND3_X1  g778(.A1(new_n972), .A2(new_n263), .A3(new_n546), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n966), .A2(new_n546), .A3(new_n968), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n981), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n981), .B2(G211gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(G1354gat));
  NOR3_X1   g783(.A1(new_n969), .A2(new_n264), .A3(new_n598), .ZN(new_n985));
  AOI21_X1  g784(.A(G218gat), .B1(new_n972), .B2(new_n934), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n985), .A2(new_n986), .ZN(G1355gat));
endmodule


