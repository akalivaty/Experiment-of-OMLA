//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT31), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G50gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G228gat), .A2(G233gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT83), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G141gat), .B(G148gat), .Z(new_n208));
  INV_X1    g007(.A(G155gat), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(KEYINPUT2), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G141gat), .B(G148gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n212), .B(new_n211), .C1(new_n216), .C2(KEYINPUT2), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT82), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT82), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224));
  AND2_X1   g023(.A1(G211gat), .A2(G218gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(G211gat), .A2(G218gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AND2_X1   g026(.A1(KEYINPUT76), .A2(G218gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(KEYINPUT76), .A2(G218gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT22), .B1(new_n230), .B2(G211gat), .ZN(new_n231));
  AND2_X1   g030(.A1(G197gat), .A2(G204gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(G197gat), .A2(G204gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n227), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT22), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT76), .B(G218gat), .ZN(new_n237));
  INV_X1    g036(.A(G211gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n227), .ZN(new_n240));
  INV_X1    g039(.A(new_n234), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT29), .B1(new_n235), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT84), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n224), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT29), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n231), .A2(new_n227), .A3(new_n234), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n240), .B1(new_n239), .B2(new_n241), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(KEYINPUT84), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n223), .B1(new_n245), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT77), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n252), .B1(new_n247), .B2(new_n248), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n235), .A2(KEYINPUT77), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n215), .A2(new_n217), .A3(new_n224), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(new_n246), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n207), .B1(new_n251), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n205), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT77), .B1(new_n235), .B2(new_n242), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n248), .A2(new_n252), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n224), .B1(new_n263), .B2(KEYINPUT29), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n260), .B1(new_n264), .B2(new_n218), .ZN(new_n265));
  OAI211_X1 g064(.A(G22gat), .B(new_n204), .C1(new_n258), .C2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT3), .B1(new_n249), .B2(KEYINPUT84), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n243), .A2(new_n244), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n222), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n257), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n206), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n254), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT3), .B1(new_n272), .B2(new_n246), .ZN(new_n273));
  INV_X1    g072(.A(new_n218), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n257), .B(new_n259), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G22gat), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n204), .A2(KEYINPUT85), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n271), .A2(new_n275), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n266), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(G22gat), .B1(new_n258), .B2(new_n265), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n271), .A2(new_n275), .A3(new_n276), .ZN(new_n281));
  INV_X1    g080(.A(new_n277), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G225gat), .A2(G233gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n215), .A2(new_n217), .A3(new_n224), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n224), .B1(new_n215), .B2(new_n217), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G127gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G134gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(KEYINPUT71), .A3(G134gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT70), .B(G134gat), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n293), .B(new_n294), .C1(new_n295), .C2(new_n290), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT1), .ZN(new_n297));
  INV_X1    g096(.A(G113gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(G120gat), .ZN(new_n299));
  INV_X1    g098(.A(G120gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(G113gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n297), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(new_n298), .B2(G120gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n300), .A2(KEYINPUT72), .A3(G113gat), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n305), .B(new_n306), .C1(G113gat), .C2(new_n300), .ZN(new_n307));
  INV_X1    g106(.A(G134gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G127gat), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n291), .A2(new_n309), .A3(new_n297), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n303), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n286), .B1(new_n289), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n296), .A2(new_n302), .B1(new_n310), .B2(new_n307), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n315), .B1(new_n222), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n274), .A2(new_n316), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(KEYINPUT4), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n313), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT5), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n312), .A2(new_n218), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n318), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n321), .B1(new_n323), .B2(new_n286), .ZN(new_n324));
  INV_X1    g123(.A(new_n221), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT82), .B1(new_n215), .B2(new_n217), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n316), .B(new_n315), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n318), .A2(KEYINPUT4), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n327), .A2(new_n328), .B1(new_n312), .B2(new_n289), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n286), .A2(KEYINPUT5), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n320), .A2(new_n324), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT0), .B(G57gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(G85gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(G1gat), .B(G29gat), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n333), .B(new_n334), .Z(new_n335));
  OAI21_X1  g134(.A(KEYINPUT86), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n316), .B1(new_n325), .B2(new_n326), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n312), .A2(new_n218), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT4), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n337), .A2(new_n314), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n218), .A2(KEYINPUT3), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(new_n312), .A3(new_n255), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n285), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n324), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n328), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(new_n342), .A3(new_n330), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT86), .ZN(new_n348));
  INV_X1    g147(.A(new_n335), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n336), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n344), .A2(new_n335), .A3(new_n346), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT6), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n347), .A2(KEYINPUT6), .A3(new_n349), .ZN(new_n357));
  INV_X1    g156(.A(G226gat), .ZN(new_n358));
  INV_X1    g157(.A(G233gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(G183gat), .A2(G190gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT65), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT65), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n368), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G169gat), .A2(G176gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT23), .ZN(new_n373));
  INV_X1    g172(.A(G169gat), .ZN(new_n374));
  INV_X1    g173(.A(G176gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n372), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n370), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n366), .A2(KEYINPUT66), .ZN(new_n381));
  NAND2_X1  g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT24), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  OR2_X1    g184(.A1(new_n364), .A2(KEYINPUT67), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n364), .A2(KEYINPUT67), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n382), .A2(KEYINPUT66), .A3(new_n383), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  AOI211_X1 g188(.A(new_n380), .B(new_n372), .C1(new_n376), .C2(new_n377), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n379), .A2(new_n380), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT68), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT26), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(new_n374), .A3(new_n375), .ZN(new_n396));
  OAI211_X1 g195(.A(KEYINPUT68), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n394), .A2(new_n371), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT27), .B(G183gat), .ZN(new_n399));
  INV_X1    g198(.A(G190gat), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT28), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AND2_X1   g200(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n403));
  OAI211_X1 g202(.A(KEYINPUT28), .B(new_n400), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n382), .B(new_n398), .C1(new_n401), .C2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n362), .B1(new_n391), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n378), .A2(KEYINPUT25), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n363), .B1(KEYINPUT66), .B2(new_n366), .ZN(new_n410));
  INV_X1    g209(.A(new_n388), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n386), .A2(new_n387), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT25), .B1(new_n370), .B2(new_n378), .ZN(new_n415));
  OAI211_X1 g214(.A(KEYINPUT78), .B(new_n406), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n361), .B1(new_n408), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n360), .A2(KEYINPUT29), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n406), .A2(KEYINPUT69), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n398), .A2(new_n382), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT69), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT28), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n404), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n421), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n379), .A2(new_n380), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n389), .A2(new_n390), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n419), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n263), .B1(new_n417), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n408), .A2(new_n418), .A3(new_n416), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(new_n360), .A3(new_n431), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n272), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT37), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n416), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT78), .B1(new_n431), .B2(new_n406), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n360), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n406), .A2(KEYINPUT69), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n422), .B1(new_n421), .B2(new_n426), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n431), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n418), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n442), .A2(new_n272), .A3(new_n446), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n434), .A2(new_n435), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n447), .B(KEYINPUT37), .C1(new_n448), .C2(new_n272), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT38), .ZN(new_n450));
  XNOR2_X1  g249(.A(G8gat), .B(G36gat), .ZN(new_n451));
  INV_X1    g250(.A(G64gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(G92gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT79), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n439), .A2(new_n449), .A3(new_n450), .A4(new_n455), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n356), .A2(new_n357), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n454), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(new_n433), .B2(new_n436), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n272), .B1(new_n442), .B2(new_n446), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n434), .A2(new_n272), .A3(new_n435), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT37), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(new_n458), .A3(new_n439), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n459), .B1(new_n464), .B2(KEYINPUT38), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n284), .B1(new_n457), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n454), .B1(new_n460), .B2(new_n461), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT30), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n467), .A2(new_n468), .B1(new_n462), .B2(new_n455), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n459), .A2(KEYINPUT80), .A3(KEYINPUT30), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT80), .B1(new_n459), .B2(KEYINPUT30), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OR3_X1    g271(.A1(new_n329), .A2(KEYINPUT39), .A3(new_n285), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n322), .A2(new_n285), .A3(new_n318), .ZN(new_n474));
  OAI211_X1 g273(.A(KEYINPUT39), .B(new_n474), .C1(new_n329), .C2(new_n285), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n473), .A2(new_n335), .A3(new_n475), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n476), .A2(KEYINPUT40), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n476), .A2(KEYINPUT40), .B1(new_n336), .B2(new_n350), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n472), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT87), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n472), .A2(new_n477), .A3(new_n478), .A4(KEYINPUT87), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n484));
  AOI211_X1 g283(.A(new_n312), .B(new_n391), .C1(new_n420), .C2(new_n427), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n316), .B1(new_n428), .B2(new_n431), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G227gat), .A2(G233gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(KEYINPUT64), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n484), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n445), .A2(new_n312), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n428), .A2(new_n316), .A3(new_n431), .ZN(new_n493));
  NAND2_X1  g292(.A1(KEYINPUT74), .A2(KEYINPUT34), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n492), .A2(new_n490), .A3(new_n493), .A4(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(KEYINPUT73), .B(G71gat), .ZN(new_n499));
  INV_X1    g298(.A(G99gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G15gat), .B(G43gat), .ZN(new_n502));
  XOR2_X1   g301(.A(new_n501), .B(new_n502), .Z(new_n503));
  AOI21_X1  g302(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(KEYINPUT33), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT32), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n489), .B1(new_n485), .B2(new_n486), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT33), .ZN(new_n510));
  INV_X1    g309(.A(new_n503), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n509), .B(KEYINPUT32), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n498), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT75), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n509), .A2(KEYINPUT32), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n509), .A2(new_n510), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n503), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n492), .A2(new_n493), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(new_n489), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n496), .B1(new_n520), .B2(new_n484), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n521), .A3(new_n512), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n514), .A2(new_n515), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT36), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n521), .B1(new_n518), .B2(new_n512), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT75), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n518), .A2(new_n521), .A3(new_n512), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n528), .A2(new_n525), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT36), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n331), .A2(new_n335), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n357), .B1(new_n354), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n532), .B(new_n469), .C1(new_n470), .C2(new_n471), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n527), .A2(new_n530), .B1(new_n284), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n483), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n284), .B1(new_n523), .B2(new_n526), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT35), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n356), .A2(new_n357), .ZN(new_n538));
  INV_X1    g337(.A(new_n455), .ZN(new_n539));
  OAI22_X1  g338(.A1(new_n459), .A2(KEYINPUT30), .B1(new_n437), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT80), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(new_n467), .B2(new_n468), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n459), .A2(KEYINPUT80), .A3(KEYINPUT30), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT88), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n538), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n357), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n547), .B1(new_n351), .B2(new_n355), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT88), .B1(new_n472), .B2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n536), .A2(new_n537), .A3(new_n546), .A4(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n514), .A2(new_n522), .A3(new_n279), .A4(new_n283), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT35), .B1(new_n551), .B2(new_n533), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT89), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT89), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n554), .B(KEYINPUT35), .C1(new_n551), .C2(new_n533), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n452), .A2(G57gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n452), .A2(G57gat), .ZN(new_n559));
  AND2_X1   g358(.A1(G71gat), .A2(G78gat), .ZN(new_n560));
  OAI22_X1  g359(.A1(new_n558), .A2(new_n559), .B1(KEYINPUT9), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G71gat), .B(G78gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT96), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(KEYINPUT96), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT21), .ZN(new_n569));
  XNOR2_X1  g368(.A(G15gat), .B(G22gat), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT16), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n570), .B1(new_n571), .B2(G1gat), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(G1gat), .B2(new_n570), .ZN(new_n573));
  INV_X1    g372(.A(G8gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(G183gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n576), .A2(G183gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n578), .B2(new_n579), .ZN(new_n584));
  XNOR2_X1  g383(.A(G127gat), .B(G155gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n568), .A2(KEYINPUT21), .ZN(new_n588));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(G211gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n590), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n579), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n580), .B1(new_n594), .B2(new_n577), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n585), .B1(new_n595), .B2(new_n582), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n587), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n593), .B1(new_n587), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G43gat), .B(G50gat), .Z(new_n600));
  INV_X1    g399(.A(KEYINPUT15), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT14), .ZN(new_n604));
  INV_X1    g403(.A(G29gat), .ZN(new_n605));
  INV_X1    g404(.A(G36gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n607), .A2(new_n608), .B1(G29gat), .B2(G36gat), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n602), .A2(new_n603), .A3(new_n609), .ZN(new_n610));
  OR3_X1    g409(.A1(new_n609), .A2(new_n601), .A3(new_n600), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT17), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT99), .B(G85gat), .ZN(new_n615));
  INV_X1    g414(.A(G92gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G85gat), .A2(G92gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT7), .ZN(new_n619));
  INV_X1    g418(.A(G106gat), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT8), .B1(new_n500), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G99gat), .B(G106gat), .Z(new_n623));
  OR2_X1    g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n610), .A2(KEYINPUT17), .A3(new_n611), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n614), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n624), .A2(new_n625), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n612), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT41), .ZN(new_n631));
  NAND2_X1  g430(.A1(G232gat), .A2(G233gat), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n628), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G134gat), .B(G162gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G190gat), .B(G218gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT100), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n632), .A2(new_n631), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n635), .B(new_n639), .Z(new_n640));
  NOR2_X1   g439(.A1(new_n599), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT91), .ZN(new_n643));
  XOR2_X1   g442(.A(G113gat), .B(G141gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G169gat), .B(G197gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT12), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n614), .A2(new_n575), .A3(new_n627), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT92), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n573), .B(G8gat), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n651), .B1(new_n652), .B2(new_n612), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n614), .A2(new_n575), .A3(new_n651), .A4(new_n627), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G229gat), .A2(G233gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n575), .B(new_n612), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n657), .B(KEYINPUT13), .ZN(new_n661));
  OAI22_X1  g460(.A1(new_n658), .A2(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT93), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n656), .A2(KEYINPUT93), .A3(new_n657), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(new_n659), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n649), .B1(new_n663), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT95), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT93), .B1(new_n656), .B2(new_n657), .ZN(new_n670));
  INV_X1    g469(.A(new_n657), .ZN(new_n671));
  AOI211_X1 g470(.A(new_n664), .B(new_n671), .C1(new_n654), .C2(new_n655), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n670), .A2(new_n672), .A3(KEYINPUT18), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n649), .B1(new_n673), .B2(KEYINPUT94), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT94), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n663), .B1(new_n667), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n669), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n662), .B1(new_n673), .B2(KEYINPUT94), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n648), .B1(new_n667), .B2(new_n675), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(new_n679), .A3(KEYINPUT95), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n668), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(G230gat), .A2(G233gat), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n568), .A2(new_n626), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n626), .A2(new_n563), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT10), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n568), .A2(KEYINPUT101), .A3(KEYINPUT10), .A4(new_n629), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n563), .B(new_n565), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n624), .A2(KEYINPUT10), .A3(new_n625), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n682), .B1(new_n686), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n682), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n683), .A2(new_n694), .A3(new_n685), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(G176gat), .B(G204gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT102), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(G120gat), .ZN(new_n699));
  INV_X1    g498(.A(G148gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n696), .A2(new_n701), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n681), .A2(new_n705), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n557), .A2(new_n641), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n532), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g509(.A1(new_n707), .A2(new_n472), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(KEYINPUT42), .Z(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n574), .B2(new_n711), .ZN(G1325gat));
  NAND2_X1  g514(.A1(new_n523), .A2(new_n526), .ZN(new_n716));
  AOI21_X1  g515(.A(G15gat), .B1(new_n707), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n527), .A2(new_n530), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G15gat), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT103), .Z(new_n721));
  AOI21_X1  g520(.A(new_n717), .B1(new_n707), .B2(new_n721), .ZN(G1326gat));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n284), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT43), .B(G22gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1327gat));
  AND3_X1   g524(.A1(new_n283), .A2(new_n266), .A3(new_n278), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n529), .A2(new_n544), .A3(new_n726), .A4(new_n532), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n554), .B1(new_n727), .B2(KEYINPUT35), .ZN(new_n728));
  INV_X1    g527(.A(new_n555), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT104), .B1(new_n730), .B2(new_n550), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n550), .A2(new_n553), .A3(KEYINPUT104), .A4(new_n555), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n535), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(new_n640), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n557), .A2(new_n640), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT44), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n706), .A2(new_n599), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(G29gat), .B1(new_n742), .B2(new_n532), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n737), .A2(new_n740), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n605), .A3(new_n708), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT45), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(G1328gat));
  OAI21_X1  g546(.A(G36gat), .B1(new_n742), .B2(new_n544), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n744), .A2(new_n606), .A3(new_n472), .ZN(new_n749));
  AND2_X1   g548(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n748), .B(new_n752), .C1(new_n750), .C2(new_n749), .ZN(G1329gat));
  INV_X1    g552(.A(new_n742), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(G43gat), .A3(new_n719), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n744), .A2(new_n716), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(G43gat), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g557(.A1(new_n754), .A2(G50gat), .A3(new_n284), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n737), .A2(new_n726), .A3(new_n740), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(G50gat), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g561(.A1(new_n641), .A2(new_n734), .A3(new_n705), .A4(new_n681), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n532), .B(KEYINPUT107), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G57gat), .ZN(G1332gat));
  INV_X1    g566(.A(KEYINPUT49), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n763), .B(new_n472), .C1(new_n768), .C2(new_n452), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n452), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1333gat));
  NAND3_X1  g570(.A1(new_n763), .A2(G71gat), .A3(new_n719), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n763), .A2(new_n716), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(KEYINPUT108), .Z(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n774), .B2(G71gat), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g575(.A1(new_n763), .A2(new_n284), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g577(.A1(new_n599), .A2(new_n681), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(KEYINPUT109), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n599), .B2(new_n681), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n705), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n739), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n708), .ZN(new_n787));
  XOR2_X1   g586(.A(new_n787), .B(KEYINPUT110), .Z(new_n788));
  INV_X1    g587(.A(new_n640), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT104), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n556), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n732), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n789), .B1(new_n792), .B2(new_n535), .ZN(new_n793));
  INV_X1    g592(.A(new_n783), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n793), .A2(KEYINPUT51), .A3(new_n794), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n705), .A2(new_n708), .A3(new_n615), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT111), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n788), .A2(new_n615), .B1(new_n800), .B2(new_n802), .ZN(G1336gat));
  INV_X1    g602(.A(new_n786), .ZN(new_n804));
  OAI21_X1  g603(.A(G92gat), .B1(new_n804), .B2(new_n544), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n799), .A2(new_n616), .A3(new_n705), .A4(new_n472), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g607(.A(G99gat), .B1(new_n804), .B2(new_n718), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n716), .A2(new_n500), .A3(new_n705), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT112), .Z(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n800), .B2(new_n811), .ZN(G1338gat));
  NAND4_X1  g611(.A1(new_n799), .A2(new_n620), .A3(new_n705), .A4(new_n284), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n483), .A2(new_n534), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n791), .B2(new_n732), .ZN(new_n815));
  INV_X1    g614(.A(new_n735), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n815), .A2(new_n789), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n738), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n284), .B(new_n785), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(G106gat), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n813), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT53), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT51), .B1(new_n793), .B2(new_n794), .ZN(new_n823));
  NOR4_X1   g622(.A1(new_n815), .A2(new_n783), .A3(new_n796), .A4(new_n789), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n705), .B(new_n284), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT53), .B1(new_n826), .B2(new_n620), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n819), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n739), .A2(KEYINPUT113), .A3(new_n284), .A4(new_n785), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(G106gat), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT114), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n833));
  AND4_X1   g632(.A1(KEYINPUT114), .A2(new_n831), .A3(new_n833), .A4(new_n813), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n822), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g636(.A(KEYINPUT115), .B(new_n822), .C1(new_n832), .C2(new_n834), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1339gat));
  NAND3_X1  g638(.A1(new_n641), .A2(new_n784), .A3(new_n681), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n677), .A2(new_n680), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n656), .A2(new_n657), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(new_n660), .B2(new_n661), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n647), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n640), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT10), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n689), .A2(new_n629), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(new_n684), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n851), .A2(new_n694), .A3(new_n687), .A4(new_n691), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n693), .A2(new_n852), .A3(KEYINPUT54), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n854), .B(new_n682), .C1(new_n686), .C2(new_n692), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n701), .A3(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT55), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n853), .A2(KEYINPUT55), .A3(new_n701), .A4(new_n855), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n703), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT116), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n702), .B1(new_n856), .B2(new_n857), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n863), .A3(new_n859), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n842), .B1(new_n848), .B2(new_n865), .ZN(new_n866));
  AND4_X1   g665(.A1(new_n863), .A2(new_n858), .A3(new_n703), .A4(new_n859), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n863), .B1(new_n862), .B2(new_n859), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n846), .B1(new_n677), .B2(new_n680), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n869), .A2(KEYINPUT117), .A3(new_n640), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n705), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n873), .B1(new_n865), .B2(new_n681), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n789), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n841), .B1(new_n876), .B2(new_n599), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(new_n472), .A3(new_n764), .ZN(new_n878));
  INV_X1    g677(.A(new_n551), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n681), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n298), .A3(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n877), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n472), .A2(new_n532), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n536), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n882), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n883), .B1(new_n298), .B2(new_n890), .ZN(G1340gat));
  NAND3_X1  g690(.A1(new_n881), .A2(new_n300), .A3(new_n705), .ZN(new_n892));
  OAI21_X1  g691(.A(G120gat), .B1(new_n887), .B2(new_n784), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g693(.A(new_n894), .B(KEYINPUT118), .Z(G1341gat));
  OR3_X1    g694(.A1(new_n880), .A2(KEYINPUT119), .A3(new_n599), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT119), .B1(new_n880), .B2(new_n599), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n290), .A3(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n599), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n888), .A2(G127gat), .A3(new_n899), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n898), .A2(new_n900), .ZN(G1342gat));
  NOR3_X1   g700(.A1(new_n880), .A2(new_n295), .A3(new_n789), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT56), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G134gat), .B1(new_n887), .B2(new_n789), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n902), .A2(new_n903), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(G1343gat));
  INV_X1    g706(.A(new_n856), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(KEYINPUT120), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n857), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n703), .B1(new_n909), .B2(new_n857), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n911), .A2(new_n681), .A3(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n873), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n789), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n899), .B1(new_n915), .B2(new_n872), .ZN(new_n916));
  OAI211_X1 g715(.A(KEYINPUT57), .B(new_n284), .C1(new_n916), .C2(new_n841), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT121), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n908), .A2(KEYINPUT120), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n702), .B1(new_n919), .B2(KEYINPUT55), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n882), .A2(new_n910), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n873), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n922), .A2(new_n789), .B1(new_n866), .B2(new_n871), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n840), .B1(new_n923), .B2(new_n899), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n924), .A2(new_n925), .A3(KEYINPUT57), .A4(new_n284), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT57), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n927), .B1(new_n877), .B2(new_n726), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n918), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n718), .A2(new_n885), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n882), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G141gat), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n719), .A2(new_n726), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n878), .A2(new_n935), .ZN(new_n936));
  OR3_X1    g735(.A1(new_n936), .A2(G141gat), .A3(new_n681), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT58), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT58), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1344gat));
  NAND3_X1  g741(.A1(new_n929), .A2(new_n705), .A3(new_n931), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(new_n944), .A3(G148gat), .ZN(new_n945));
  OAI21_X1  g744(.A(KEYINPUT57), .B1(new_n877), .B2(new_n726), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n848), .A2(new_n860), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n899), .B1(new_n915), .B2(new_n947), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n927), .B(new_n284), .C1(new_n948), .C2(new_n841), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n946), .A2(new_n705), .A3(new_n931), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G148gat), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT59), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n945), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n878), .A2(new_n700), .A3(new_n705), .A4(new_n935), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT122), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n953), .A2(new_n954), .A3(KEYINPUT122), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1345gat));
  NAND3_X1  g758(.A1(new_n932), .A2(G155gat), .A3(new_n899), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n209), .B1(new_n936), .B2(new_n599), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(G1346gat));
  NAND3_X1  g761(.A1(new_n932), .A2(G162gat), .A3(new_n640), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n210), .B1(new_n936), .B2(new_n789), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n963), .A2(new_n964), .ZN(G1347gat));
  NOR2_X1   g764(.A1(new_n765), .A2(new_n544), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n966), .A2(KEYINPUT124), .A3(new_n716), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT124), .B1(new_n966), .B2(new_n716), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n968), .A2(new_n284), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n884), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(G169gat), .B1(new_n970), .B2(new_n681), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n877), .A2(new_n708), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n972), .A2(new_n472), .A3(new_n879), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n974), .A2(new_n374), .A3(new_n882), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT123), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n971), .B1(new_n977), .B2(new_n978), .ZN(G1348gat));
  NOR3_X1   g778(.A1(new_n970), .A2(new_n375), .A3(new_n784), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n974), .A2(new_n705), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n980), .B1(new_n981), .B2(new_n375), .ZN(G1349gat));
  OAI21_X1  g781(.A(G183gat), .B1(new_n970), .B2(new_n599), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n899), .A2(new_n399), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n983), .B1(new_n973), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g785(.A(G190gat), .B1(new_n970), .B2(new_n789), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n988));
  OR2_X1    g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  NAND2_X1  g794(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n996));
  NAND4_X1  g795(.A1(new_n989), .A2(new_n995), .A3(new_n996), .A4(new_n990), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n974), .A2(new_n400), .A3(new_n640), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n994), .A2(new_n997), .A3(new_n998), .ZN(G1351gat));
  NAND3_X1  g798(.A1(new_n972), .A2(new_n472), .A3(new_n935), .ZN(new_n1000));
  INV_X1    g799(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g800(.A(G197gat), .B1(new_n1001), .B2(new_n882), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n946), .A2(new_n949), .ZN(new_n1003));
  INV_X1    g802(.A(G197gat), .ZN(new_n1004));
  AND2_X1   g803(.A1(new_n966), .A2(new_n718), .ZN(new_n1005));
  XNOR2_X1  g804(.A(new_n1005), .B(KEYINPUT127), .ZN(new_n1006));
  NOR4_X1   g805(.A1(new_n1003), .A2(new_n1004), .A3(new_n681), .A4(new_n1006), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n1002), .A2(new_n1007), .ZN(G1352gat));
  NOR3_X1   g807(.A1(new_n1000), .A2(G204gat), .A3(new_n784), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n1010));
  OR2_X1    g809(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g810(.A(new_n1003), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1012), .A2(new_n705), .ZN(new_n1013));
  OAI21_X1  g812(.A(G204gat), .B1(new_n1013), .B2(new_n1006), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1011), .A2(new_n1014), .A3(new_n1015), .ZN(G1353gat));
  NAND3_X1  g815(.A1(new_n1012), .A2(new_n899), .A3(new_n1005), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1017), .A2(G211gat), .ZN(new_n1018));
  XOR2_X1   g817(.A(new_n1018), .B(KEYINPUT63), .Z(new_n1019));
  NAND3_X1  g818(.A1(new_n1001), .A2(new_n238), .A3(new_n899), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1019), .A2(new_n1020), .ZN(G1354gat));
  AOI21_X1  g820(.A(G218gat), .B1(new_n1001), .B2(new_n640), .ZN(new_n1022));
  NOR3_X1   g821(.A1(new_n1006), .A2(new_n789), .A3(new_n237), .ZN(new_n1023));
  AOI21_X1  g822(.A(new_n1022), .B1(new_n1012), .B2(new_n1023), .ZN(G1355gat));
endmodule


