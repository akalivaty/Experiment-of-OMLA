

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U547 ( .A1(n724), .A2(G1341), .ZN(n511) );
  AND2_X1 U548 ( .A1(n685), .A2(n684), .ZN(n687) );
  INV_X1 U549 ( .A(KEYINPUT29), .ZN(n707) );
  NOR2_X1 U550 ( .A1(G1384), .A2(G164), .ZN(n752) );
  NOR2_X1 U551 ( .A1(G651), .A2(G543), .ZN(n642) );
  NOR2_X1 U552 ( .A1(G651), .A2(n628), .ZN(n646) );
  NOR2_X1 U553 ( .A1(n521), .A2(n520), .ZN(G160) );
  INV_X1 U554 ( .A(G2105), .ZN(n517) );
  AND2_X2 U555 ( .A1(n517), .A2(G2104), .ZN(n868) );
  NAND2_X1 U556 ( .A1(G101), .A2(n868), .ZN(n512) );
  XOR2_X1 U557 ( .A(KEYINPUT66), .B(n512), .Z(n513) );
  XNOR2_X1 U558 ( .A(n513), .B(KEYINPUT23), .ZN(n516) );
  NOR2_X1 U559 ( .A1(G2104), .A2(G2105), .ZN(n514) );
  XOR2_X2 U560 ( .A(KEYINPUT17), .B(n514), .Z(n867) );
  NAND2_X1 U561 ( .A1(G137), .A2(n867), .ZN(n515) );
  NAND2_X1 U562 ( .A1(n516), .A2(n515), .ZN(n521) );
  AND2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n871) );
  NAND2_X1 U564 ( .A1(G113), .A2(n871), .ZN(n519) );
  NOR2_X1 U565 ( .A1(G2104), .A2(n517), .ZN(n872) );
  NAND2_X1 U566 ( .A1(G125), .A2(n872), .ZN(n518) );
  NAND2_X1 U567 ( .A1(n519), .A2(n518), .ZN(n520) );
  NAND2_X1 U568 ( .A1(G138), .A2(n867), .ZN(n523) );
  NAND2_X1 U569 ( .A1(G126), .A2(n872), .ZN(n522) );
  NAND2_X1 U570 ( .A1(n523), .A2(n522), .ZN(n527) );
  NAND2_X1 U571 ( .A1(G114), .A2(n871), .ZN(n525) );
  NAND2_X1 U572 ( .A1(G102), .A2(n868), .ZN(n524) );
  NAND2_X1 U573 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U574 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U575 ( .A(KEYINPUT88), .B(n528), .ZN(G164) );
  NAND2_X1 U576 ( .A1(n642), .A2(G89), .ZN(n529) );
  XNOR2_X1 U577 ( .A(n529), .B(KEYINPUT4), .ZN(n531) );
  XOR2_X1 U578 ( .A(G543), .B(KEYINPUT0), .Z(n628) );
  INV_X1 U579 ( .A(G651), .ZN(n533) );
  NOR2_X1 U580 ( .A1(n628), .A2(n533), .ZN(n639) );
  NAND2_X1 U581 ( .A1(G76), .A2(n639), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U583 ( .A(KEYINPUT5), .B(n532), .ZN(n541) );
  NAND2_X1 U584 ( .A1(G51), .A2(n646), .ZN(n537) );
  NOR2_X1 U585 ( .A1(G543), .A2(n533), .ZN(n535) );
  XNOR2_X1 U586 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n534) );
  XNOR2_X1 U587 ( .A(n535), .B(n534), .ZN(n643) );
  NAND2_X1 U588 ( .A1(n643), .A2(G63), .ZN(n536) );
  NAND2_X1 U589 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U590 ( .A(n538), .B(KEYINPUT6), .ZN(n539) );
  XOR2_X1 U591 ( .A(KEYINPUT72), .B(n539), .Z(n540) );
  NAND2_X1 U592 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U593 ( .A(KEYINPUT7), .B(n542), .ZN(G168) );
  XOR2_X1 U594 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U595 ( .A1(G85), .A2(n642), .ZN(n544) );
  NAND2_X1 U596 ( .A1(G60), .A2(n643), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U598 ( .A1(G72), .A2(n639), .ZN(n546) );
  NAND2_X1 U599 ( .A1(G47), .A2(n646), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U601 ( .A1(n548), .A2(n547), .ZN(G290) );
  XOR2_X1 U602 ( .A(G2438), .B(G2454), .Z(n550) );
  XNOR2_X1 U603 ( .A(G2435), .B(G2430), .ZN(n549) );
  XNOR2_X1 U604 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U605 ( .A(n551), .B(G2427), .Z(n553) );
  XNOR2_X1 U606 ( .A(G1348), .B(G1341), .ZN(n552) );
  XNOR2_X1 U607 ( .A(n553), .B(n552), .ZN(n557) );
  XOR2_X1 U608 ( .A(G2443), .B(G2446), .Z(n555) );
  XNOR2_X1 U609 ( .A(KEYINPUT106), .B(G2451), .ZN(n554) );
  XNOR2_X1 U610 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U611 ( .A(n557), .B(n556), .Z(n558) );
  AND2_X1 U612 ( .A1(G14), .A2(n558), .ZN(G401) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U614 ( .A1(G111), .A2(n871), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G99), .A2(n868), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(n563) );
  NAND2_X1 U617 ( .A1(n872), .A2(G123), .ZN(n561) );
  XOR2_X1 U618 ( .A(KEYINPUT18), .B(n561), .Z(n562) );
  NOR2_X1 U619 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U620 ( .A1(n867), .A2(G135), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n565), .A2(n564), .ZN(n910) );
  XNOR2_X1 U622 ( .A(G2096), .B(n910), .ZN(n566) );
  OR2_X1 U623 ( .A1(G2100), .A2(n566), .ZN(G156) );
  INV_X1 U624 ( .A(G132), .ZN(G219) );
  INV_X1 U625 ( .A(G82), .ZN(G220) );
  NAND2_X1 U626 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U627 ( .A(n567), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U628 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n569) );
  INV_X1 U629 ( .A(G223), .ZN(n818) );
  NAND2_X1 U630 ( .A1(G567), .A2(n818), .ZN(n568) );
  XNOR2_X1 U631 ( .A(n569), .B(n568), .ZN(G234) );
  NAND2_X1 U632 ( .A1(G56), .A2(n643), .ZN(n570) );
  XOR2_X1 U633 ( .A(KEYINPUT14), .B(n570), .Z(n576) );
  NAND2_X1 U634 ( .A1(n642), .A2(G81), .ZN(n571) );
  XNOR2_X1 U635 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U636 ( .A1(G68), .A2(n639), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT13), .B(n574), .Z(n575) );
  NOR2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n646), .A2(G43), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n578), .A2(n577), .ZN(n979) );
  INV_X1 U642 ( .A(G860), .ZN(n607) );
  OR2_X1 U643 ( .A1(n979), .A2(n607), .ZN(G153) );
  NAND2_X1 U644 ( .A1(G90), .A2(n642), .ZN(n580) );
  NAND2_X1 U645 ( .A1(G77), .A2(n639), .ZN(n579) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(KEYINPUT9), .B(n581), .ZN(n585) );
  NAND2_X1 U648 ( .A1(G64), .A2(n643), .ZN(n583) );
  NAND2_X1 U649 ( .A1(G52), .A2(n646), .ZN(n582) );
  AND2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(G301) );
  NAND2_X1 U652 ( .A1(G92), .A2(n642), .ZN(n587) );
  NAND2_X1 U653 ( .A1(G66), .A2(n643), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U655 ( .A1(G79), .A2(n639), .ZN(n589) );
  NAND2_X1 U656 ( .A1(G54), .A2(n646), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U658 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U659 ( .A(KEYINPUT15), .B(n592), .Z(n981) );
  NOR2_X1 U660 ( .A1(n981), .A2(G868), .ZN(n593) );
  XNOR2_X1 U661 ( .A(n593), .B(KEYINPUT71), .ZN(n595) );
  NAND2_X1 U662 ( .A1(G868), .A2(G301), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G91), .A2(n642), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G78), .A2(n639), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n643), .A2(G65), .ZN(n598) );
  XOR2_X1 U668 ( .A(KEYINPUT68), .B(n598), .Z(n599) );
  NOR2_X1 U669 ( .A1(n600), .A2(n599), .ZN(n602) );
  NAND2_X1 U670 ( .A1(n646), .A2(G53), .ZN(n601) );
  NAND2_X1 U671 ( .A1(n602), .A2(n601), .ZN(G299) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n603) );
  XOR2_X1 U673 ( .A(KEYINPUT73), .B(n603), .Z(n605) );
  INV_X1 U674 ( .A(G868), .ZN(n652) );
  NOR2_X1 U675 ( .A1(G286), .A2(n652), .ZN(n604) );
  NOR2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U677 ( .A(KEYINPUT74), .B(n606), .ZN(G297) );
  NAND2_X1 U678 ( .A1(n607), .A2(G559), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n608), .A2(n981), .ZN(n609) );
  XNOR2_X1 U680 ( .A(n609), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n979), .ZN(n612) );
  NAND2_X1 U682 ( .A1(n981), .A2(G868), .ZN(n610) );
  NOR2_X1 U683 ( .A1(G559), .A2(n610), .ZN(n611) );
  NOR2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U685 ( .A(KEYINPUT75), .B(n613), .Z(G282) );
  NAND2_X1 U686 ( .A1(G559), .A2(n981), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n979), .B(n614), .ZN(n661) );
  NOR2_X1 U688 ( .A1(n661), .A2(G860), .ZN(n623) );
  NAND2_X1 U689 ( .A1(G80), .A2(n639), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G67), .A2(n643), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U692 ( .A1(G93), .A2(n642), .ZN(n617) );
  XNOR2_X1 U693 ( .A(KEYINPUT77), .B(n617), .ZN(n618) );
  NOR2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n646), .A2(G55), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n655) );
  XOR2_X1 U697 ( .A(n655), .B(KEYINPUT76), .Z(n622) );
  XNOR2_X1 U698 ( .A(n623), .B(n622), .ZN(G145) );
  NAND2_X1 U699 ( .A1(G49), .A2(n646), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U702 ( .A1(n643), .A2(n626), .ZN(n627) );
  XNOR2_X1 U703 ( .A(n627), .B(KEYINPUT78), .ZN(n630) );
  NAND2_X1 U704 ( .A1(G87), .A2(n628), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n630), .A2(n629), .ZN(G288) );
  NAND2_X1 U706 ( .A1(G88), .A2(n642), .ZN(n631) );
  XNOR2_X1 U707 ( .A(n631), .B(KEYINPUT82), .ZN(n638) );
  NAND2_X1 U708 ( .A1(G75), .A2(n639), .ZN(n633) );
  NAND2_X1 U709 ( .A1(G50), .A2(n646), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U711 ( .A1(G62), .A2(n643), .ZN(n634) );
  XNOR2_X1 U712 ( .A(KEYINPUT81), .B(n634), .ZN(n635) );
  NOR2_X1 U713 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(G303) );
  XOR2_X1 U715 ( .A(KEYINPUT79), .B(KEYINPUT2), .Z(n641) );
  NAND2_X1 U716 ( .A1(G73), .A2(n639), .ZN(n640) );
  XNOR2_X1 U717 ( .A(n641), .B(n640), .ZN(n651) );
  NAND2_X1 U718 ( .A1(G86), .A2(n642), .ZN(n645) );
  NAND2_X1 U719 ( .A1(G61), .A2(n643), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n646), .A2(G48), .ZN(n647) );
  XOR2_X1 U722 ( .A(KEYINPUT80), .B(n647), .Z(n648) );
  NOR2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n651), .A2(n650), .ZN(G305) );
  NAND2_X1 U725 ( .A1(n652), .A2(n655), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n653), .B(KEYINPUT84), .ZN(n664) );
  XOR2_X1 U727 ( .A(G299), .B(G288), .Z(n654) );
  XNOR2_X1 U728 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U729 ( .A(KEYINPUT19), .B(n656), .ZN(n658) );
  XNOR2_X1 U730 ( .A(G290), .B(KEYINPUT83), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n659), .B(G303), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n660), .B(G305), .ZN(n890) );
  XOR2_X1 U734 ( .A(n890), .B(n661), .Z(n662) );
  NAND2_X1 U735 ( .A1(G868), .A2(n662), .ZN(n663) );
  NAND2_X1 U736 ( .A1(n664), .A2(n663), .ZN(G295) );
  XOR2_X1 U737 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n668) );
  NAND2_X1 U738 ( .A1(G2084), .A2(G2078), .ZN(n665) );
  XOR2_X1 U739 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U740 ( .A1(n666), .A2(G2090), .ZN(n667) );
  XNOR2_X1 U741 ( .A(n668), .B(n667), .ZN(n669) );
  NAND2_X1 U742 ( .A1(G2072), .A2(n669), .ZN(G158) );
  XNOR2_X1 U743 ( .A(KEYINPUT86), .B(G44), .ZN(n670) );
  XNOR2_X1 U744 ( .A(n670), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U745 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  NOR2_X1 U746 ( .A1(G220), .A2(G219), .ZN(n671) );
  XOR2_X1 U747 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U748 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U749 ( .A1(G96), .A2(n673), .ZN(n822) );
  NAND2_X1 U750 ( .A1(G2106), .A2(n822), .ZN(n678) );
  NAND2_X1 U751 ( .A1(G69), .A2(G120), .ZN(n674) );
  NOR2_X1 U752 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U753 ( .A1(n675), .A2(G108), .ZN(n676) );
  XOR2_X1 U754 ( .A(KEYINPUT87), .B(n676), .Z(n823) );
  NAND2_X1 U755 ( .A1(G567), .A2(n823), .ZN(n677) );
  NAND2_X1 U756 ( .A1(n678), .A2(n677), .ZN(n824) );
  NAND2_X1 U757 ( .A1(G483), .A2(G661), .ZN(n679) );
  NOR2_X1 U758 ( .A1(n824), .A2(n679), .ZN(n821) );
  NAND2_X1 U759 ( .A1(n821), .A2(G36), .ZN(G176) );
  INV_X1 U760 ( .A(G301), .ZN(G171) );
  NAND2_X1 U761 ( .A1(G160), .A2(G40), .ZN(n751) );
  INV_X1 U762 ( .A(n751), .ZN(n680) );
  NAND2_X1 U763 ( .A1(n680), .A2(n752), .ZN(n681) );
  XNOR2_X2 U764 ( .A(n681), .B(KEYINPUT64), .ZN(n724) );
  INV_X1 U765 ( .A(G1996), .ZN(n931) );
  NOR2_X1 U766 ( .A1(n724), .A2(n931), .ZN(n683) );
  XNOR2_X1 U767 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n682) );
  XNOR2_X1 U768 ( .A(n683), .B(n682), .ZN(n685) );
  NOR2_X1 U769 ( .A1(n511), .A2(n979), .ZN(n684) );
  NOR2_X1 U770 ( .A1(n687), .A2(n981), .ZN(n686) );
  XOR2_X1 U771 ( .A(n686), .B(KEYINPUT98), .Z(n699) );
  NAND2_X1 U772 ( .A1(n687), .A2(n981), .ZN(n691) );
  NOR2_X1 U773 ( .A1(G2067), .A2(n724), .ZN(n689) );
  INV_X1 U774 ( .A(n724), .ZN(n709) );
  NOR2_X1 U775 ( .A1(G1348), .A2(n709), .ZN(n688) );
  NOR2_X1 U776 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U777 ( .A1(n691), .A2(n690), .ZN(n697) );
  INV_X1 U778 ( .A(G2072), .ZN(n930) );
  NOR2_X1 U779 ( .A1(n724), .A2(n930), .ZN(n693) );
  XOR2_X1 U780 ( .A(KEYINPUT97), .B(KEYINPUT27), .Z(n692) );
  XNOR2_X1 U781 ( .A(n693), .B(n692), .ZN(n695) );
  NAND2_X1 U782 ( .A1(n724), .A2(G1956), .ZN(n694) );
  NAND2_X1 U783 ( .A1(n695), .A2(n694), .ZN(n701) );
  NAND2_X1 U784 ( .A1(G299), .A2(n701), .ZN(n696) );
  XNOR2_X1 U785 ( .A(n696), .B(KEYINPUT28), .ZN(n700) );
  AND2_X1 U786 ( .A1(n697), .A2(n700), .ZN(n698) );
  NAND2_X1 U787 ( .A1(n699), .A2(n698), .ZN(n706) );
  INV_X1 U788 ( .A(n700), .ZN(n704) );
  NOR2_X1 U789 ( .A1(G299), .A2(n701), .ZN(n702) );
  XNOR2_X1 U790 ( .A(n702), .B(KEYINPUT99), .ZN(n703) );
  OR2_X1 U791 ( .A1(n704), .A2(n703), .ZN(n705) );
  AND2_X1 U792 ( .A1(n706), .A2(n705), .ZN(n708) );
  XNOR2_X1 U793 ( .A(n708), .B(n707), .ZN(n713) );
  XNOR2_X1 U794 ( .A(G2078), .B(KEYINPUT25), .ZN(n929) );
  NAND2_X1 U795 ( .A1(n709), .A2(n929), .ZN(n711) );
  INV_X1 U796 ( .A(G1961), .ZN(n952) );
  NAND2_X1 U797 ( .A1(n724), .A2(n952), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U799 ( .A1(n714), .A2(G171), .ZN(n712) );
  NAND2_X1 U800 ( .A1(n713), .A2(n712), .ZN(n723) );
  NOR2_X1 U801 ( .A1(G171), .A2(n714), .ZN(n719) );
  NAND2_X1 U802 ( .A1(n724), .A2(G8), .ZN(n808) );
  NOR2_X1 U803 ( .A1(G1966), .A2(n808), .ZN(n735) );
  NOR2_X1 U804 ( .A1(n724), .A2(G2084), .ZN(n732) );
  NOR2_X1 U805 ( .A1(n735), .A2(n732), .ZN(n715) );
  NAND2_X1 U806 ( .A1(G8), .A2(n715), .ZN(n716) );
  XNOR2_X1 U807 ( .A(KEYINPUT30), .B(n716), .ZN(n717) );
  NOR2_X1 U808 ( .A1(G168), .A2(n717), .ZN(n718) );
  NOR2_X1 U809 ( .A1(n719), .A2(n718), .ZN(n721) );
  XOR2_X1 U810 ( .A(KEYINPUT31), .B(KEYINPUT100), .Z(n720) );
  XNOR2_X1 U811 ( .A(n721), .B(n720), .ZN(n722) );
  NAND2_X1 U812 ( .A1(n723), .A2(n722), .ZN(n733) );
  NAND2_X1 U813 ( .A1(n733), .A2(G286), .ZN(n729) );
  NOR2_X1 U814 ( .A1(n724), .A2(G2090), .ZN(n726) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n808), .ZN(n725) );
  NOR2_X1 U816 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U817 ( .A1(n727), .A2(G303), .ZN(n728) );
  NAND2_X1 U818 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U819 ( .A1(n730), .A2(G8), .ZN(n731) );
  XNOR2_X1 U820 ( .A(KEYINPUT32), .B(n731), .ZN(n739) );
  NAND2_X1 U821 ( .A1(G8), .A2(n732), .ZN(n737) );
  XNOR2_X1 U822 ( .A(KEYINPUT101), .B(n733), .ZN(n734) );
  NOR2_X1 U823 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U824 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U825 ( .A1(n739), .A2(n738), .ZN(n804) );
  NOR2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n746) );
  NOR2_X1 U827 ( .A1(G1971), .A2(G303), .ZN(n740) );
  NOR2_X1 U828 ( .A1(n746), .A2(n740), .ZN(n986) );
  NAND2_X1 U829 ( .A1(n804), .A2(n986), .ZN(n743) );
  INV_X1 U830 ( .A(n808), .ZN(n741) );
  NAND2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n985) );
  AND2_X1 U832 ( .A1(n741), .A2(n985), .ZN(n742) );
  AND2_X1 U833 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U834 ( .A1(KEYINPUT33), .A2(n744), .ZN(n745) );
  XNOR2_X1 U835 ( .A(n745), .B(KEYINPUT102), .ZN(n749) );
  NAND2_X1 U836 ( .A1(n746), .A2(KEYINPUT33), .ZN(n747) );
  NOR2_X1 U837 ( .A1(n808), .A2(n747), .ZN(n748) );
  NOR2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n787) );
  XNOR2_X1 U839 ( .A(G1981), .B(KEYINPUT103), .ZN(n750) );
  XNOR2_X1 U840 ( .A(n750), .B(G305), .ZN(n976) );
  NOR2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n799) );
  NAND2_X1 U842 ( .A1(G140), .A2(n867), .ZN(n754) );
  NAND2_X1 U843 ( .A1(G104), .A2(n868), .ZN(n753) );
  NAND2_X1 U844 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U845 ( .A(KEYINPUT34), .B(n755), .ZN(n760) );
  NAND2_X1 U846 ( .A1(G116), .A2(n871), .ZN(n757) );
  NAND2_X1 U847 ( .A1(G128), .A2(n872), .ZN(n756) );
  NAND2_X1 U848 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U849 ( .A(KEYINPUT35), .B(n758), .Z(n759) );
  NOR2_X1 U850 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U851 ( .A(KEYINPUT36), .B(n761), .ZN(n886) );
  XNOR2_X1 U852 ( .A(G2067), .B(KEYINPUT37), .ZN(n788) );
  NOR2_X1 U853 ( .A1(n886), .A2(n788), .ZN(n908) );
  NAND2_X1 U854 ( .A1(n799), .A2(n908), .ZN(n762) );
  XNOR2_X1 U855 ( .A(n762), .B(KEYINPUT90), .ZN(n795) );
  XNOR2_X1 U856 ( .A(G1986), .B(G290), .ZN(n994) );
  NAND2_X1 U857 ( .A1(n994), .A2(n799), .ZN(n763) );
  XOR2_X1 U858 ( .A(KEYINPUT89), .B(n763), .Z(n764) );
  NAND2_X1 U859 ( .A1(n795), .A2(n764), .ZN(n785) );
  NAND2_X1 U860 ( .A1(n868), .A2(G105), .ZN(n765) );
  XNOR2_X1 U861 ( .A(n765), .B(KEYINPUT38), .ZN(n767) );
  NAND2_X1 U862 ( .A1(G117), .A2(n871), .ZN(n766) );
  NAND2_X1 U863 ( .A1(n767), .A2(n766), .ZN(n770) );
  NAND2_X1 U864 ( .A1(G129), .A2(n872), .ZN(n768) );
  XNOR2_X1 U865 ( .A(KEYINPUT93), .B(n768), .ZN(n769) );
  NOR2_X1 U866 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U867 ( .A(KEYINPUT94), .B(n771), .ZN(n774) );
  NAND2_X1 U868 ( .A1(n867), .A2(G141), .ZN(n772) );
  XOR2_X1 U869 ( .A(KEYINPUT95), .B(n772), .Z(n773) );
  NAND2_X1 U870 ( .A1(n774), .A2(n773), .ZN(n855) );
  NAND2_X1 U871 ( .A1(G1996), .A2(n855), .ZN(n775) );
  XNOR2_X1 U872 ( .A(n775), .B(KEYINPUT96), .ZN(n784) );
  XNOR2_X1 U873 ( .A(KEYINPUT92), .B(G1991), .ZN(n934) );
  NAND2_X1 U874 ( .A1(G107), .A2(n871), .ZN(n777) );
  NAND2_X1 U875 ( .A1(G95), .A2(n868), .ZN(n776) );
  NAND2_X1 U876 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U877 ( .A1(G131), .A2(n867), .ZN(n778) );
  XNOR2_X1 U878 ( .A(KEYINPUT91), .B(n778), .ZN(n779) );
  NOR2_X1 U879 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U880 ( .A1(n872), .A2(G119), .ZN(n781) );
  NAND2_X1 U881 ( .A1(n782), .A2(n781), .ZN(n856) );
  NAND2_X1 U882 ( .A1(n934), .A2(n856), .ZN(n783) );
  NAND2_X1 U883 ( .A1(n784), .A2(n783), .ZN(n924) );
  AND2_X1 U884 ( .A1(n799), .A2(n924), .ZN(n791) );
  NOR2_X1 U885 ( .A1(n785), .A2(n791), .ZN(n801) );
  AND2_X1 U886 ( .A1(n976), .A2(n801), .ZN(n786) );
  NAND2_X1 U887 ( .A1(n787), .A2(n786), .ZN(n816) );
  NAND2_X1 U888 ( .A1(n886), .A2(n788), .ZN(n914) );
  NOR2_X1 U889 ( .A1(G1996), .A2(n855), .ZN(n917) );
  NOR2_X1 U890 ( .A1(G1986), .A2(G290), .ZN(n789) );
  NOR2_X1 U891 ( .A1(n934), .A2(n856), .ZN(n913) );
  NOR2_X1 U892 ( .A1(n789), .A2(n913), .ZN(n790) );
  NOR2_X1 U893 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U894 ( .A(n792), .B(KEYINPUT104), .ZN(n793) );
  NOR2_X1 U895 ( .A1(n917), .A2(n793), .ZN(n794) );
  XNOR2_X1 U896 ( .A(KEYINPUT39), .B(n794), .ZN(n796) );
  NAND2_X1 U897 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U898 ( .A1(n914), .A2(n797), .ZN(n798) );
  NAND2_X1 U899 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U900 ( .A(KEYINPUT105), .B(n800), .Z(n814) );
  INV_X1 U901 ( .A(n801), .ZN(n812) );
  NOR2_X1 U902 ( .A1(G2090), .A2(G303), .ZN(n802) );
  NAND2_X1 U903 ( .A1(G8), .A2(n802), .ZN(n803) );
  NAND2_X1 U904 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U905 ( .A1(n805), .A2(n808), .ZN(n810) );
  NOR2_X1 U906 ( .A1(G1981), .A2(G305), .ZN(n806) );
  XOR2_X1 U907 ( .A(n806), .B(KEYINPUT24), .Z(n807) );
  OR2_X1 U908 ( .A1(n808), .A2(n807), .ZN(n809) );
  AND2_X1 U909 ( .A1(n810), .A2(n809), .ZN(n811) );
  OR2_X1 U910 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U911 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U912 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U913 ( .A(n817), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n818), .ZN(G217) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n819) );
  NAND2_X1 U916 ( .A1(G661), .A2(n819), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n820) );
  NAND2_X1 U918 ( .A1(n821), .A2(n820), .ZN(G188) );
  XNOR2_X1 U919 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  XOR2_X1 U920 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  INV_X1 U922 ( .A(G108), .ZN(G238) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  NOR2_X1 U924 ( .A1(n823), .A2(n822), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U926 ( .A(KEYINPUT109), .B(n824), .ZN(G319) );
  XOR2_X1 U927 ( .A(KEYINPUT43), .B(KEYINPUT111), .Z(n826) );
  XNOR2_X1 U928 ( .A(G2100), .B(KEYINPUT110), .ZN(n825) );
  XNOR2_X1 U929 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U930 ( .A(n827), .B(G2096), .Z(n829) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2072), .ZN(n828) );
  XNOR2_X1 U932 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U933 ( .A(KEYINPUT42), .B(G2090), .Z(n831) );
  XNOR2_X1 U934 ( .A(G2084), .B(G2078), .ZN(n830) );
  XNOR2_X1 U935 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U936 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U937 ( .A(G2678), .B(KEYINPUT112), .ZN(n834) );
  XNOR2_X1 U938 ( .A(n835), .B(n834), .ZN(G227) );
  XOR2_X1 U939 ( .A(G1976), .B(G1971), .Z(n837) );
  XNOR2_X1 U940 ( .A(G1966), .B(G1961), .ZN(n836) );
  XNOR2_X1 U941 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U942 ( .A(G1981), .B(G1956), .Z(n839) );
  XNOR2_X1 U943 ( .A(G1991), .B(G1996), .ZN(n838) );
  XNOR2_X1 U944 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U945 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U946 ( .A(KEYINPUT113), .B(G2474), .ZN(n842) );
  XNOR2_X1 U947 ( .A(n843), .B(n842), .ZN(n845) );
  XOR2_X1 U948 ( .A(G1986), .B(KEYINPUT41), .Z(n844) );
  XNOR2_X1 U949 ( .A(n845), .B(n844), .ZN(G229) );
  NAND2_X1 U950 ( .A1(G100), .A2(n868), .ZN(n846) );
  XNOR2_X1 U951 ( .A(n846), .B(KEYINPUT114), .ZN(n853) );
  NAND2_X1 U952 ( .A1(G136), .A2(n867), .ZN(n848) );
  NAND2_X1 U953 ( .A1(G112), .A2(n871), .ZN(n847) );
  NAND2_X1 U954 ( .A1(n848), .A2(n847), .ZN(n851) );
  NAND2_X1 U955 ( .A1(n872), .A2(G124), .ZN(n849) );
  XOR2_X1 U956 ( .A(KEYINPUT44), .B(n849), .Z(n850) );
  NOR2_X1 U957 ( .A1(n851), .A2(n850), .ZN(n852) );
  NAND2_X1 U958 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U959 ( .A(KEYINPUT115), .B(n854), .ZN(G162) );
  XOR2_X1 U960 ( .A(n856), .B(n855), .Z(n857) );
  XNOR2_X1 U961 ( .A(G164), .B(n857), .ZN(n866) );
  NAND2_X1 U962 ( .A1(G118), .A2(n871), .ZN(n859) );
  NAND2_X1 U963 ( .A1(G130), .A2(n872), .ZN(n858) );
  NAND2_X1 U964 ( .A1(n859), .A2(n858), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G142), .A2(n867), .ZN(n861) );
  NAND2_X1 U966 ( .A1(G106), .A2(n868), .ZN(n860) );
  NAND2_X1 U967 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U968 ( .A(KEYINPUT45), .B(n862), .Z(n863) );
  NOR2_X1 U969 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U970 ( .A(n866), .B(n865), .Z(n879) );
  NAND2_X1 U971 ( .A1(G139), .A2(n867), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G103), .A2(n868), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n877) );
  NAND2_X1 U974 ( .A1(G115), .A2(n871), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G127), .A2(n872), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n903) );
  XNOR2_X1 U979 ( .A(G160), .B(n903), .ZN(n878) );
  XNOR2_X1 U980 ( .A(n879), .B(n878), .ZN(n888) );
  XNOR2_X1 U981 ( .A(KEYINPUT46), .B(KEYINPUT118), .ZN(n881) );
  XNOR2_X1 U982 ( .A(n910), .B(KEYINPUT117), .ZN(n880) );
  XNOR2_X1 U983 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U984 ( .A(n882), .B(KEYINPUT116), .Z(n884) );
  XNOR2_X1 U985 ( .A(G162), .B(KEYINPUT48), .ZN(n883) );
  XNOR2_X1 U986 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U987 ( .A(n886), .B(n885), .Z(n887) );
  XNOR2_X1 U988 ( .A(n888), .B(n887), .ZN(n889) );
  NOR2_X1 U989 ( .A1(G37), .A2(n889), .ZN(G395) );
  XOR2_X1 U990 ( .A(KEYINPUT119), .B(n890), .Z(n892) );
  XNOR2_X1 U991 ( .A(G171), .B(G286), .ZN(n891) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n979), .B(n981), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U995 ( .A1(G37), .A2(n895), .ZN(G397) );
  NOR2_X1 U996 ( .A1(G227), .A2(G229), .ZN(n897) );
  XNOR2_X1 U997 ( .A(KEYINPUT49), .B(KEYINPUT120), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U999 ( .A1(G401), .A2(n898), .ZN(n899) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n899), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(KEYINPUT121), .B(n900), .ZN(n902) );
  NOR2_X1 U1002 ( .A1(G395), .A2(G397), .ZN(n901) );
  NAND2_X1 U1003 ( .A1(n902), .A2(n901), .ZN(G225) );
  INV_X1 U1004 ( .A(G225), .ZN(G308) );
  INV_X1 U1005 ( .A(G303), .ZN(G166) );
  XOR2_X1 U1006 ( .A(G2072), .B(n903), .Z(n905) );
  XOR2_X1 U1007 ( .A(G164), .B(G2078), .Z(n904) );
  NOR2_X1 U1008 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1009 ( .A(KEYINPUT50), .B(n906), .Z(n907) );
  NOR2_X1 U1010 ( .A1(n908), .A2(n907), .ZN(n922) );
  XNOR2_X1 U1011 ( .A(G160), .B(G2084), .ZN(n909) );
  XNOR2_X1 U1012 ( .A(n909), .B(KEYINPUT122), .ZN(n911) );
  NAND2_X1 U1013 ( .A1(n911), .A2(n910), .ZN(n912) );
  NOR2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n915), .A2(n914), .ZN(n920) );
  XOR2_X1 U1016 ( .A(G2090), .B(G162), .Z(n916) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n918), .B(KEYINPUT51), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(KEYINPUT52), .B(n925), .ZN(n926) );
  INV_X1 U1023 ( .A(KEYINPUT55), .ZN(n948) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n948), .ZN(n927) );
  NAND2_X1 U1025 ( .A1(n927), .A2(G29), .ZN(n1008) );
  XNOR2_X1 U1026 ( .A(G2090), .B(G35), .ZN(n943) );
  XOR2_X1 U1027 ( .A(G2067), .B(G26), .Z(n928) );
  NAND2_X1 U1028 ( .A1(n928), .A2(G28), .ZN(n940) );
  XNOR2_X1 U1029 ( .A(G27), .B(n929), .ZN(n938) );
  XNOR2_X1 U1030 ( .A(n930), .B(G33), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(n931), .B(G32), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(G25), .B(n934), .ZN(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1037 ( .A(KEYINPUT53), .B(n941), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n946) );
  XOR2_X1 U1039 ( .A(G2084), .B(G34), .Z(n944) );
  XNOR2_X1 U1040 ( .A(KEYINPUT54), .B(n944), .ZN(n945) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(n948), .B(n947), .ZN(n950) );
  INV_X1 U1043 ( .A(G29), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1045 ( .A1(G11), .A2(n951), .ZN(n1006) );
  XNOR2_X1 U1046 ( .A(G5), .B(n952), .ZN(n962) );
  XNOR2_X1 U1047 ( .A(G1971), .B(G22), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G23), .B(G1976), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1050 ( .A(KEYINPUT126), .B(n955), .Z(n957) );
  XNOR2_X1 U1051 ( .A(G1986), .B(G24), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1053 ( .A(KEYINPUT58), .B(n958), .Z(n960) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G21), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n972) );
  XOR2_X1 U1057 ( .A(G1348), .B(KEYINPUT59), .Z(n963) );
  XNOR2_X1 U1058 ( .A(G4), .B(n963), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(G20), .B(G1956), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(G1341), .B(G19), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(G1981), .B(G6), .ZN(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(KEYINPUT60), .B(n970), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1067 ( .A(KEYINPUT61), .B(n973), .Z(n974) );
  NOR2_X1 U1068 ( .A1(G16), .A2(n974), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(KEYINPUT127), .B(n975), .ZN(n1004) );
  XNOR2_X1 U1070 ( .A(KEYINPUT56), .B(G16), .ZN(n1002) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G168), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(n978), .B(KEYINPUT57), .ZN(n1000) );
  XNOR2_X1 U1074 ( .A(G1341), .B(KEYINPUT125), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(n980), .B(n979), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(G1348), .B(n981), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n998) );
  XNOR2_X1 U1078 ( .A(G299), .B(G1956), .ZN(n991) );
  INV_X1 U1079 ( .A(G1971), .ZN(n984) );
  NOR2_X1 U1080 ( .A1(G166), .A2(n984), .ZN(n988) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(KEYINPUT123), .B(n989), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(KEYINPUT124), .B(n992), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(G1961), .B(G301), .ZN(n993) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1095 ( .A(KEYINPUT62), .B(n1009), .Z(G311) );
  INV_X1 U1096 ( .A(G311), .ZN(G150) );
endmodule

