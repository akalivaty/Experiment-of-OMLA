//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1213,
    new_n1214, new_n1215, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  INV_X1    g0005(.A(G58), .ZN(new_n206));
  INV_X1    g0006(.A(G232), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  INV_X1    g0008(.A(G264), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G50), .B2(G226), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(KEYINPUT64), .ZN(new_n214));
  AND2_X1   g0014(.A1(new_n213), .A2(KEYINPUT64), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n211), .B(new_n212), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n205), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  NAND2_X1  g0022(.A1(new_n202), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n205), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT0), .ZN(new_n232));
  NAND4_X1  g0032(.A1(new_n222), .A2(new_n228), .A3(new_n229), .A4(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n245), .B(KEYINPUT67), .Z(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT66), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G68), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n246), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OR2_X1    g0054(.A1(new_n254), .A2(KEYINPUT68), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n254), .A2(KEYINPUT68), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n255), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n256), .A2(new_n254), .ZN(new_n261));
  INV_X1    g0061(.A(G226), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT69), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n262), .A2(KEYINPUT69), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT70), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G222), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G223), .A2(G1698), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n276), .B(new_n256), .C1(G77), .C2(new_n272), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n267), .A2(G190), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT75), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n267), .A2(new_n277), .ZN(new_n280));
  INV_X1    g0080(.A(G200), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n278), .B(new_n279), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n225), .ZN(new_n284));
  INV_X1    g0084(.A(G50), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n226), .B1(new_n201), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n286), .B(KEYINPUT72), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT71), .B1(G20), .B2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NOR3_X1   g0089(.A1(KEYINPUT71), .A2(G20), .A3(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G150), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n226), .A2(G33), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n291), .A2(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n284), .B1(new_n287), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G1), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(G13), .A3(G20), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n285), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n284), .B1(new_n297), .B2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G50), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n296), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OR3_X1    g0104(.A1(new_n304), .A2(KEYINPUT74), .A3(KEYINPUT9), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT74), .B1(new_n304), .B2(KEYINPUT9), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n282), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n304), .A2(KEYINPUT9), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n307), .A2(new_n312), .A3(new_n309), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n280), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n316), .B(new_n303), .C1(G169), .C2(new_n280), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n261), .A2(G238), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n207), .A2(G1698), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n272), .B(new_n319), .C1(G226), .C2(G1698), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G97), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n256), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n260), .B(new_n318), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT13), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n323), .B1(new_n320), .B2(new_n321), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n255), .A2(new_n258), .A3(new_n259), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT13), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(new_n318), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G169), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n332), .A2(KEYINPUT14), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n331), .A2(new_n315), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n332), .A2(KEYINPUT14), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n291), .ZN(new_n338));
  INV_X1    g0138(.A(G68), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n338), .A2(G50), .B1(G20), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n217), .B2(new_n294), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n284), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT11), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n299), .A2(new_n339), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT12), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n341), .A2(KEYINPUT11), .A3(new_n284), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n301), .A2(G68), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n344), .A2(new_n346), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n331), .A2(G200), .ZN(new_n350));
  INV_X1    g0150(.A(new_n331), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n349), .B1(new_n351), .B2(G190), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n337), .A2(new_n349), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n269), .A2(new_n271), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G107), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n207), .A2(G1698), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(G238), .B2(G1698), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n355), .B1(new_n357), .B2(new_n354), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT73), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n256), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n327), .B1(G244), .B2(new_n261), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(G169), .ZN(new_n364));
  INV_X1    g0164(.A(new_n293), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n338), .A2(new_n365), .B1(G20), .B2(G77), .ZN(new_n366));
  XOR2_X1   g0166(.A(KEYINPUT15), .B(G87), .Z(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n366), .B1(new_n294), .B2(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(new_n284), .B1(new_n217), .B2(new_n299), .ZN(new_n370));
  INV_X1    g0170(.A(new_n301), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(new_n217), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n362), .B2(G179), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n364), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n314), .A2(new_n317), .A3(new_n353), .A4(new_n375), .ZN(new_n376));
  XNOR2_X1  g0176(.A(G58), .B(G68), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G20), .ZN(new_n378));
  INV_X1    g0178(.A(G159), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n378), .B1(new_n291), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n270), .A2(KEYINPUT76), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT76), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G33), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n384), .A3(KEYINPUT3), .ZN(new_n385));
  AOI21_X1  g0185(.A(G20), .B1(new_n385), .B2(new_n269), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT7), .ZN(new_n387));
  OAI21_X1  g0187(.A(G68), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n269), .ZN(new_n389));
  XNOR2_X1  g0189(.A(KEYINPUT76), .B(G33), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n389), .B1(new_n390), .B2(KEYINPUT3), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n391), .A2(KEYINPUT7), .A3(G20), .ZN(new_n392));
  OAI211_X1 g0192(.A(KEYINPUT16), .B(new_n381), .C1(new_n388), .C2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n387), .B1(new_n272), .B2(G20), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n382), .A2(new_n384), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(KEYINPUT77), .A3(new_n268), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n226), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT3), .B1(new_n382), .B2(new_n384), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT77), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n271), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT7), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n394), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n380), .B1(new_n402), .B2(G68), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n284), .B(new_n393), .C1(new_n403), .C2(KEYINPUT16), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n293), .A2(new_n298), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n301), .B2(new_n293), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n262), .A2(G1698), .ZN(new_n407));
  OR2_X1    g0207(.A1(G223), .A2(G1698), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n385), .A2(new_n407), .A3(new_n269), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G87), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n256), .ZN(new_n412));
  INV_X1    g0212(.A(G190), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n261), .A2(G232), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n412), .A2(new_n413), .A3(new_n414), .A4(new_n260), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n323), .B1(new_n409), .B2(new_n410), .ZN(new_n416));
  INV_X1    g0216(.A(new_n414), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n416), .A2(new_n327), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n415), .B1(new_n418), .B2(G200), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n404), .A2(new_n406), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT78), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT78), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n404), .A2(new_n422), .A3(new_n419), .A4(new_n406), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(KEYINPUT17), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n404), .A2(new_n406), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n418), .A2(G179), .ZN(new_n430));
  INV_X1    g0230(.A(G169), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n430), .B1(new_n431), .B2(new_n418), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n429), .A2(KEYINPUT18), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT18), .B1(new_n429), .B2(new_n432), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n372), .B1(new_n363), .B2(G190), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n281), .B2(new_n363), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n428), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n376), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n284), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n297), .A2(G33), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n298), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT79), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n444), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G107), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n299), .A2(new_n208), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n448), .B1(KEYINPUT25), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G87), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G20), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n385), .A2(KEYINPUT22), .A3(new_n269), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G116), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(new_n382), .B2(new_n384), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n226), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n208), .A2(G20), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT23), .ZN(new_n458));
  XNOR2_X1  g0258(.A(new_n457), .B(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n452), .A2(new_n269), .A3(new_n271), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT22), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n453), .A2(new_n456), .A3(new_n459), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT85), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT24), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n226), .A2(new_n455), .B1(new_n460), .B2(new_n461), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT85), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n466), .A2(new_n467), .A3(new_n459), .A4(new_n453), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n464), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n465), .B1(new_n464), .B2(new_n468), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n284), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT86), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(KEYINPUT86), .B(new_n284), .C1(new_n469), .C2(new_n470), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n450), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n449), .A2(KEYINPUT25), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n391), .A2(KEYINPUT87), .A3(G257), .A4(G1698), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n385), .A2(G257), .A3(G1698), .A4(new_n269), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT87), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n385), .A2(G250), .A3(new_n273), .A4(new_n269), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n395), .A2(G294), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT88), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT88), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n482), .A2(new_n488), .A3(new_n485), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n256), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n253), .A2(G1), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT81), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n492), .B(new_n493), .C1(KEYINPUT5), .C2(new_n252), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n297), .A2(G45), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT81), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n258), .A2(new_n491), .A3(new_n494), .A4(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n497), .A3(new_n491), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n323), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(new_n209), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n490), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n431), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n490), .A2(new_n502), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(new_n315), .A3(new_n498), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n477), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(G190), .A3(new_n498), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n503), .A2(G200), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n475), .A2(new_n508), .A3(new_n509), .A4(new_n476), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n209), .A2(G1698), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n391), .B(new_n512), .C1(G257), .C2(G1698), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n354), .A2(G303), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n323), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n499), .A2(G270), .A3(new_n323), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n498), .ZN(new_n517));
  OR2_X1    g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OR2_X1    g0318(.A1(new_n443), .A2(new_n454), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n299), .A2(new_n454), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  INV_X1    g0321(.A(G97), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n226), .C1(G33), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n454), .A2(G20), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n284), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT20), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n525), .A2(new_n526), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n519), .B(new_n520), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n518), .A2(new_n531), .A3(new_n315), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(G169), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n515), .A2(new_n517), .ZN(new_n534));
  OAI211_X1 g0334(.A(KEYINPUT84), .B(KEYINPUT21), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n529), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n536), .A2(new_n527), .B1(new_n454), .B2(new_n299), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n431), .B1(new_n537), .B2(new_n519), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT84), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT21), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n540), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n518), .A2(new_n538), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n532), .B1(new_n535), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n256), .B1(new_n257), .B2(new_n492), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n492), .A2(G250), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G238), .A2(G1698), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n218), .B2(G1698), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n455), .B1(new_n391), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n548), .B1(new_n551), .B2(new_n323), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G200), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n367), .A2(new_n298), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n391), .A2(new_n226), .A3(G68), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT19), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n556), .A2(new_n226), .A3(G33), .A4(G97), .ZN(new_n557));
  NOR3_X1   g0357(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n226), .B2(new_n321), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n557), .B1(new_n559), .B2(new_n556), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n554), .B1(new_n561), .B2(new_n284), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n445), .A2(G87), .A3(new_n446), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n553), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT83), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n552), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G190), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n553), .A2(new_n562), .A3(KEYINPUT83), .A4(new_n563), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n447), .A2(new_n367), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n562), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT82), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n567), .A2(G179), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n567), .B2(new_n431), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n571), .A2(KEYINPUT82), .A3(new_n562), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n534), .A2(G190), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n579), .B(new_n531), .C1(new_n281), .C2(new_n534), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n545), .A2(new_n570), .A3(new_n578), .A4(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n391), .A2(G244), .A3(new_n273), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT4), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n272), .A2(G250), .A3(G1698), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n583), .A2(G1698), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n586), .A2(new_n269), .A3(new_n271), .A4(G244), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n587), .B(KEYINPUT80), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n584), .A2(new_n585), .A3(new_n588), .A4(new_n521), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n256), .ZN(new_n590));
  INV_X1    g0390(.A(G257), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n500), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n498), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G200), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT6), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n522), .A2(new_n208), .ZN(new_n597));
  NOR2_X1   g0397(.A1(G97), .A2(G107), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n208), .A2(KEYINPUT6), .A3(G97), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n226), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n402), .B2(G107), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n217), .B2(new_n291), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n603), .A2(new_n284), .B1(new_n522), .B2(new_n299), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n447), .A2(G97), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n590), .A2(G190), .A3(new_n498), .A4(new_n593), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n595), .A2(new_n604), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n291), .A2(new_n217), .ZN(new_n608));
  AOI211_X1 g0408(.A(new_n608), .B(new_n601), .C1(new_n402), .C2(G107), .ZN(new_n609));
  OAI221_X1 g0409(.A(new_n605), .B1(G97), .B2(new_n298), .C1(new_n609), .C2(new_n441), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n594), .A2(new_n431), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n590), .A2(new_n315), .A3(new_n498), .A4(new_n593), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n581), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n440), .A2(new_n511), .A3(new_n615), .ZN(G372));
  AND2_X1   g0416(.A1(new_n337), .A2(new_n349), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n375), .B1(new_n350), .B2(new_n352), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n428), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n436), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n314), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT90), .B1(new_n621), .B2(new_n317), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT90), .ZN(new_n623));
  INV_X1    g0423(.A(new_n317), .ZN(new_n624));
  AOI211_X1 g0424(.A(new_n623), .B(new_n624), .C1(new_n620), .C2(new_n314), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n576), .A2(new_n572), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n578), .A2(new_n570), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT26), .B1(new_n628), .B2(new_n613), .ZN(new_n629));
  INV_X1    g0429(.A(new_n545), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n475), .A2(new_n476), .B1(new_n431), .B2(new_n503), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n630), .B1(new_n631), .B2(new_n506), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n562), .A2(KEYINPUT89), .A3(new_n563), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT89), .B1(new_n562), .B2(new_n563), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n568), .B(new_n553), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n607), .A2(new_n613), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n510), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n627), .B(new_n629), .C1(new_n632), .C2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n635), .A2(new_n611), .A3(new_n610), .A4(new_n612), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n440), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n626), .A2(new_n642), .ZN(G369));
  INV_X1    g0443(.A(new_n477), .ZN(new_n644));
  INV_X1    g0444(.A(G13), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(G20), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n297), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n511), .B1(new_n644), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n507), .B2(new_n653), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n531), .A2(new_n653), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n630), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n545), .A2(new_n580), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n657), .B1(new_n658), .B2(new_n656), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n545), .A2(new_n652), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n511), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g0464(.A(new_n652), .B(KEYINPUT91), .Z(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n631), .A2(new_n506), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n662), .A2(new_n668), .ZN(G399));
  INV_X1    g0469(.A(new_n230), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G41), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n558), .A2(new_n454), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n671), .A2(new_n672), .A3(new_n297), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT92), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  INV_X1    g0476(.A(new_n671), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n675), .B(new_n676), .C1(new_n223), .C2(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT29), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n641), .A2(new_n680), .A3(new_n666), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n628), .A2(new_n613), .A3(KEYINPUT26), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n627), .B(new_n684), .C1(new_n632), .C2(new_n637), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n653), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT29), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n615), .A2(new_n507), .A3(new_n510), .A4(new_n666), .ZN(new_n689));
  INV_X1    g0489(.A(new_n498), .ZN(new_n690));
  AOI211_X1 g0490(.A(new_n690), .B(new_n592), .C1(new_n589), .C2(new_n256), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n691), .A2(G179), .A3(new_n534), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(new_n503), .A3(new_n552), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n518), .A2(new_n575), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n694), .A2(new_n691), .A3(new_n502), .A4(new_n490), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n505), .A2(KEYINPUT30), .A3(new_n691), .A4(new_n694), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n693), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n652), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n699), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n689), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n688), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n679), .B1(new_n707), .B2(G1), .ZN(G364));
  NOR2_X1   g0508(.A1(new_n226), .A2(G190), .ZN(new_n709));
  NOR2_X1   g0509(.A1(G179), .A2(G200), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n379), .ZN(new_n712));
  XOR2_X1   g0512(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n713));
  XNOR2_X1  g0513(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n226), .A2(new_n413), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n315), .A2(G200), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n709), .A2(new_n716), .ZN(new_n718));
  OAI221_X1 g0518(.A(new_n714), .B1(new_n206), .B2(new_n717), .C1(new_n217), .C2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n281), .A2(G179), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n451), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n226), .A2(new_n315), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G200), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n413), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n226), .B1(new_n710), .B2(G190), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n726), .A2(new_n285), .B1(new_n727), .B2(new_n522), .ZN(new_n728));
  NOR4_X1   g0528(.A1(new_n719), .A2(new_n354), .A3(new_n722), .A4(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n724), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n730), .A2(KEYINPUT97), .A3(new_n413), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT97), .B1(new_n730), .B2(new_n413), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n720), .A2(new_n709), .ZN(new_n734));
  OAI221_X1 g0534(.A(new_n729), .B1(new_n339), .B2(new_n733), .C1(new_n208), .C2(new_n734), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT98), .ZN(new_n736));
  INV_X1    g0536(.A(G294), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n354), .B1(new_n727), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G322), .ZN(new_n739));
  INV_X1    g0539(.A(G311), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n717), .A2(new_n739), .B1(new_n718), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n711), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n741), .B1(G329), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G283), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n743), .B1(new_n744), .B2(new_n734), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n738), .B(new_n745), .C1(G326), .C2(new_n725), .ZN(new_n746));
  INV_X1    g0546(.A(G303), .ZN(new_n747));
  XOR2_X1   g0547(.A(KEYINPUT33), .B(G317), .Z(new_n748));
  OAI221_X1 g0548(.A(new_n746), .B1(new_n747), .B2(new_n721), .C1(new_n733), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n736), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT99), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n225), .B1(G20), .B2(new_n431), .ZN(new_n752));
  INV_X1    g0552(.A(new_n391), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n230), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT93), .Z(new_n755));
  NAND2_X1  g0555(.A1(new_n224), .A2(new_n253), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n755), .B(new_n756), .C1(new_n250), .C2(new_n253), .ZN(new_n757));
  INV_X1    g0557(.A(G355), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n272), .A2(new_n230), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n757), .B1(G116), .B2(new_n230), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT94), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n752), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT95), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n751), .A2(new_n752), .B1(new_n762), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n297), .B1(new_n646), .B2(G45), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n671), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n766), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n770), .B(new_n773), .C1(new_n659), .C2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT100), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n661), .A2(new_n773), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G330), .B2(new_n659), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n776), .A2(new_n778), .ZN(G396));
  NAND2_X1  g0579(.A1(new_n641), .A2(new_n666), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n372), .A2(new_n652), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n438), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n375), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n374), .A2(new_n653), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n785), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n666), .B(new_n787), .C1(new_n638), .C2(new_n640), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n705), .ZN(new_n790));
  INV_X1    g0590(.A(new_n773), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n786), .A2(new_n706), .A3(new_n788), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n752), .ZN(new_n794));
  INV_X1    g0594(.A(new_n717), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n725), .A2(G137), .B1(new_n795), .B2(G143), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n796), .B1(new_n379), .B2(new_n718), .C1(new_n733), .C2(new_n292), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT34), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n742), .A2(G132), .ZN(new_n799));
  INV_X1    g0599(.A(new_n734), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G68), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n285), .B2(new_n721), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT101), .ZN(new_n803));
  INV_X1    g0603(.A(new_n727), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n753), .B1(G58), .B2(new_n804), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n798), .A2(new_n799), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n726), .A2(new_n747), .B1(new_n727), .B2(new_n522), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n717), .A2(new_n737), .B1(new_n718), .B2(new_n454), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n354), .B1(new_n721), .B2(new_n208), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n734), .A2(new_n451), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n807), .A2(new_n808), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n811), .B1(new_n744), .B2(new_n733), .C1(new_n740), .C2(new_n711), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n794), .B1(new_n806), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n752), .A2(new_n764), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n813), .B1(new_n217), .B2(new_n814), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n773), .B(new_n815), .C1(new_n787), .C2(new_n765), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n793), .A2(new_n816), .ZN(G384));
  INV_X1    g0617(.A(KEYINPUT105), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n424), .B(new_n426), .C1(new_n434), .C2(new_n433), .ZN(new_n819));
  INV_X1    g0619(.A(new_n650), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n429), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n421), .A2(new_n423), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT37), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n429), .A2(new_n432), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n823), .A2(new_n824), .A3(new_n825), .A4(new_n821), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(new_n821), .A3(new_n420), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(KEYINPUT37), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n819), .A2(new_n822), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n818), .B1(new_n829), .B2(KEYINPUT38), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n822), .B1(new_n427), .B2(new_n435), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n826), .A2(new_n828), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT38), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n833), .A2(KEYINPUT105), .A3(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT39), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n381), .B1(new_n388), .B2(new_n392), .ZN(new_n837));
  NOR2_X1   g0637(.A1(KEYINPUT103), .A2(KEYINPUT16), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n381), .B1(KEYINPUT103), .B2(KEYINPUT16), .C1(new_n388), .C2(new_n392), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n839), .A2(new_n840), .A3(new_n284), .ZN(new_n841));
  AND3_X1   g0641(.A1(new_n841), .A2(KEYINPUT104), .A3(new_n406), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT104), .B1(new_n841), .B2(new_n406), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n819), .A2(new_n820), .A3(new_n844), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n432), .A2(new_n820), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n844), .A2(new_n846), .B1(new_n421), .B2(new_n423), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n826), .B1(new_n847), .B2(new_n824), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n845), .A2(new_n848), .A3(KEYINPUT38), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n830), .A2(new_n835), .A3(new_n836), .A4(new_n849), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n845), .A2(KEYINPUT38), .A3(new_n848), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT38), .B1(new_n845), .B2(new_n848), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT39), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT106), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT106), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n850), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n617), .A2(new_n653), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n435), .A2(new_n650), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n788), .A2(new_n784), .ZN(new_n863));
  INV_X1    g0663(.A(new_n349), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(new_n653), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n353), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n851), .A2(new_n852), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n861), .A2(new_n862), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n622), .A2(new_n625), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n440), .B2(new_n688), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n872), .B(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n830), .A2(new_n835), .A3(new_n849), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n699), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n689), .A2(new_n702), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n867), .A2(new_n787), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT40), .ZN(new_n880));
  OR3_X1    g0680(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n880), .B1(new_n879), .B2(new_n869), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n440), .A2(new_n878), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n883), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(G330), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n875), .B(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n297), .B2(new_n646), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n599), .A2(new_n600), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT102), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n454), .B1(new_n890), .B2(KEYINPUT35), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n891), .B(new_n227), .C1(KEYINPUT35), .C2(new_n890), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT36), .ZN(new_n893));
  OAI21_X1  g0693(.A(G77), .B1(new_n206), .B2(new_n339), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n223), .A2(new_n894), .B1(G50), .B2(new_n339), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(G1), .A3(new_n645), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n888), .A2(new_n893), .A3(new_n896), .ZN(G367));
  OR3_X1    g0697(.A1(new_n633), .A2(new_n634), .A3(new_n653), .ZN(new_n898));
  OR3_X1    g0698(.A1(new_n898), .A2(KEYINPUT107), .A3(new_n627), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT107), .B1(new_n898), .B2(new_n627), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n898), .A2(new_n627), .A3(new_n635), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(KEYINPUT43), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT109), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n613), .A2(new_n665), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n610), .A2(new_n665), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n607), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n906), .B1(new_n909), .B2(new_n613), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n905), .B1(new_n662), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n662), .A2(new_n905), .A3(new_n910), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n904), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n902), .A2(KEYINPUT43), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT42), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT108), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n667), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n668), .A2(new_n910), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n511), .A2(new_n910), .A3(new_n663), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n906), .B1(new_n921), .B2(new_n918), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n920), .B(new_n922), .C1(KEYINPUT108), .C2(new_n917), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n912), .A2(new_n904), .A3(new_n913), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n915), .A2(new_n916), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n916), .ZN(new_n926));
  INV_X1    g0726(.A(new_n924), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n926), .B1(new_n927), .B2(new_n914), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n671), .B(KEYINPUT41), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n664), .B1(new_n655), .B2(new_n663), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(new_n660), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n932), .A2(new_n706), .A3(new_n688), .ZN(new_n933));
  INV_X1    g0733(.A(new_n910), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n668), .A2(new_n934), .B1(KEYINPUT110), .B2(KEYINPUT44), .ZN(new_n935));
  NOR2_X1   g0735(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT111), .Z(new_n937));
  XNOR2_X1  g0737(.A(new_n935), .B(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n662), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n668), .A2(new_n934), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT45), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n938), .A2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n662), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n933), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n930), .B1(new_n945), .B2(new_n707), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n925), .B(new_n928), .C1(new_n946), .C2(new_n772), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n368), .A2(new_n230), .ZN(new_n948));
  INV_X1    g0748(.A(new_n241), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n768), .B(new_n948), .C1(new_n755), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n725), .A2(G143), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n339), .B2(new_n727), .ZN(new_n952));
  INV_X1    g0752(.A(G137), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n718), .A2(new_n285), .B1(new_n711), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n734), .A2(new_n217), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n272), .B1(new_n717), .B2(new_n292), .ZN(new_n956));
  NOR4_X1   g0756(.A1(new_n952), .A2(new_n954), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n957), .B1(new_n206), .B2(new_n721), .C1(new_n379), .C2(new_n733), .ZN(new_n958));
  INV_X1    g0758(.A(new_n733), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(G294), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n721), .A2(new_n454), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n961), .A2(KEYINPUT46), .B1(new_n208), .B2(new_n727), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(G311), .B2(new_n725), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n391), .B1(new_n961), .B2(KEYINPUT46), .ZN(new_n964));
  INV_X1    g0764(.A(G317), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n717), .A2(new_n747), .B1(new_n711), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G97), .B2(new_n800), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n960), .A2(new_n963), .A3(new_n964), .A4(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n718), .A2(new_n744), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n958), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT47), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n950), .B1(new_n971), .B2(new_n752), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n972), .B(new_n773), .C1(new_n774), .C2(new_n902), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n947), .A2(new_n973), .ZN(G387));
  INV_X1    g0774(.A(KEYINPUT112), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n933), .B2(new_n677), .ZN(new_n976));
  INV_X1    g0776(.A(new_n932), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n707), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(KEYINPUT112), .A3(new_n671), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n976), .B(new_n979), .C1(new_n707), .C2(new_n977), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n772), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n755), .B1(new_n238), .B2(new_n253), .ZN(new_n982));
  INV_X1    g0782(.A(new_n672), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n982), .B1(new_n983), .B2(new_n759), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n339), .A2(new_n217), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n365), .A2(new_n285), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n672), .B1(new_n986), .B2(KEYINPUT50), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n987), .B(new_n253), .C1(KEYINPUT50), .C2(new_n986), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n984), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n670), .A2(new_n208), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n768), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n725), .A2(G322), .B1(new_n795), .B2(G317), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n747), .B2(new_n718), .C1(new_n733), .C2(new_n740), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT48), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n744), .B2(new_n727), .C1(new_n737), .C2(new_n721), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT49), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n742), .A2(G326), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n995), .A2(new_n996), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n391), .B1(G116), .B2(new_n800), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n718), .A2(new_n339), .B1(new_n711), .B2(new_n292), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n804), .A2(new_n367), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n522), .B2(new_n734), .C1(new_n726), .C2(new_n379), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1002), .B(new_n1004), .C1(G50), .C2(new_n795), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n721), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(G77), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1005), .B(new_n1007), .C1(new_n293), .C2(new_n733), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1001), .B1(new_n753), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n991), .B1(new_n1009), .B2(new_n752), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1010), .B(new_n773), .C1(new_n655), .C2(new_n774), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n980), .A2(new_n981), .A3(new_n1011), .ZN(G393));
  INV_X1    g0812(.A(new_n718), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n810), .B1(new_n365), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n339), .B2(new_n721), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n753), .B(new_n1015), .C1(G77), .C2(new_n804), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n742), .A2(G143), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n725), .A2(G150), .B1(new_n795), .B2(G159), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT51), .Z(new_n1019));
  NAND2_X1  g0819(.A1(new_n959), .A2(G50), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n272), .B1(new_n800), .B2(G107), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n744), .B2(new_n721), .C1(new_n739), .C2(new_n711), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT114), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n725), .A2(G317), .B1(new_n795), .B2(G311), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT52), .Z(new_n1026));
  AOI22_X1  g0826(.A1(new_n959), .A2(G303), .B1(G294), .B2(new_n1013), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n727), .A2(new_n454), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1021), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n752), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n755), .A2(new_n245), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n768), .B1(G97), .B2(new_n670), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n791), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT113), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1031), .B(new_n1035), .C1(new_n910), .C2(new_n774), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n944), .A2(new_n942), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1036), .B1(new_n1037), .B2(new_n771), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT115), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1037), .A2(new_n978), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT116), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n677), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1037), .A2(KEYINPUT116), .A3(new_n978), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1043), .A2(new_n945), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1040), .A2(new_n1045), .ZN(G390));
  AND3_X1   g0846(.A1(new_n850), .A2(new_n856), .A3(new_n853), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n856), .B1(new_n850), .B2(new_n853), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n764), .ZN(new_n1050));
  INV_X1    g0850(.A(G128), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n272), .B1(new_n727), .B2(new_n379), .C1(new_n726), .C2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G132), .B2(new_n795), .ZN(new_n1053));
  XOR2_X1   g0853(.A(KEYINPUT54), .B(G143), .Z(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1055), .A2(new_n718), .B1(new_n734), .B2(new_n285), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT53), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n721), .B2(new_n292), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1006), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1053), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(G125), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1061), .B1(new_n1062), .B2(new_n711), .C1(new_n953), .C2(new_n733), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n801), .B1(new_n454), .B2(new_n717), .C1(new_n737), .C2(new_n711), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G97), .B2(new_n1013), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n959), .A2(G107), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n804), .A2(G77), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n272), .B(new_n722), .C1(G283), .C2(new_n725), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n794), .B1(new_n1063), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n293), .B2(new_n814), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1050), .A2(new_n773), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(G330), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n785), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n867), .A2(new_n704), .A3(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n353), .B(new_n865), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n685), .A2(new_n653), .A3(new_n783), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(new_n784), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1079), .A2(new_n876), .A3(new_n860), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n868), .A2(new_n859), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1076), .B(new_n1080), .C1(new_n1049), .C2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n867), .A2(new_n878), .A3(new_n1075), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1077), .B1(new_n788), .B2(new_n784), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n855), .B(new_n857), .C1(new_n860), .C2(new_n1085), .ZN(new_n1086));
  OR3_X1    g0886(.A1(new_n1079), .A2(new_n860), .A3(new_n876), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n772), .B1(new_n1082), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(KEYINPUT118), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1076), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1085), .A2(new_n860), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1091), .B(new_n1087), .C1(new_n858), .C2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1080), .B1(new_n1049), .B2(new_n1081), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1093), .B1(new_n1094), .B2(new_n1084), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT118), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1095), .A2(new_n1096), .A3(new_n772), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1073), .B1(new_n1090), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n704), .A2(new_n1075), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n1077), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1100), .A2(KEYINPUT117), .A3(new_n1083), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT117), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1099), .A2(new_n1102), .A3(new_n1077), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n863), .A3(new_n1103), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1078), .A2(new_n784), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n878), .A2(new_n1075), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1105), .B(new_n1076), .C1(new_n867), .C2(new_n1106), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n688), .A2(new_n440), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n884), .A2(G330), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n626), .A3(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1095), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n1083), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n874), .A2(new_n1110), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1115), .A2(new_n1117), .A3(new_n1093), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1113), .A2(new_n1118), .A3(new_n671), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1098), .A2(new_n1119), .ZN(G378));
  NAND2_X1  g0920(.A1(new_n314), .A2(new_n317), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n304), .A2(new_n650), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1122), .B(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1124), .B(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n881), .A2(new_n882), .A3(G330), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n872), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n870), .B1(new_n860), .B2(new_n858), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1128), .B1(new_n1131), .B2(new_n862), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1127), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n872), .A2(new_n1129), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1131), .A2(new_n862), .A3(new_n1128), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n1126), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1133), .A2(new_n772), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n814), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n773), .B1(new_n1138), .B2(G50), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT120), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n726), .A2(new_n1062), .B1(new_n727), .B2(new_n292), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n1055), .A2(new_n721), .B1(new_n1051), .B2(new_n717), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n959), .C2(G132), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n953), .B2(new_n718), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT119), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1145), .A2(KEYINPUT59), .ZN(new_n1146));
  AOI211_X1 g0946(.A(G41), .B(new_n1146), .C1(G159), .C2(new_n800), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n742), .A2(G124), .ZN(new_n1148));
  AOI211_X1 g0948(.A(G33), .B(new_n1148), .C1(new_n1145), .C2(KEYINPUT59), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n252), .B1(new_n384), .B2(new_n268), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1147), .A2(new_n1149), .B1(new_n285), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n733), .A2(new_n522), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n717), .A2(new_n208), .B1(new_n711), .B2(new_n744), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n734), .A2(new_n206), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1155), .B(new_n753), .C1(new_n368), .C2(new_n718), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1007), .B1(new_n339), .B2(new_n727), .C1(new_n726), .C2(new_n454), .ZN(new_n1157));
  NOR4_X1   g0957(.A1(new_n1152), .A2(new_n1156), .A3(new_n1157), .A4(G41), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT58), .Z(new_n1159));
  AND2_X1   g0959(.A1(new_n1151), .A2(new_n1159), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1140), .B1(new_n794), .B2(new_n1160), .C1(new_n1126), .C2(new_n765), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1137), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1113), .A2(new_n874), .A3(new_n1110), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1163), .A2(new_n1133), .A3(KEYINPUT57), .A4(new_n1136), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n671), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1134), .A2(new_n1126), .A3(new_n1135), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1126), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT57), .B1(new_n1168), .B2(new_n1163), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1162), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT122), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(KEYINPUT122), .B(new_n1162), .C1(new_n1165), .C2(new_n1169), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(G375));
  NAND2_X1  g0974(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1175), .A2(new_n1117), .A3(new_n929), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n959), .A2(G116), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n272), .B(new_n955), .C1(G294), .C2(new_n725), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n717), .A2(new_n744), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n721), .A2(new_n522), .B1(new_n718), .B2(new_n208), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(G303), .C2(new_n742), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1177), .A2(new_n1003), .A3(new_n1178), .A4(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n959), .A2(new_n1054), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G137), .A2(new_n795), .B1(new_n1013), .B2(G150), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n753), .B1(G128), .B2(new_n742), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n727), .A2(new_n285), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1186), .B(new_n1154), .C1(G132), .C2(new_n725), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n721), .A2(new_n379), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1182), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n752), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(G68), .B2(new_n1138), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n791), .B(new_n1192), .C1(new_n1077), .C2(new_n764), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1116), .B2(new_n772), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1176), .A2(new_n1194), .ZN(G381));
  INV_X1    g0995(.A(KEYINPUT123), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n1095), .A2(new_n1096), .A3(new_n772), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1096), .B1(new_n1095), .B2(new_n772), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1072), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1113), .A2(new_n1118), .A3(new_n671), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1196), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1098), .A2(KEYINPUT123), .A3(new_n1119), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1040), .A2(new_n947), .A3(new_n1045), .A4(new_n973), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(G384), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1176), .A2(new_n1207), .A3(new_n1194), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(G393), .A2(G396), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1206), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  OR3_X1    g1011(.A1(G375), .A2(new_n1204), .A3(new_n1211), .ZN(G407));
  NAND2_X1  g1012(.A1(new_n1211), .A2(G343), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1213), .A2(new_n1172), .A3(new_n1173), .A4(new_n1203), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(G213), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT124), .Z(G409));
  NAND2_X1  g1016(.A1(G390), .A2(G387), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1205), .ZN(new_n1218));
  AND2_X1   g1018(.A1(G393), .A2(G396), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1219), .A2(new_n1210), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1217), .B(new_n1205), .C1(new_n1210), .C2(new_n1219), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n651), .A2(G213), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT125), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1163), .A2(new_n1133), .A3(new_n929), .A4(new_n1136), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(new_n1137), .A3(new_n1161), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1199), .A2(new_n1196), .A3(new_n1200), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT123), .B1(new_n1098), .B2(new_n1119), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1225), .B(new_n1227), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1230));
  OAI211_X1 g1030(.A(G378), .B(new_n1162), .C1(new_n1165), .C2(new_n1169), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1225), .B1(new_n1203), .B2(new_n1227), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1224), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n651), .A2(G213), .A3(G2897), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT126), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT60), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1175), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1108), .A2(new_n1111), .A3(KEYINPUT60), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1239), .A2(new_n671), .A3(new_n1117), .A4(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1194), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1237), .B1(new_n1242), .B2(new_n1207), .ZN(new_n1243));
  AOI211_X1 g1043(.A(KEYINPUT126), .B(G384), .C1(new_n1241), .C2(new_n1194), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1242), .A2(new_n1207), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1236), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .A4(new_n1235), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1234), .A2(new_n1251), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1253), .B(new_n1224), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT62), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(KEYINPUT62), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1223), .B1(new_n1255), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1254), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1227), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT125), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1250), .B1(new_n1263), .B2(new_n1224), .ZN(new_n1264));
  OAI21_X1  g1064(.A(KEYINPUT63), .B1(new_n1260), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT63), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1223), .B1(new_n1254), .B2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1265), .A2(new_n1257), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1259), .A2(new_n1268), .ZN(G405));
  INV_X1    g1069(.A(KEYINPUT127), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1221), .A2(new_n1270), .A3(new_n1222), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1270), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1204), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1231), .ZN(new_n1275));
  OR3_X1    g1075(.A1(new_n1274), .A2(new_n1253), .A3(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1253), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1273), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1273), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(G402));
endmodule


