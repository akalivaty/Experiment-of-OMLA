//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1170, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1216, new_n1217, new_n1218;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  OR3_X1    g0010(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT64), .ZN(new_n211));
  OAI21_X1  g0011(.A(KEYINPUT64), .B1(new_n209), .B2(new_n210), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT0), .Z(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G58), .A2(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n217), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G97), .B2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(G116), .B2(G270), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G77), .A2(G244), .ZN(new_n227));
  AOI22_X1  g0027(.A1(new_n226), .A2(new_n227), .B1(new_n212), .B2(new_n211), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT65), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n210), .ZN(new_n232));
  INV_X1    g0032(.A(G58), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(new_n201), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G50), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n216), .B(new_n230), .C1(new_n232), .C2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT66), .B(G250), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G257), .ZN(new_n243));
  XOR2_X1   g0043(.A(G264), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  NOR2_X1   g0046(.A1(new_n201), .A2(new_n202), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n203), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT67), .ZN(new_n250));
  XOR2_X1   g0050(.A(G50), .B(G58), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G87), .B(G97), .Z(new_n253));
  XNOR2_X1  g0053(.A(G107), .B(G116), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  XNOR2_X1  g0056(.A(KEYINPUT68), .B(G41), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n209), .B(G274), .C1(new_n257), .C2(G45), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G77), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G222), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(G1698), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT69), .ZN(new_n270));
  INV_X1    g0070(.A(G223), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n265), .B(new_n268), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  OAI211_X1 g0073(.A(G1), .B(G13), .C1(new_n260), .C2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n259), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G226), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G179), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(G20), .B1(new_n234), .B2(G50), .ZN(new_n284));
  INV_X1    g0084(.A(G150), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n260), .A2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n284), .B1(new_n285), .B2(new_n287), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n231), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n291), .A2(new_n293), .B1(new_n219), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n293), .B1(new_n209), .B2(G20), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n296), .B1(new_n219), .B2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n283), .B(new_n299), .C1(G169), .C2(new_n281), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT72), .ZN(new_n302));
  INV_X1    g0102(.A(G190), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n302), .B1(new_n280), .B2(new_n303), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n276), .A2(KEYINPUT72), .A3(G190), .A4(new_n279), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n299), .B(KEYINPUT9), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n280), .A2(G200), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n306), .A2(KEYINPUT71), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT71), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n304), .B2(new_n305), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT10), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n312), .A2(new_n313), .A3(new_n307), .A4(new_n308), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n301), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n271), .A2(new_n267), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n266), .B(new_n316), .C1(G226), .C2(new_n267), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G87), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n274), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n259), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n274), .A2(G232), .A3(new_n277), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n321), .B(KEYINPUT76), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n320), .A2(G179), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n320), .B2(new_n322), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT77), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT77), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n320), .A2(new_n322), .A3(G179), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n317), .A2(new_n318), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n275), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n322), .A2(new_n330), .A3(new_n258), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n327), .B(new_n328), .C1(new_n331), .C2(new_n324), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT7), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n266), .B2(G20), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n262), .A2(G33), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n337));
  OAI211_X1 g0137(.A(KEYINPUT7), .B(new_n210), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n201), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G159), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n287), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G58), .A2(G68), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n210), .B1(new_n234), .B2(new_n342), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n339), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT75), .B1(new_n344), .B2(KEYINPUT16), .ZN(new_n345));
  INV_X1    g0145(.A(new_n293), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n344), .B2(KEYINPUT16), .ZN(new_n347));
  INV_X1    g0147(.A(new_n341), .ZN(new_n348));
  INV_X1    g0148(.A(new_n343), .ZN(new_n349));
  NOR3_X1   g0149(.A1(new_n266), .A2(new_n334), .A3(G20), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT7), .B1(new_n264), .B2(new_n210), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n348), .B(new_n349), .C1(new_n352), .C2(new_n201), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT75), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT16), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n345), .A2(new_n347), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n290), .A2(new_n294), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n297), .B2(new_n290), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n333), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT18), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT18), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n333), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT78), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n331), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n331), .A2(G190), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n357), .A2(new_n368), .A3(new_n369), .A4(new_n359), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT17), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n370), .A2(new_n371), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n366), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n357), .A2(new_n359), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n375), .A2(KEYINPUT17), .A3(new_n368), .A4(new_n369), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n370), .A2(new_n371), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(KEYINPUT78), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n365), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n278), .A2(G244), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n266), .A2(G232), .A3(new_n267), .ZN(new_n381));
  INV_X1    g0181(.A(G238), .ZN(new_n382));
  OAI221_X1 g0182(.A(new_n381), .B1(new_n206), .B2(new_n266), .C1(new_n270), .C2(new_n382), .ZN(new_n383));
  AOI211_X1 g0183(.A(new_n259), .B(new_n380), .C1(new_n383), .C2(new_n275), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n282), .ZN(new_n385));
  XOR2_X1   g0185(.A(KEYINPUT15), .B(G87), .Z(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n288), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n286), .B(KEYINPUT70), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n387), .B1(new_n210), .B2(new_n202), .C1(new_n388), .C2(new_n290), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(new_n293), .B1(new_n202), .B2(new_n295), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n202), .B2(new_n298), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n385), .B(new_n391), .C1(G169), .C2(new_n384), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n315), .A2(new_n379), .A3(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n261), .A2(new_n263), .A3(G226), .A4(new_n267), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n261), .A2(new_n263), .A3(G232), .A4(G1698), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G97), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT73), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT73), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(G33), .A3(G97), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n394), .A2(new_n395), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n275), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n278), .A2(G238), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n258), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT13), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT74), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT13), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n402), .A2(new_n407), .A3(new_n258), .A4(new_n403), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n404), .A2(KEYINPUT74), .A3(KEYINPUT13), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT14), .B1(new_n411), .B2(new_n324), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT14), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n409), .A2(new_n413), .A3(G169), .A4(new_n410), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n405), .A2(G179), .A3(new_n408), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n289), .A2(new_n202), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n287), .A2(new_n219), .B1(new_n210), .B2(G68), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n293), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n419), .B(KEYINPUT11), .ZN(new_n420));
  OR3_X1    g0220(.A1(new_n294), .A2(KEYINPUT12), .A3(G68), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT12), .B1(new_n294), .B2(G68), .ZN(new_n422));
  AOI22_X1  g0222(.A1(G68), .A2(new_n297), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n416), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n424), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n405), .A2(G190), .A3(new_n408), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n426), .B(new_n427), .C1(new_n411), .C2(new_n367), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n391), .B1(new_n384), .B2(G190), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n367), .B2(new_n384), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n425), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n393), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n295), .A2(new_n205), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n346), .B(new_n294), .C1(G1), .C2(new_n260), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n433), .B1(new_n434), .B2(new_n205), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT81), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G97), .A2(G107), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(G97), .A2(G107), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n438), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n207), .A2(KEYINPUT81), .A3(new_n439), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n437), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OR2_X1    g0244(.A1(KEYINPUT80), .A2(G97), .ZN(new_n445));
  NAND2_X1  g0245(.A1(KEYINPUT80), .A2(G97), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n206), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT6), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT79), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT79), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT6), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(G20), .B1(new_n444), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT82), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n287), .A2(new_n202), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n455), .B1(new_n454), .B2(new_n457), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n352), .A2(new_n206), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n436), .B1(new_n461), .B2(new_n346), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT4), .ZN(new_n463));
  INV_X1    g0263(.A(G244), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n463), .B1(new_n264), .B2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .A4(new_n267), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n266), .A2(G250), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n267), .B1(new_n469), .B2(KEYINPUT4), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n275), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT84), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(G41), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n209), .A2(G45), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT5), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n475), .B1(new_n257), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n476), .A2(KEYINPUT83), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n476), .A2(KEYINPUT83), .ZN(new_n479));
  OAI211_X1 g0279(.A(KEYINPUT84), .B(new_n273), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n474), .A2(new_n477), .A3(G274), .A4(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n474), .A2(new_n477), .A3(new_n480), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(G257), .A3(new_n274), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n471), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n324), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n471), .A2(new_n483), .A3(new_n282), .A4(new_n481), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n462), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n484), .A2(G200), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n303), .B2(new_n484), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n488), .B1(new_n462), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n261), .A2(new_n263), .A3(G244), .A4(G1698), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT85), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n266), .A2(KEYINPUT85), .A3(G244), .A4(G1698), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n266), .A2(G238), .A3(new_n267), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G116), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n494), .A2(new_n495), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n275), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n475), .A2(G274), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n475), .A2(new_n224), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(new_n274), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n303), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n502), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n498), .B2(new_n275), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(G200), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n434), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G87), .ZN(new_n508));
  INV_X1    g0308(.A(new_n386), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n295), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n397), .A2(new_n399), .A3(KEYINPUT19), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n210), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n445), .A2(new_n446), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(new_n223), .A3(new_n206), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n266), .A2(new_n210), .A3(G68), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT19), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n513), .B2(new_n289), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT87), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n515), .A2(KEYINPUT87), .A3(new_n516), .A4(new_n518), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n293), .A3(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n506), .A2(new_n508), .A3(new_n510), .A4(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n266), .A2(new_n210), .A3(G87), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT22), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n266), .A2(KEYINPUT22), .A3(new_n210), .A4(G87), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n288), .A2(G116), .ZN(new_n530));
  NAND2_X1  g0330(.A1(KEYINPUT93), .A2(KEYINPUT23), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(G20), .A3(new_n206), .ZN(new_n532));
  NOR2_X1   g0332(.A1(KEYINPUT93), .A2(KEYINPUT23), .ZN(new_n533));
  XNOR2_X1  g0333(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n529), .A2(KEYINPUT24), .A3(new_n530), .A4(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n527), .A2(new_n534), .A3(new_n530), .A4(new_n528), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT24), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n535), .A2(new_n293), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT25), .B1(new_n294), .B2(G107), .ZN(new_n540));
  OR3_X1    g0340(.A1(new_n294), .A2(KEYINPUT25), .A3(G107), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n540), .B(new_n541), .C1(new_n434), .C2(new_n206), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT94), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n482), .A2(G264), .A3(new_n274), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n266), .B1(G250), .B2(G1698), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n267), .A2(G257), .ZN(new_n547));
  INV_X1    g0347(.A(G294), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n546), .A2(new_n547), .B1(new_n260), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n275), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n545), .A2(new_n550), .A3(new_n481), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G200), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n545), .A2(new_n550), .A3(G190), .A4(new_n481), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n539), .A2(new_n544), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n524), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n539), .A2(new_n544), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n551), .A2(new_n324), .ZN(new_n557));
  OR2_X1    g0357(.A1(new_n551), .A2(G179), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n491), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(G116), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n346), .B1(G20), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT91), .ZN(new_n563));
  OR2_X1    g0363(.A1(new_n563), .A2(KEYINPUT20), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n445), .A2(new_n260), .A3(new_n446), .ZN(new_n565));
  AOI21_X1  g0365(.A(G20), .B1(G33), .B2(G283), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(KEYINPUT90), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT90), .B1(new_n565), .B2(new_n566), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n562), .B(new_n564), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n563), .A2(KEYINPUT20), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n569), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n567), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n574), .A2(new_n563), .A3(KEYINPUT20), .A4(new_n562), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT89), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n294), .B2(G116), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n295), .A2(KEYINPUT89), .A3(new_n561), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n507), .A2(G116), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n324), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(G303), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n274), .B1(new_n264), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n267), .A2(G257), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G264), .A2(G1698), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n266), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n482), .A2(G270), .A3(new_n274), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT88), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n588), .A2(new_n589), .A3(new_n481), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n588), .B2(new_n481), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n581), .A2(new_n592), .A3(KEYINPUT21), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT92), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n581), .A2(new_n592), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n581), .A2(new_n592), .A3(KEYINPUT92), .A4(KEYINPUT21), .ZN(new_n599));
  INV_X1    g0399(.A(new_n592), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n576), .A2(new_n580), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(G179), .A3(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n595), .A2(new_n598), .A3(new_n599), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(G190), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n592), .A2(G200), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n604), .A2(new_n580), .A3(new_n605), .A4(new_n576), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n507), .A2(new_n386), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n523), .A2(new_n510), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n505), .A2(G179), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n324), .B2(new_n505), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT86), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n610), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n432), .A2(new_n560), .A3(new_n608), .A4(new_n616), .ZN(G372));
  INV_X1    g0417(.A(new_n392), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n428), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n619), .A2(new_n425), .B1(new_n374), .B2(new_n378), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n328), .B1(new_n331), .B2(new_n324), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n360), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n363), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n360), .A2(KEYINPUT18), .A3(new_n621), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n310), .B2(new_n314), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n628), .A2(new_n301), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n610), .A2(new_n612), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n462), .A2(new_n630), .A3(new_n524), .A4(new_n487), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT95), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n485), .A2(new_n486), .ZN(new_n636));
  INV_X1    g0436(.A(new_n459), .ZN(new_n637));
  INV_X1    g0437(.A(new_n460), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n293), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n636), .B1(new_n641), .B2(new_n436), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n616), .A2(new_n642), .A3(KEYINPUT26), .A4(new_n524), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n631), .A2(KEYINPUT95), .A3(new_n632), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n635), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n462), .A2(new_n490), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(new_n642), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n630), .A2(new_n524), .A3(new_n554), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n647), .B(new_n648), .C1(new_n603), .C2(new_n559), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n645), .A2(new_n649), .A3(new_n630), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n432), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n629), .A2(new_n651), .ZN(G369));
  INV_X1    g0452(.A(G13), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(G20), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT27), .B1(new_n655), .B2(G1), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n654), .A2(new_n657), .A3(new_n209), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT96), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n601), .A2(new_n665), .ZN(new_n666));
  MUX2_X1   g0466(.A(new_n603), .B(new_n608), .S(new_n666), .Z(new_n667));
  AND2_X1   g0467(.A1(new_n667), .A2(G330), .ZN(new_n668));
  INV_X1    g0468(.A(new_n554), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n556), .B2(new_n665), .ZN(new_n670));
  MUX2_X1   g0470(.A(new_n670), .B(new_n665), .S(new_n559), .Z(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n665), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n559), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n603), .A2(new_n673), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(new_n674), .A3(new_n676), .ZN(G399));
  INV_X1    g0477(.A(new_n214), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n257), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n514), .A2(G116), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n679), .A2(new_n209), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n236), .B2(new_n679), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT28), .Z(new_n683));
  NAND2_X1  g0483(.A1(new_n650), .A2(new_n673), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT29), .ZN(new_n685));
  INV_X1    g0485(.A(new_n611), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n545), .A2(new_n550), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n484), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n600), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n484), .A2(new_n551), .ZN(new_n692));
  INV_X1    g0492(.A(new_n505), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n592), .A2(new_n692), .A3(new_n282), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  OAI22_X1  g0495(.A1(new_n695), .A2(KEYINPUT97), .B1(new_n690), .B2(new_n689), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n695), .A2(KEYINPUT97), .ZN(new_n697));
  OAI211_X1 g0497(.A(KEYINPUT31), .B(new_n665), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n689), .A2(new_n690), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n665), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n608), .A2(new_n560), .A3(new_n616), .A4(new_n673), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n698), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n646), .A2(new_n642), .A3(new_n555), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n603), .B2(new_n559), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n616), .A2(new_n632), .A3(new_n524), .A4(new_n642), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n642), .A2(new_n524), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n709), .A2(KEYINPUT26), .B1(new_n610), .B2(new_n612), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n673), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n685), .A2(new_n705), .A3(new_n713), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT98), .Z(new_n715));
  OAI21_X1  g0515(.A(new_n683), .B1(new_n715), .B2(G1), .ZN(G364));
  AOI21_X1  g0516(.A(new_n209), .B1(new_n654), .B2(G45), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n679), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n668), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(G330), .B2(new_n667), .ZN(new_n721));
  INV_X1    g0521(.A(new_n719), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n214), .A2(G355), .A3(new_n266), .ZN(new_n723));
  INV_X1    g0523(.A(G45), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n252), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n678), .A2(new_n266), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(G45), .B2(new_n235), .ZN(new_n727));
  OAI221_X1 g0527(.A(new_n723), .B1(G116), .B2(new_n214), .C1(new_n725), .C2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n231), .B1(G20), .B2(new_n324), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n728), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n210), .A2(new_n303), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n367), .A2(G179), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n582), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G179), .A2(G200), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n210), .B1(new_n739), .B2(G190), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n264), .B1(new_n740), .B2(new_n548), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n282), .A2(new_n367), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n210), .A2(G190), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT100), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n744), .A2(KEYINPUT100), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  XNOR2_X1  g0549(.A(KEYINPUT33), .B(G317), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n738), .B(new_n741), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n282), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n735), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G322), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n752), .A2(new_n743), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(KEYINPUT99), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n756), .A2(KEYINPUT99), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G311), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n735), .A2(new_n742), .ZN(new_n763));
  INV_X1    g0563(.A(G326), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n743), .A2(new_n739), .ZN(new_n765));
  INV_X1    g0565(.A(G329), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n763), .A2(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n743), .A2(new_n736), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n767), .B1(G283), .B2(new_n769), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n751), .A2(new_n755), .A3(new_n762), .A4(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n761), .A2(G77), .B1(G58), .B2(new_n754), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n763), .A2(new_n219), .B1(new_n737), .B2(new_n223), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n768), .A2(new_n206), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n740), .A2(new_n205), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n773), .A2(new_n774), .A3(new_n775), .A4(new_n264), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n772), .B(new_n776), .C1(new_n201), .C2(new_n748), .ZN(new_n777));
  INV_X1    g0577(.A(new_n765), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G159), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT32), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n771), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT101), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n722), .B(new_n734), .C1(new_n782), .C2(new_n732), .ZN(new_n783));
  INV_X1    g0583(.A(new_n731), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n783), .B1(new_n667), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n721), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(G396));
  NOR2_X1   g0587(.A1(new_n392), .A2(new_n665), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n391), .A2(new_n665), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n430), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n788), .B1(new_n392), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n684), .B(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(new_n705), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n722), .ZN(new_n794));
  INV_X1    g0594(.A(G283), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n264), .B1(new_n760), .B2(new_n561), .C1(new_n795), .C2(new_n748), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n775), .B1(G294), .B2(new_n754), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT102), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n582), .B2(new_n763), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n797), .A2(new_n798), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n768), .A2(new_n223), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n796), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n206), .B2(new_n737), .C1(new_n804), .C2(new_n765), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n737), .A2(new_n219), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n749), .A2(G150), .B1(G143), .B2(new_n754), .ZN(new_n807));
  INV_X1    g0607(.A(G137), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n807), .B1(new_n808), .B2(new_n763), .C1(new_n340), .C2(new_n760), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT34), .Z(new_n810));
  AOI211_X1 g0610(.A(new_n806), .B(new_n810), .C1(G132), .C2(new_n778), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n811), .B1(new_n233), .B2(new_n740), .C1(new_n201), .C2(new_n768), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n805), .B1(new_n812), .B2(new_n264), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n722), .B1(new_n813), .B2(new_n732), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n732), .A2(new_n729), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n814), .B1(G77), .B2(new_n815), .C1(new_n730), .C2(new_n791), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n794), .A2(new_n816), .ZN(G384));
  NAND3_X1  g0617(.A1(new_n650), .A2(new_n673), .A3(new_n791), .ZN(new_n818));
  INV_X1    g0618(.A(new_n788), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n665), .A2(new_n424), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n425), .A2(new_n428), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n416), .A2(new_n424), .A3(new_n665), .ZN(new_n823));
  AND3_X1   g0623(.A1(new_n822), .A2(KEYINPUT103), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(KEYINPUT103), .B1(new_n822), .B2(new_n823), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n820), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(KEYINPUT104), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n347), .B1(KEYINPUT16), .B2(new_n344), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n359), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n621), .ZN(new_n832));
  INV_X1    g0632(.A(new_n663), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n832), .A2(new_n834), .A3(new_n370), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT37), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n663), .B(KEYINPUT105), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n360), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n361), .A2(new_n838), .A3(new_n370), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n836), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n379), .B2(new_n834), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT38), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(KEYINPUT38), .B(new_n842), .C1(new_n379), .C2(new_n834), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT104), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n820), .A2(new_n848), .A3(new_n827), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n829), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n845), .A2(KEYINPUT39), .A3(new_n846), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n622), .A2(new_n838), .A3(new_n370), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n839), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n853), .A2(new_n841), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n372), .A2(new_n373), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n838), .B1(new_n855), .B2(new_n625), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n844), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n846), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT39), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n851), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n425), .A2(new_n665), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n625), .A2(new_n837), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n850), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n713), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n684), .A2(KEYINPUT29), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n432), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n868), .A2(new_n629), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n865), .B(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT107), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n700), .A2(new_n871), .A3(new_n701), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n665), .B1(KEYINPUT107), .B2(KEYINPUT31), .C1(new_n695), .C2(new_n699), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n703), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n791), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n875), .A2(new_n826), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(new_n847), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n827), .A2(new_n791), .A3(new_n874), .ZN(new_n879));
  INV_X1    g0679(.A(new_n858), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT40), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(new_n432), .A3(new_n874), .ZN(new_n883));
  INV_X1    g0683(.A(G330), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n878), .B2(new_n881), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n432), .A2(G330), .A3(new_n874), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n883), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n870), .B(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n209), .B2(new_n654), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n444), .A2(new_n453), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n561), .B1(new_n891), .B2(KEYINPUT35), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n892), .B(new_n232), .C1(KEYINPUT35), .C2(new_n891), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT36), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n342), .A2(G77), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n235), .A2(new_n895), .B1(G50), .B2(new_n201), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(G1), .A3(new_n653), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n890), .A2(new_n894), .A3(new_n897), .ZN(G367));
  AOI21_X1  g0698(.A(new_n264), .B1(new_n769), .B2(G77), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT114), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n760), .B2(new_n219), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n899), .A2(KEYINPUT114), .B1(new_n808), .B2(new_n765), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n740), .A2(new_n201), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n340), .B2(new_n748), .ZN(new_n905));
  INV_X1    g0705(.A(new_n763), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n901), .B(new_n905), .C1(G143), .C2(new_n906), .ZN(new_n907));
  OAI221_X1 g0707(.A(new_n907), .B1(new_n233), .B2(new_n737), .C1(new_n285), .C2(new_n753), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n763), .A2(new_n804), .B1(new_n753), .B2(new_n582), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT112), .Z(new_n910));
  NOR2_X1   g0710(.A1(new_n768), .A2(new_n513), .ZN(new_n911));
  INV_X1    g0711(.A(new_n737), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(KEYINPUT46), .A3(G116), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n264), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n740), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(G107), .ZN(new_n917));
  INV_X1    g0717(.A(G317), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n760), .A2(new_n795), .B1(new_n918), .B2(new_n765), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(G294), .B2(new_n749), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n915), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT46), .B1(new_n912), .B2(G116), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT113), .Z(new_n923));
  OAI21_X1  g0723(.A(new_n908), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT47), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n732), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n523), .A2(new_n510), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n434), .A2(new_n223), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n665), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n524), .A3(new_n630), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n630), .B2(new_n929), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n931), .A2(new_n784), .ZN(new_n932));
  INV_X1    g0732(.A(new_n726), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n733), .B1(new_n214), .B2(new_n509), .C1(new_n933), .C2(new_n245), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n926), .A2(new_n719), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT111), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n679), .B(KEYINPUT41), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n676), .A2(new_n674), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n673), .B1(new_n641), .B2(new_n436), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n491), .A2(new_n939), .B1(new_n488), .B2(new_n673), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT44), .Z(new_n943));
  NOR2_X1   g0743(.A1(new_n938), .A2(new_n941), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT45), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n943), .A2(new_n672), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n672), .B1(new_n943), .B2(new_n945), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n672), .ZN(new_n950));
  INV_X1    g0750(.A(new_n668), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT110), .B1(new_n671), .B2(new_n675), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(new_n676), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n950), .A2(KEYINPUT110), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n715), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n949), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n715), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n936), .B(new_n937), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n957), .B1(new_n948), .B2(new_n954), .ZN(new_n959));
  INV_X1    g0759(.A(new_n937), .ZN(new_n960));
  OAI21_X1  g0760(.A(KEYINPUT111), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n718), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n931), .B(KEYINPUT43), .Z(new_n963));
  NOR3_X1   g0763(.A1(new_n676), .A2(new_n491), .A3(new_n939), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT42), .Z(new_n965));
  XOR2_X1   g0765(.A(new_n940), .B(KEYINPUT108), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n559), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n665), .B1(new_n967), .B2(new_n488), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n963), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(KEYINPUT109), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(KEYINPUT109), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n965), .A2(new_n968), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n970), .B(new_n971), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n966), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n672), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n974), .B(new_n976), .Z(new_n977));
  OAI21_X1  g0777(.A(new_n935), .B1(new_n962), .B2(new_n977), .ZN(G387));
  NAND2_X1  g0778(.A1(new_n954), .A2(new_n718), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n748), .A2(new_n290), .B1(new_n509), .B2(new_n740), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n760), .A2(new_n201), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n266), .B1(new_n768), .B2(new_n205), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n763), .A2(new_n340), .B1(new_n765), .B2(new_n285), .ZN(new_n983));
  NOR4_X1   g0783(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n984), .B1(new_n219), .B2(new_n753), .C1(new_n202), .C2(new_n737), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n761), .A2(G303), .B1(G322), .B2(new_n906), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n804), .B2(new_n748), .C1(new_n918), .C2(new_n753), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT48), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n795), .B2(new_n740), .C1(new_n548), .C2(new_n737), .ZN(new_n989));
  XNOR2_X1  g0789(.A(KEYINPUT116), .B(KEYINPUT49), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n264), .B1(new_n765), .B2(new_n764), .C1(new_n561), .C2(new_n768), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n985), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n732), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n680), .A2(new_n214), .A3(new_n266), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n680), .B(KEYINPUT115), .ZN(new_n996));
  INV_X1    g0796(.A(new_n290), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n219), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT50), .ZN(new_n999));
  NOR4_X1   g0799(.A1(new_n996), .A2(G45), .A3(new_n247), .A4(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n726), .B1(new_n241), .B2(new_n724), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n995), .B1(G107), .B2(new_n214), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n722), .B1(new_n1002), .B2(new_n733), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n994), .B(new_n1003), .C1(new_n671), .C2(new_n784), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n715), .A2(new_n954), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n679), .B1(new_n715), .B2(new_n954), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n979), .B(new_n1004), .C1(new_n1005), .C2(new_n1006), .ZN(G393));
  AOI22_X1  g0807(.A1(new_n749), .A2(G50), .B1(G77), .B2(new_n916), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n290), .B2(new_n760), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT117), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n763), .A2(new_n285), .B1(new_n753), .B2(new_n340), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT51), .Z(new_n1012));
  AOI211_X1 g0812(.A(new_n264), .B(new_n802), .C1(G143), .C2(new_n778), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n201), .B2(new_n737), .ZN(new_n1014));
  NOR3_X1   g0814(.A1(new_n1010), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G317), .A2(new_n906), .B1(new_n754), .B2(G311), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n264), .B1(new_n1016), .B2(KEYINPUT52), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1017), .A2(new_n774), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n761), .A2(G294), .B1(G322), .B2(new_n778), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n749), .A2(G303), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1016), .A2(KEYINPUT52), .B1(G116), .B2(new_n916), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G283), .B2(new_n912), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n732), .B1(new_n1015), .B2(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n733), .B1(new_n214), .B2(new_n513), .C1(new_n933), .C2(new_n255), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1024), .A2(new_n719), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n975), .B2(new_n731), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n948), .B2(new_n718), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n679), .B1(new_n1005), .B2(new_n948), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n1029), .B2(new_n956), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT118), .ZN(G390));
  INV_X1    g0831(.A(KEYINPUT124), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n768), .A2(new_n201), .B1(new_n765), .B2(new_n548), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n760), .A2(new_n513), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G87), .B2(new_n912), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n266), .B1(new_n1033), .B2(new_n1032), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n749), .A2(G107), .B1(G77), .B2(new_n916), .ZN(new_n1037));
  AND3_X1   g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n561), .B2(new_n753), .C1(new_n795), .C2(new_n763), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n749), .A2(G137), .B1(G159), .B2(new_n916), .ZN(new_n1040));
  XOR2_X1   g0840(.A(KEYINPUT54), .B(G143), .Z(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1040), .B1(new_n760), .B2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT123), .Z(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G128), .B2(new_n906), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n737), .A2(new_n285), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT53), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n264), .B1(new_n754), .B2(G132), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n769), .A2(G50), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(G125), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n765), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1039), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n722), .B1(new_n1053), .B2(new_n732), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n997), .B2(new_n815), .C1(new_n861), .C2(new_n730), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n862), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n828), .A2(new_n1056), .B1(new_n851), .B2(new_n860), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n790), .A2(new_n392), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n711), .A2(new_n673), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n819), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n827), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n862), .B(KEYINPUT119), .Z(new_n1062));
  AND3_X1   g0862(.A1(new_n1061), .A2(new_n858), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(KEYINPUT120), .B1(new_n1057), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1061), .A2(new_n858), .A3(new_n1062), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT120), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n862), .B1(new_n820), .B2(new_n827), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1065), .B(new_n1066), .C1(new_n861), .C2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n879), .A2(new_n884), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1064), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT121), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n827), .A2(new_n704), .A3(G330), .A4(new_n791), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1073), .B(new_n1065), .C1(new_n861), .C2(new_n1067), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1064), .A2(new_n1068), .A3(KEYINPUT121), .A4(new_n1069), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1055), .B1(new_n1076), .B2(new_n717), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n826), .B1(new_n875), .B2(new_n884), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1078), .A2(new_n819), .A3(new_n1073), .A4(new_n1059), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n704), .A2(G330), .A3(new_n791), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n876), .A2(G330), .B1(new_n1080), .B2(new_n826), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n820), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n868), .A2(new_n629), .A3(new_n886), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT122), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n868), .A2(new_n629), .A3(KEYINPUT122), .A4(new_n886), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1083), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .A4(new_n1088), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1089), .A2(new_n679), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1088), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1076), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1077), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(G378));
  NAND2_X1  g0894(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1089), .A2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n315), .B(KEYINPUT55), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n833), .A2(new_n299), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1098), .B(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(KEYINPUT125), .B(KEYINPUT56), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n865), .A2(new_n885), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n865), .A2(new_n885), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n865), .A2(new_n885), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1104), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n1110), .A3(new_n1105), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1097), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT57), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1097), .A2(new_n1112), .A3(KEYINPUT57), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n679), .A3(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n768), .A2(new_n233), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G107), .A2(new_n754), .B1(new_n778), .B2(G283), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1119), .B1(new_n202), .B2(new_n737), .C1(new_n561), .C2(new_n763), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1118), .B(new_n1120), .C1(new_n386), .C2(new_n761), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n903), .A2(new_n266), .A3(new_n257), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(new_n205), .C2(new_n748), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT58), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n219), .B1(G33), .B2(G41), .C1(new_n266), .C2(new_n257), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1042), .A2(new_n737), .ZN(new_n1126));
  INV_X1    g0926(.A(G128), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n763), .A2(new_n1051), .B1(new_n753), .B2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1126), .B(new_n1128), .C1(new_n749), .C2(G132), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n808), .B2(new_n760), .C1(new_n285), .C2(new_n740), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT59), .ZN(new_n1131));
  AOI211_X1 g0931(.A(G33), .B(G41), .C1(new_n778), .C2(G124), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n340), .B2(new_n768), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1124), .B(new_n1125), .C1(new_n1131), .C2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n722), .B1(new_n1134), .B2(new_n732), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1135), .B1(G50), .B2(new_n815), .C1(new_n1104), .C2(new_n730), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT126), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n718), .B2(new_n1112), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1117), .A2(new_n1138), .ZN(G375));
  NAND2_X1  g0939(.A1(new_n826), .A2(new_n729), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n719), .B1(G68), .B2(new_n815), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n749), .A2(G116), .B1(G303), .B2(new_n778), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(G283), .A2(new_n754), .B1(new_n769), .B2(G77), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1142), .B(new_n1143), .C1(new_n205), .C2(new_n737), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G107), .B2(new_n761), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n266), .B1(new_n916), .B2(new_n386), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1145), .B(new_n1146), .C1(new_n548), .C2(new_n763), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT127), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n761), .A2(G150), .B1(G137), .B2(new_n754), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n264), .B1(new_n778), .B2(G128), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(new_n219), .C2(new_n740), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G159), .B2(new_n912), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1118), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n906), .A2(G132), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n749), .A2(new_n1041), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1148), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1141), .B1(new_n1157), .B2(new_n732), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1083), .A2(new_n718), .B1(new_n1140), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1083), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1095), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n937), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1159), .B1(new_n1162), .B2(new_n1088), .ZN(G381));
  OR2_X1    g0963(.A1(G387), .A2(G390), .ZN(new_n1164));
  OR2_X1    g0964(.A1(G393), .A2(G396), .ZN(new_n1165));
  NOR4_X1   g0965(.A1(new_n1164), .A2(G384), .A3(G381), .A4(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1117), .A2(new_n1093), .A3(new_n1138), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(G407));
  OAI21_X1  g0969(.A(new_n1168), .B1(new_n1166), .B2(new_n664), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(G213), .ZN(G409));
  XNOR2_X1  g0971(.A(G393), .B(new_n786), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(G387), .A2(G390), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(G387), .A2(G390), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1173), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1164), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1093), .B1(new_n1117), .B2(new_n1138), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n960), .B1(new_n1089), .B2(new_n1096), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1112), .B1(new_n1182), .B2(new_n718), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1093), .A2(new_n1183), .A3(new_n1136), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT60), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1091), .B(new_n679), .C1(new_n1186), .C2(new_n1161), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT60), .B1(new_n1095), .B2(new_n1160), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1159), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1189), .A2(new_n794), .A3(new_n816), .ZN(new_n1190));
  OAI211_X1 g0990(.A(G384), .B(new_n1159), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n664), .A2(G213), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NOR4_X1   g0994(.A1(new_n1181), .A2(new_n1185), .A3(new_n1192), .A4(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT62), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1181), .A2(new_n1194), .A3(new_n1185), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1194), .A2(G2897), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1192), .B(new_n1198), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n1195), .A2(new_n1196), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT61), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(G375), .A2(G378), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1192), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1202), .A2(new_n1203), .A3(new_n1193), .A4(new_n1184), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1201), .B1(new_n1204), .B2(KEYINPUT62), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1180), .B1(new_n1200), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT61), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1195), .A2(KEYINPUT63), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT63), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1202), .A2(new_n1193), .A3(new_n1184), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1194), .A2(G2897), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1192), .B(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1209), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1207), .B(new_n1208), .C1(new_n1213), .C2(new_n1195), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1206), .A2(new_n1214), .ZN(G405));
  OAI21_X1  g1015(.A(new_n1203), .B1(new_n1168), .B2(new_n1181), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1202), .A2(new_n1167), .A3(new_n1192), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(new_n1179), .ZN(G402));
endmodule


