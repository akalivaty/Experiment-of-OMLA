//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1239, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT64), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g0017(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n209), .ZN(new_n221));
  INV_X1    g0021(.A(new_n201), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G50), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT65), .Z(new_n224));
  AOI21_X1  g0024(.A(new_n214), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G226), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI22_X1  g0028(.A1(new_n202), .A2(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(G116), .B2(G270), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT66), .B(G68), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT67), .B(G238), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n230), .B(new_n231), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  AOI22_X1  g0034(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT68), .Z(new_n236));
  OAI21_X1  g0036(.A(new_n211), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g0037(.A(new_n225), .B1(KEYINPUT1), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g0038(.A(new_n238), .B1(KEYINPUT1), .B2(new_n237), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT69), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G264), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G58), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1698), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G222), .ZN(new_n261));
  INV_X1    g0061(.A(G77), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n258), .A2(new_n259), .ZN(new_n263));
  INV_X1    g0063(.A(G223), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(G1698), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n261), .B1(new_n262), .B2(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  INV_X1    g0067(.A(new_n218), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT70), .A2(G41), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT70), .A2(G41), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n274), .A2(new_n275), .A3(G45), .ZN(new_n276));
  AND2_X1   g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n208), .B(G274), .C1(new_n277), .C2(new_n215), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n267), .A2(G1), .A3(G13), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n226), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n272), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G200), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n272), .A2(G190), .A3(new_n284), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(KEYINPUT74), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n217), .A2(new_n289), .A3(new_n218), .A4(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n208), .A2(G20), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(G50), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n289), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n202), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT8), .B(G58), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n209), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(G150), .ZN(new_n299));
  NOR2_X1   g0099(.A1(G20), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n297), .A2(new_n298), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(G20), .B2(new_n203), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n217), .A2(new_n218), .A3(new_n290), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n294), .B(new_n296), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT9), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n305), .B(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT10), .B1(new_n288), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n305), .B(KEYINPUT9), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n287), .A2(KEYINPUT74), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT10), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .A4(new_n286), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n285), .A2(new_n314), .ZN(new_n315));
  XOR2_X1   g0115(.A(KEYINPUT71), .B(G179), .Z(new_n316));
  OAI211_X1 g0116(.A(new_n315), .B(new_n305), .C1(new_n316), .C2(new_n285), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  XOR2_X1   g0119(.A(KEYINPUT8), .B(G58), .Z(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n293), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n321), .A2(new_n291), .B1(new_n289), .B2(new_n320), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT79), .ZN(new_n323));
  INV_X1    g0123(.A(G58), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n222), .B1(new_n232), .B2(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n325), .A2(G20), .B1(G159), .B2(new_n300), .ZN(new_n326));
  AND2_X1   g0126(.A1(KEYINPUT3), .A2(G33), .ZN(new_n327));
  NOR2_X1   g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT7), .B1(new_n329), .B2(new_n209), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n259), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(G68), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n326), .A2(new_n333), .A3(KEYINPUT16), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n217), .A2(new_n218), .A3(new_n290), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n258), .A2(new_n209), .A3(new_n259), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT78), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(new_n340), .A3(new_n331), .ZN(new_n341));
  INV_X1    g0141(.A(G68), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT66), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT66), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G68), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n332), .A2(KEYINPUT78), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n341), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT16), .B1(new_n348), .B2(new_n326), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n323), .B1(new_n336), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n226), .A2(G1698), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n351), .B1(G223), .B2(G1698), .C1(new_n327), .C2(new_n328), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G33), .A2(G87), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT80), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n353), .B(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n270), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G232), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n276), .A2(new_n278), .B1(new_n282), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n314), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n316), .ZN(new_n362));
  NOR3_X1   g0162(.A1(new_n356), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n350), .A2(new_n365), .A3(KEYINPUT18), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT18), .B1(new_n350), .B2(new_n365), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n357), .A2(new_n360), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n356), .B2(new_n359), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n373), .B(new_n323), .C1(new_n336), .C2(new_n349), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT17), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n374), .B(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n368), .A2(new_n376), .ZN(new_n377));
  XOR2_X1   g0177(.A(KEYINPUT15), .B(G87), .Z(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n298), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n297), .A2(new_n301), .B1(new_n209), .B2(new_n262), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n335), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n292), .A2(G77), .A3(new_n293), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n295), .A2(new_n262), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT72), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G244), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n276), .A2(new_n278), .B1(new_n282), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n260), .A2(G232), .ZN(new_n389));
  INV_X1    g0189(.A(G107), .ZN(new_n390));
  OAI221_X1 g0190(.A(new_n389), .B1(new_n390), .B2(new_n263), .C1(new_n265), .C2(new_n233), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n388), .B1(new_n391), .B2(new_n271), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n386), .B1(new_n393), .B2(G200), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n369), .B2(new_n393), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n314), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n392), .A2(new_n362), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n397), .A3(new_n386), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n399), .A2(KEYINPUT73), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(KEYINPUT73), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n319), .A2(new_n377), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G97), .ZN(new_n404));
  INV_X1    g0204(.A(G1698), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n226), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n358), .A2(G1698), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n406), .B(new_n407), .C1(new_n327), .C2(new_n328), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n270), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G238), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n276), .A2(new_n278), .B1(new_n282), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT75), .B(KEYINPUT13), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n409), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT13), .B1(new_n409), .B2(new_n411), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT76), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g0217(.A(KEYINPUT76), .B(KEYINPUT13), .C1(new_n409), .C2(new_n411), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n414), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G179), .ZN(new_n420));
  INV_X1    g0220(.A(new_n411), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n408), .A2(new_n404), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n271), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n423), .A3(new_n412), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n413), .B1(new_n409), .B2(new_n411), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT14), .B1(new_n426), .B2(G169), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT14), .ZN(new_n428));
  AOI211_X1 g0228(.A(new_n428), .B(new_n314), .C1(new_n424), .C2(new_n425), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n420), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n232), .A2(G20), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n257), .A2(G20), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n432), .A2(G77), .B1(new_n300), .B2(G50), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n335), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT11), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT12), .B1(new_n295), .B2(new_n342), .ZN(new_n438));
  INV_X1    g0238(.A(new_n431), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n208), .A2(KEYINPUT12), .A3(G13), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n434), .A2(KEYINPUT11), .A3(new_n335), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n292), .A2(G68), .A3(new_n293), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n437), .A2(new_n441), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n430), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n419), .A2(G190), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(G200), .B2(new_n426), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT77), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT81), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n403), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT81), .B1(new_n402), .B2(new_n450), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(G264), .B(G1698), .C1(new_n327), .C2(new_n328), .ZN(new_n457));
  OAI211_X1 g0257(.A(G257), .B(new_n405), .C1(new_n327), .C2(new_n328), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n258), .A2(G303), .A3(new_n259), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n271), .ZN(new_n461));
  OR2_X1    g0261(.A1(KEYINPUT70), .A2(G41), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT5), .B1(new_n462), .B2(new_n273), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT5), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n208), .B(G45), .C1(new_n464), .C2(G41), .ZN(new_n465));
  OAI211_X1 g0265(.A(G270), .B(new_n280), .C1(new_n463), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n462), .A2(new_n273), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n465), .B1(new_n467), .B2(new_n464), .ZN(new_n468));
  INV_X1    g0268(.A(new_n280), .ZN(new_n469));
  INV_X1    g0269(.A(G274), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n461), .A2(new_n466), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n208), .A2(G33), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n304), .A2(G116), .A3(new_n289), .A4(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n295), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(G20), .B1(G33), .B2(G283), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n257), .A2(G97), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n478), .A2(new_n479), .B1(G20), .B2(new_n476), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n480), .A2(new_n335), .A3(KEYINPUT20), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT20), .B1(new_n480), .B2(new_n335), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n475), .B(new_n477), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n473), .A2(new_n483), .A3(G169), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT21), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n464), .B1(new_n274), .B2(new_n275), .ZN(new_n487));
  INV_X1    g0287(.A(new_n465), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n469), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n489), .A2(G270), .B1(new_n468), .B2(new_n471), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n314), .B1(new_n490), .B2(new_n461), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(KEYINPUT21), .A3(new_n483), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT84), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n461), .A2(G179), .A3(new_n472), .A4(new_n466), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n493), .B1(new_n495), .B2(new_n483), .ZN(new_n496));
  INV_X1    g0296(.A(new_n483), .ZN(new_n497));
  NOR3_X1   g0297(.A1(new_n497), .A2(KEYINPUT84), .A3(new_n494), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n486), .B(new_n492), .C1(new_n496), .C2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n483), .B1(G200), .B2(new_n473), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(new_n369), .B2(new_n473), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  OAI211_X1 g0304(.A(G250), .B(G1698), .C1(new_n327), .C2(new_n328), .ZN(new_n505));
  OAI211_X1 g0305(.A(G244), .B(new_n405), .C1(new_n327), .C2(new_n328), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n504), .B(new_n505), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT4), .B1(new_n260), .B2(G244), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n271), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n489), .A2(G257), .B1(new_n468), .B2(new_n471), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n314), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n510), .A2(new_n511), .A3(new_n362), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n341), .A2(G107), .A3(new_n347), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n390), .A2(KEYINPUT6), .A3(G97), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n227), .A2(new_n390), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n517), .A2(new_n205), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n516), .B1(new_n518), .B2(KEYINPUT6), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(G20), .B1(G77), .B2(new_n300), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n304), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n295), .A2(new_n227), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n292), .A2(new_n474), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(new_n227), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n513), .B(new_n514), .C1(new_n521), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n515), .A2(new_n520), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n335), .ZN(new_n527));
  INV_X1    g0327(.A(new_n524), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n510), .A2(new_n511), .A3(new_n369), .ZN(new_n529));
  AOI21_X1  g0329(.A(G200), .B1(new_n510), .B2(new_n511), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n527), .B(new_n528), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(G244), .B(G1698), .C1(new_n327), .C2(new_n328), .ZN(new_n533));
  OAI211_X1 g0333(.A(G238), .B(new_n405), .C1(new_n327), .C2(new_n328), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n534), .C1(new_n257), .C2(new_n476), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n271), .ZN(new_n536));
  INV_X1    g0336(.A(G250), .ZN(new_n537));
  INV_X1    g0337(.A(G45), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(G1), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n208), .A2(new_n470), .A3(G45), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n280), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n314), .ZN(new_n543));
  INV_X1    g0343(.A(new_n541), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n535), .B2(new_n271), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n362), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n378), .A2(new_n289), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT19), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n209), .B1(new_n404), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(G87), .B2(new_n206), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n209), .B(G68), .C1(new_n327), .C2(new_n328), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n548), .B1(new_n298), .B2(new_n227), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n547), .B1(new_n553), .B2(new_n335), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n292), .A2(new_n378), .A3(new_n474), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n554), .A2(KEYINPUT82), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT82), .B1(new_n554), .B2(new_n555), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n543), .B(new_n546), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT83), .B1(new_n542), .B2(new_n369), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT83), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n545), .A2(new_n560), .A3(G190), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n292), .A2(G87), .A3(new_n474), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n542), .A2(G200), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n559), .A2(new_n561), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n558), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n209), .B(G87), .C1(new_n327), .C2(new_n328), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT22), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT22), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n263), .A2(new_n569), .A3(new_n209), .A4(G87), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT24), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n257), .A2(new_n476), .A3(G20), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT23), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n209), .B2(G107), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n390), .A2(KEYINPUT23), .A3(G20), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n571), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n572), .B1(new_n571), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n335), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n523), .A2(new_n390), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT25), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n289), .B2(G107), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n295), .A2(KEYINPUT25), .A3(new_n390), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(G264), .B(new_n280), .C1(new_n463), .C2(new_n465), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n472), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n537), .A2(new_n405), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n228), .A2(G1698), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n327), .C2(new_n328), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT85), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G294), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n271), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n592), .B1(new_n591), .B2(new_n593), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT86), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n588), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT86), .B1(new_n595), .B2(new_n596), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n314), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT87), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n489), .A2(new_n602), .A3(G264), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n587), .A2(KEYINPUT87), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n603), .B(new_n604), .C1(new_n596), .C2(new_n595), .ZN(new_n605));
  INV_X1    g0405(.A(G179), .ZN(new_n606));
  INV_X1    g0406(.A(new_n472), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n586), .B1(new_n601), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n580), .A2(new_n585), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n371), .B1(new_n605), .B2(new_n607), .ZN(new_n611));
  INV_X1    g0411(.A(new_n596), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n612), .A2(new_n598), .A3(new_n271), .A4(new_n594), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n472), .A2(new_n587), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n600), .A2(new_n613), .A3(new_n614), .A4(new_n369), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n532), .A2(new_n566), .A3(new_n609), .A4(new_n617), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n456), .A2(new_n503), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g0419(.A(new_n619), .B(KEYINPUT88), .Z(G372));
  NAND2_X1  g0420(.A1(new_n398), .A2(KEYINPUT91), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT91), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n396), .A2(new_n397), .A3(new_n622), .A4(new_n386), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n448), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n376), .B1(new_n624), .B2(new_n445), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT90), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n366), .B2(new_n367), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n350), .A2(new_n365), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT18), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n350), .A2(new_n365), .A3(KEYINPUT18), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(KEYINPUT90), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n313), .B1(new_n625), .B2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n634), .A2(new_n317), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n525), .A2(new_n531), .A3(new_n558), .A4(new_n565), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n586), .B1(new_n615), .B2(new_n611), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT89), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT89), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n532), .A2(new_n566), .A3(new_n639), .A4(new_n617), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n500), .A2(new_n609), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n558), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n558), .A2(new_n565), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(new_n525), .ZN(new_n646));
  INV_X1    g0446(.A(new_n525), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n647), .A2(KEYINPUT26), .A3(new_n558), .A4(new_n565), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n643), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n635), .B1(new_n456), .B2(new_n651), .ZN(G369));
  NAND3_X1  g0452(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n653));
  OAI21_X1  g0453(.A(G213), .B1(new_n653), .B2(KEYINPUT27), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT92), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n653), .A2(KEYINPUT92), .A3(KEYINPUT27), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(new_n497), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n499), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n503), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n609), .A2(new_n617), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n610), .B2(new_n663), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n609), .B2(new_n663), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n500), .A2(new_n662), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n613), .A2(new_n614), .ZN(new_n675));
  INV_X1    g0475(.A(new_n600), .ZN(new_n676));
  OAI21_X1  g0476(.A(G169), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n594), .A2(new_n271), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n678), .A2(new_n612), .B1(KEYINPUT87), .B2(new_n587), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n679), .A2(G179), .A3(new_n472), .A4(new_n603), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n677), .A2(new_n680), .B1(new_n580), .B2(new_n585), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n674), .A2(new_n670), .B1(new_n681), .B2(new_n663), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n673), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT93), .ZN(G399));
  INV_X1    g0484(.A(new_n212), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n467), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n223), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT94), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT28), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n662), .B1(new_n642), .B2(new_n649), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(KEYINPUT29), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n636), .A2(new_n637), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT97), .B1(new_n499), .B2(new_n681), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT97), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT84), .B1(new_n497), .B2(new_n494), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n495), .A2(new_n493), .A3(new_n483), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT21), .B1(new_n491), .B2(new_n483), .ZN(new_n701));
  AND4_X1   g0501(.A1(KEYINPUT21), .A2(new_n473), .A3(new_n483), .A4(G169), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n609), .A2(new_n697), .A3(new_n700), .A4(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n695), .A2(new_n696), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n662), .B1(new_n705), .B2(new_n649), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n694), .B1(KEYINPUT29), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G330), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n669), .A2(new_n636), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n703), .A2(new_n700), .A3(new_n502), .A4(new_n663), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n709), .A2(KEYINPUT96), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT96), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n618), .B2(new_n710), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n662), .A2(KEYINPUT31), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n545), .A2(new_n490), .A3(G179), .A4(new_n461), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n717), .A2(new_n605), .A3(new_n512), .ZN(new_n718));
  AND4_X1   g0518(.A1(new_n362), .A2(new_n512), .A3(new_n473), .A4(new_n542), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n679), .A2(new_n472), .A3(new_n603), .ZN(new_n720));
  AOI22_X1  g0520(.A1(KEYINPUT30), .A2(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n679), .A2(new_n603), .A3(new_n510), .A4(new_n511), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n717), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n716), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT95), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n718), .B2(KEYINPUT30), .ZN(new_n727));
  OAI211_X1 g0527(.A(KEYINPUT95), .B(new_n722), .C1(new_n723), .C2(new_n717), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n719), .A2(new_n720), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n718), .A2(KEYINPUT30), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n727), .A2(new_n728), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n662), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT31), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n725), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n708), .B1(new_n715), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n707), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n692), .B1(new_n736), .B2(G1), .ZN(G364));
  AND2_X1   g0537(.A1(new_n209), .A2(G13), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n208), .B1(new_n738), .B2(G45), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n686), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n668), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(G330), .B2(new_n666), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n212), .A2(new_n263), .ZN(new_n744));
  INV_X1    g0544(.A(G355), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n744), .A2(new_n745), .B1(G116), .B2(new_n212), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n685), .A2(new_n263), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n224), .B2(new_n538), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n251), .A2(new_n538), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n220), .B1(G20), .B2(new_n314), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n741), .B1(new_n751), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n209), .A2(new_n371), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n316), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n369), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n209), .A2(new_n369), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n316), .A2(new_n371), .A3(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(G50), .A2(new_n761), .B1(new_n764), .B2(G58), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n209), .A2(G190), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n316), .A2(new_n371), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n765), .B1(new_n262), .B2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT98), .Z(new_n769));
  NOR2_X1   g0569(.A1(new_n371), .A2(G179), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G87), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n762), .A2(new_n770), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n263), .B1(new_n771), .B2(new_n390), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G179), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n766), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  OR3_X1    g0577(.A1(new_n776), .A2(KEYINPUT32), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(KEYINPUT32), .B1(new_n776), .B2(new_n777), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n209), .B1(new_n775), .B2(G190), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n778), .B(new_n779), .C1(new_n227), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n760), .A2(G190), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n774), .B(new_n781), .C1(G68), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n769), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G303), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n329), .B1(new_n773), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G283), .ZN(new_n787));
  INV_X1    g0587(.A(G329), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n771), .A2(new_n787), .B1(new_n776), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n780), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n786), .B(new_n789), .C1(G294), .C2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(KEYINPUT33), .B(G317), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n782), .A2(new_n792), .B1(new_n764), .B2(G322), .ZN(new_n793));
  INV_X1    g0593(.A(new_n767), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n761), .A2(G326), .B1(new_n794), .B2(G311), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n791), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n784), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n758), .B1(new_n797), .B2(new_n752), .ZN(new_n798));
  INV_X1    g0598(.A(new_n755), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n666), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n743), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G396));
  NAND4_X1  g0602(.A1(new_n621), .A2(new_n386), .A3(new_n623), .A4(new_n662), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n386), .A2(new_n662), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n395), .A2(new_n398), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n693), .B(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n735), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n741), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n808), .B2(new_n807), .ZN(new_n810));
  INV_X1    g0610(.A(new_n752), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n754), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT99), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n741), .B1(new_n813), .B2(G77), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n329), .B1(new_n776), .B2(new_n815), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n773), .A2(new_n390), .B1(new_n771), .B2(new_n772), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n816), .B(new_n817), .C1(G97), .C2(new_n790), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G303), .A2(new_n761), .B1(new_n764), .B2(G294), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n782), .A2(G283), .B1(new_n794), .B2(G116), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G137), .A2(new_n761), .B1(new_n782), .B2(G150), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT100), .ZN(new_n823));
  INV_X1    g0623(.A(G143), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n824), .B2(new_n763), .C1(new_n777), .C2(new_n767), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT34), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n263), .B1(new_n773), .B2(new_n202), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n771), .A2(new_n342), .B1(new_n776), .B2(new_n829), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n828), .B(new_n830), .C1(G58), .C2(new_n790), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n825), .B2(new_n826), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n821), .B1(new_n827), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n814), .B1(new_n833), .B2(new_n752), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n754), .B2(new_n806), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n810), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G384));
  AOI21_X1  g0637(.A(new_n659), .B1(new_n627), .B2(new_n632), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT103), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n444), .A2(new_n839), .A3(new_n662), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n839), .B1(new_n444), .B2(new_n662), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n412), .B1(new_n421), .B2(new_n423), .ZN(new_n844));
  OAI21_X1  g0644(.A(G169), .B1(new_n844), .B2(new_n414), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n428), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n426), .A2(KEYINPUT14), .A3(G169), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n846), .A2(new_n847), .B1(new_n419), .B2(G179), .ZN(new_n848));
  INV_X1    g0648(.A(new_n444), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n448), .B(new_n843), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT104), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT104), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n445), .A2(new_n852), .A3(new_n448), .A4(new_n843), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n848), .A2(new_n448), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n855), .A2(new_n444), .A3(new_n662), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n693), .A2(new_n806), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n398), .A2(new_n662), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n858), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT38), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT16), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n201), .B1(new_n346), .B2(G58), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n865), .A2(new_n209), .B1(new_n777), .B2(new_n301), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n342), .B1(new_n339), .B2(new_n331), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(new_n334), .A3(new_n335), .ZN(new_n869));
  INV_X1    g0669(.A(new_n322), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n660), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n630), .A2(new_n631), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n374), .B(KEYINPUT17), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n350), .A2(new_n659), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n628), .A2(new_n876), .A3(new_n877), .A4(new_n374), .ZN(new_n878));
  INV_X1    g0678(.A(new_n374), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n364), .A2(new_n660), .B1(new_n869), .B2(new_n870), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT37), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n863), .B1(new_n875), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n871), .B1(new_n368), .B2(new_n376), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n878), .A2(new_n881), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n838), .B1(new_n862), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n883), .A2(new_n886), .A3(KEYINPUT39), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n445), .A2(new_n662), .ZN(new_n890));
  INV_X1    g0690(.A(new_n886), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n628), .A2(new_n876), .A3(new_n374), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n876), .A2(new_n626), .A3(new_n374), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT37), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n892), .B1(KEYINPUT37), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT105), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n350), .A2(new_n659), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(new_n879), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n898), .B(new_n628), .C1(new_n626), .C2(new_n877), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT105), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT37), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n627), .A2(new_n632), .A3(new_n874), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n897), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n896), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n891), .B1(new_n905), .B2(new_n863), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n889), .B(new_n890), .C1(new_n906), .C2(KEYINPUT39), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n888), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n455), .A2(new_n707), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n635), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n908), .B(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n905), .A2(new_n863), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n886), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n731), .A2(KEYINPUT31), .A3(new_n662), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT31), .B1(new_n731), .B2(new_n662), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n715), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n803), .A2(new_n805), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n854), .B2(new_n856), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n917), .A2(KEYINPUT40), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n913), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n917), .A2(new_n919), .A3(new_n887), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n455), .A2(new_n917), .ZN(new_n926));
  OAI21_X1  g0726(.A(G330), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n925), .B2(new_n926), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n911), .A2(new_n928), .B1(new_n208), .B2(new_n738), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n911), .B2(new_n928), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n931), .A2(G116), .A3(new_n221), .A4(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(KEYINPUT101), .B(KEYINPUT36), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n933), .B(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n223), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n936), .B(G77), .C1(new_n324), .C2(new_n232), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n342), .A2(G50), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT102), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n208), .B(G13), .C1(new_n937), .C2(new_n939), .ZN(new_n940));
  OR3_X1    g0740(.A1(new_n930), .A2(new_n935), .A3(new_n940), .ZN(G367));
  OR2_X1    g0741(.A1(new_n663), .A2(new_n563), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n566), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n943), .A2(KEYINPUT106), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n558), .A2(new_n942), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(KEYINPUT106), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(new_n799), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n247), .A2(new_n748), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n756), .B1(new_n212), .B2(new_n379), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n741), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI22_X1  g0751(.A1(G150), .A2(new_n764), .B1(new_n794), .B2(G50), .ZN(new_n952));
  INV_X1    g0752(.A(new_n761), .ZN(new_n953));
  INV_X1    g0753(.A(new_n782), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n952), .B1(new_n824), .B2(new_n953), .C1(new_n777), .C2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n780), .A2(new_n342), .ZN(new_n956));
  INV_X1    g0756(.A(G137), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n263), .B1(new_n776), .B2(new_n957), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n773), .A2(new_n324), .B1(new_n771), .B2(new_n262), .ZN(new_n959));
  NOR4_X1   g0759(.A1(new_n955), .A2(new_n956), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n782), .A2(G294), .B1(new_n794), .B2(G283), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n815), .B2(new_n953), .ZN(new_n962));
  INV_X1    g0762(.A(new_n773), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n963), .A2(KEYINPUT46), .A3(G116), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT46), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n773), .B2(new_n476), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n964), .B(new_n966), .C1(new_n390), .C2(new_n780), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n763), .A2(new_n785), .ZN(new_n968));
  INV_X1    g0768(.A(G317), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n329), .B1(new_n776), .B2(new_n969), .C1(new_n227), .C2(new_n771), .ZN(new_n970));
  NOR4_X1   g0770(.A1(new_n962), .A2(new_n967), .A3(new_n968), .A4(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n960), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT47), .Z(new_n973));
  AOI21_X1  g0773(.A(new_n951), .B1(new_n973), .B2(new_n752), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n948), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n662), .B1(new_n521), .B2(new_n524), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n532), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n647), .A2(new_n662), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n682), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT45), .Z(new_n981));
  NOR2_X1   g0781(.A1(new_n682), .A2(new_n979), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT44), .ZN(new_n983));
  AND3_X1   g0783(.A1(new_n981), .A2(new_n673), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n673), .B1(new_n981), .B2(new_n983), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n674), .A2(new_n670), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n672), .B2(new_n674), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(new_n668), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n736), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n736), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n686), .B(KEYINPUT41), .Z(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n740), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n979), .A2(new_n670), .A3(new_n674), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT42), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n525), .B1(new_n977), .B2(new_n609), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n663), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(KEYINPUT42), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT107), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(KEYINPUT43), .B2(new_n947), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n947), .B(KEYINPUT43), .Z(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(new_n1004), .B2(new_n1002), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n979), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n673), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1005), .B(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n975), .B1(new_n995), .B2(new_n1008), .ZN(G387));
  NAND2_X1  g0809(.A1(new_n990), .A2(new_n740), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n688), .B(new_n538), .C1(new_n342), .C2(new_n262), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT108), .ZN(new_n1012));
  OAI21_X1  g0812(.A(KEYINPUT50), .B1(new_n297), .B2(G50), .ZN(new_n1013));
  OR3_X1    g0813(.A1(new_n297), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1011), .A2(KEYINPUT108), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n747), .B1(new_n1015), .B2(new_n1016), .C1(new_n243), .C2(new_n538), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(G107), .B2(new_n212), .C1(new_n688), .C2(new_n744), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n686), .B(new_n740), .C1(new_n1018), .C2(new_n756), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n776), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G77), .A2(new_n963), .B1(new_n1020), .B2(G150), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1021), .B(new_n263), .C1(new_n227), .C2(new_n771), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n782), .A2(new_n320), .B1(new_n794), .B2(G68), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n202), .B2(new_n763), .C1(new_n777), .C2(new_n953), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1022), .B(new_n1024), .C1(new_n378), .C2(new_n790), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n963), .A2(G294), .B1(new_n790), .B2(G283), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n785), .A2(new_n767), .B1(new_n763), .B2(new_n969), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1027), .A2(KEYINPUT109), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(KEYINPUT109), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G311), .A2(new_n782), .B1(new_n761), .B2(G322), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT48), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1026), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT110), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n1032), .B2(new_n1031), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(KEYINPUT49), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n263), .B1(new_n1020), .B2(G326), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n476), .B2(new_n771), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n1035), .B2(KEYINPUT49), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1025), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1019), .B1(new_n672), .B2(new_n799), .C1(new_n1040), .C2(new_n811), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n991), .A2(new_n686), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n736), .A2(new_n990), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1010), .B(new_n1041), .C1(new_n1042), .C2(new_n1043), .ZN(G393));
  NOR2_X1   g0844(.A1(new_n748), .A2(new_n254), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n756), .B1(new_n227), .B2(new_n212), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G283), .A2(new_n963), .B1(new_n1020), .B2(G322), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1047), .B(new_n329), .C1(new_n390), .C2(new_n771), .ZN(new_n1048));
  INV_X1    g0848(.A(G294), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n954), .A2(new_n785), .B1(new_n1049), .B2(new_n767), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1048), .B(new_n1050), .C1(G116), .C2(new_n790), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n953), .A2(new_n969), .B1(new_n815), .B2(new_n763), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT52), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n953), .A2(new_n299), .B1(new_n777), .B2(new_n763), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT51), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n954), .A2(new_n202), .B1(new_n297), .B2(new_n767), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n780), .A2(new_n262), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n263), .B1(new_n771), .B2(new_n772), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n773), .A2(new_n232), .B1(new_n776), .B2(new_n824), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1051), .A2(new_n1053), .B1(new_n1055), .B2(new_n1060), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n741), .B1(new_n1045), .B2(new_n1046), .C1(new_n1061), .C2(new_n811), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT111), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n799), .B2(new_n979), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n987), .B2(new_n739), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n987), .A2(new_n991), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n991), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n687), .B1(new_n1067), .B2(new_n986), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1065), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(G390));
  AOI21_X1  g0870(.A(KEYINPUT96), .B1(new_n709), .B2(new_n711), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n669), .A2(new_n710), .A3(new_n636), .A4(new_n713), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n734), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(G330), .A3(new_n806), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n708), .B1(new_n715), .B2(new_n916), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1074), .A2(new_n858), .B1(new_n1075), .B2(new_n919), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n860), .B1(new_n693), .B2(new_n806), .ZN(new_n1077));
  OAI21_X1  g0877(.A(KEYINPUT112), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT112), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1077), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n857), .B1(new_n735), .B2(new_n806), .ZN(new_n1081));
  AND3_X1   g0881(.A1(new_n917), .A2(G330), .A3(new_n919), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1079), .B(new_n1080), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1078), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n735), .A2(new_n806), .A3(new_n857), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n705), .A2(new_n649), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1086), .A2(new_n663), .A3(new_n806), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1085), .A2(new_n861), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n857), .B1(new_n1075), .B2(new_n806), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1084), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n455), .A2(new_n1075), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n909), .A2(new_n1092), .A3(new_n635), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n889), .B1(new_n906), .B2(KEYINPUT39), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1077), .A2(new_n858), .B1(new_n445), .B2(new_n662), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1087), .A2(new_n861), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n890), .B1(new_n1098), .B2(new_n857), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1096), .A2(new_n1097), .B1(new_n913), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n1085), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1082), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1095), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1074), .A2(new_n858), .ZN(new_n1105));
  AOI221_X4 g0905(.A(new_n1105), .B1(new_n1099), .B2(new_n913), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1099), .A2(new_n913), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1102), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1093), .B1(new_n1084), .B2(new_n1090), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1104), .A2(new_n686), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(G125), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n263), .B1(new_n776), .B2(new_n1114), .C1(new_n202), .C2(new_n771), .ZN(new_n1115));
  OR3_X1    g0915(.A1(new_n773), .A2(KEYINPUT53), .A3(new_n299), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT53), .B1(new_n773), .B2(new_n299), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(new_n777), .C2(new_n780), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1115), .B(new_n1118), .C1(G128), .C2(new_n761), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT54), .B(G143), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n829), .A2(new_n763), .B1(new_n767), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G137), .B2(new_n782), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n771), .A2(new_n342), .B1(new_n776), .B2(new_n1049), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n329), .B1(new_n773), .B2(new_n772), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n1057), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n953), .A2(new_n787), .B1(new_n227), .B2(new_n767), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n954), .A2(new_n390), .B1(new_n476), .B2(new_n763), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1119), .A2(new_n1122), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n741), .B1(new_n320), .B2(new_n813), .C1(new_n1129), .C2(new_n811), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n1096), .B2(new_n753), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n1110), .B2(new_n740), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1113), .A2(new_n1132), .ZN(G378));
  INV_X1    g0933(.A(KEYINPUT57), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n708), .B1(new_n922), .B2(new_n923), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n305), .A2(new_n659), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n318), .B(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1137), .B(new_n1139), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n921), .A2(new_n1135), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(new_n921), .B2(new_n1135), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n908), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT117), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1140), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n924), .A2(G330), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n917), .A2(new_n919), .A3(KEYINPUT40), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n906), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1145), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n888), .A2(new_n907), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n921), .A2(new_n1135), .A3(new_n1140), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1143), .A2(new_n1144), .A3(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1149), .A2(new_n1150), .A3(KEYINPUT117), .A4(new_n1151), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1093), .B1(new_n1110), .B2(new_n1091), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1134), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1150), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1159));
  OAI21_X1  g0959(.A(KEYINPUT57), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(KEYINPUT118), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n1078), .B2(new_n1083), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1094), .B1(new_n1103), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT118), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1134), .B1(new_n1143), .B2(new_n1152), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1157), .A2(new_n1161), .A3(new_n686), .A4(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1153), .A2(new_n740), .A3(new_n1154), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n761), .A2(G116), .B1(new_n794), .B2(new_n378), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n227), .B2(new_n954), .C1(new_n390), .C2(new_n763), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n773), .A2(new_n262), .B1(new_n776), .B2(new_n787), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n467), .A2(new_n263), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n324), .B2(new_n771), .ZN(new_n1174));
  NOR4_X1   g0974(.A1(new_n1171), .A2(new_n956), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT58), .Z(new_n1176));
  AOI22_X1  g0976(.A1(new_n761), .A2(G125), .B1(G150), .B2(new_n790), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT113), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n767), .A2(new_n957), .B1(new_n773), .B2(new_n1120), .ZN(new_n1179));
  INV_X1    g0979(.A(G128), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n954), .A2(new_n829), .B1(new_n1180), .B2(new_n763), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT59), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(G33), .A2(G41), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n771), .B2(new_n777), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G124), .B2(new_n1020), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1176), .B1(new_n1184), .B2(new_n1188), .C1(new_n1173), .C2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT114), .Z(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n752), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT115), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n741), .B1(new_n813), .B2(G50), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT116), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1193), .B(new_n1195), .C1(new_n754), .C2(new_n1145), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1169), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1168), .A2(new_n1197), .ZN(G375));
  OAI21_X1  g0998(.A(KEYINPUT119), .B1(new_n1163), .B2(new_n739), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT119), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1091), .A2(new_n1200), .A3(new_n740), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n741), .B1(new_n813), .B2(G68), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G97), .A2(new_n963), .B1(new_n1020), .B2(G303), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n787), .B2(new_n763), .C1(new_n379), .C2(new_n780), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n329), .B1(new_n771), .B2(new_n262), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT120), .Z(new_n1206));
  NOR2_X1   g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n782), .A2(G116), .B1(new_n794), .B2(G107), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(new_n1049), .C2(new_n953), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n263), .B1(new_n771), .B2(new_n324), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n773), .A2(new_n777), .B1(new_n776), .B2(new_n1180), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(G50), .C2(new_n790), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G132), .A2(new_n761), .B1(new_n764), .B2(G137), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1120), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n782), .A2(new_n1214), .B1(new_n794), .B2(G150), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1209), .A2(new_n1216), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1217), .A2(KEYINPUT121), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n811), .B1(new_n1217), .B2(KEYINPUT121), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1202), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n857), .B2(new_n754), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1199), .A2(new_n1201), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1163), .A2(new_n1093), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1095), .A2(new_n1224), .A3(new_n994), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(G381));
  NAND2_X1  g1026(.A1(G378), .A2(KEYINPUT123), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT123), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1113), .A2(new_n1228), .A3(new_n1132), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(G375), .A2(new_n1230), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT122), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n975), .B(new_n1069), .C1(new_n995), .C2(new_n1008), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1233), .A2(G381), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1231), .A2(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT124), .ZN(G407));
  INV_X1    g1037(.A(G213), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1231), .B2(new_n661), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(G407), .A2(new_n1239), .ZN(G409));
  XNOR2_X1  g1040(.A(G393), .B(new_n801), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(G387), .A2(G390), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT125), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1234), .A2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1241), .B1(new_n1243), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1241), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1242), .A2(new_n1244), .A3(new_n1234), .A4(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT61), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1238), .A2(G343), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1168), .A2(G378), .A3(new_n1197), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1164), .A2(new_n994), .A3(new_n1154), .A4(new_n1153), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n740), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1196), .A3(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1227), .A2(new_n1256), .A3(new_n1229), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1252), .B1(new_n1253), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1252), .A2(G2897), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1163), .A2(KEYINPUT60), .A3(new_n1093), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n686), .ZN(new_n1262));
  OAI21_X1  g1062(.A(KEYINPUT60), .B1(new_n1163), .B2(new_n1093), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n1224), .B2(new_n1263), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1264), .A2(new_n836), .A3(new_n1222), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1224), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(new_n686), .A3(new_n1261), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G384), .B1(new_n1267), .B2(new_n1223), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1260), .B1(new_n1265), .B2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n836), .B1(new_n1264), .B2(new_n1222), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1267), .A2(G384), .A3(new_n1223), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(new_n1271), .A3(new_n1259), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1251), .B1(new_n1258), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT62), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1275), .B1(new_n1258), .B2(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1274), .A2(new_n1278), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n1252), .B(new_n1276), .C1(new_n1253), .C2(new_n1257), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1275), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1250), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1258), .A2(KEYINPUT63), .A3(new_n1277), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1283), .B(new_n1251), .C1(new_n1258), .C2(new_n1273), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1250), .B1(new_n1280), .B2(KEYINPUT63), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT126), .B1(new_n1282), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT126), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1258), .A2(new_n1277), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1249), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1274), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1292), .A3(new_n1283), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1289), .A2(KEYINPUT62), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1294), .A2(new_n1274), .A3(new_n1278), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1288), .B(new_n1293), .C1(new_n1295), .C2(new_n1250), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1287), .A2(new_n1296), .ZN(G405));
  NAND2_X1  g1097(.A1(new_n1276), .A2(KEYINPUT127), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1249), .B(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(G375), .ZN(new_n1300));
  OAI221_X1 g1100(.A(new_n1253), .B1(KEYINPUT127), .B2(new_n1276), .C1(new_n1300), .C2(new_n1230), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1299), .B(new_n1301), .ZN(G402));
endmodule


