//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n564, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT67), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT68), .Z(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n463), .B(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(G137), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n469), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n470), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n472), .A2(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n469), .A2(KEYINPUT70), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n466), .A2(new_n468), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n478), .A2(G2105), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n478), .A2(new_n470), .A3(new_n481), .ZN(new_n485));
  OAI221_X1 g060(.A(new_n477), .B1(new_n482), .B2(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  INV_X1    g062(.A(KEYINPUT71), .ZN(new_n488));
  NAND2_X1  g063(.A1(G114), .A2(G2104), .ZN(new_n489));
  INV_X1    g064(.A(G126), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n479), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n462), .A2(G102), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR4_X1   g070(.A1(new_n479), .A2(KEYINPUT4), .A3(new_n495), .A4(G2105), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n495), .A2(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n469), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n488), .B1(new_n494), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n469), .A2(new_n498), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n469), .A2(new_n497), .A3(new_n498), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n491), .A2(G2105), .B1(G102), .B2(new_n462), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(KEYINPUT71), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n501), .A2(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n509), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT6), .B1(new_n511), .B2(KEYINPUT72), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n512), .A2(new_n519), .ZN(G166));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n516), .B1(new_n515), .B2(G651), .ZN(new_n522));
  NOR3_X1   g097(.A1(new_n511), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n514), .A2(new_n517), .A3(KEYINPUT73), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n524), .A2(G543), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT74), .B(G51), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n518), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(new_n509), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n528), .A2(new_n532), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND4_X1  g111(.A1(new_n524), .A2(G52), .A3(G543), .A4(new_n525), .ZN(new_n537));
  INV_X1    g112(.A(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT5), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT5), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n518), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G90), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n509), .A2(G64), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G651), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n550));
  OAI211_X1 g125(.A(new_n537), .B(new_n544), .C1(new_n549), .C2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  NAND3_X1  g127(.A1(new_n524), .A2(G543), .A3(new_n525), .ZN(new_n553));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n543), .A2(G81), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n542), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G651), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G188));
  NAND4_X1  g143(.A1(new_n524), .A2(G53), .A3(G543), .A4(new_n525), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n525), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n571), .A2(new_n572), .A3(G53), .A4(new_n524), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n542), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(G91), .A2(new_n543), .B1(new_n577), .B2(G651), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G166), .ZN(G303));
  NAND2_X1  g155(.A1(new_n543), .A2(G87), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(KEYINPUT76), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n509), .A2(G74), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n581), .A2(KEYINPUT76), .B1(G651), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n526), .A2(G49), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(new_n509), .A2(G61), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n511), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n589), .A2(KEYINPUT77), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n589), .A2(KEYINPUT77), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n509), .A2(G86), .ZN(new_n592));
  NAND2_X1  g167(.A1(G48), .A2(G543), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n590), .A2(new_n591), .B1(new_n518), .B2(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n511), .B1(new_n596), .B2(KEYINPUT78), .ZN(new_n597));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G60), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n542), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT78), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n597), .A2(new_n602), .B1(G85), .B2(new_n543), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n526), .A2(G47), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT79), .B(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n542), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G651), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n524), .A2(G54), .A3(G543), .A4(new_n525), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n509), .A2(G92), .A3(new_n514), .A4(new_n517), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n610), .B(new_n611), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT80), .Z(new_n617));
  OAI21_X1  g192(.A(new_n606), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n606), .B1(new_n617), .B2(G868), .ZN(G321));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(G299), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n620), .B2(G168), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(new_n620), .B2(G168), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n617), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n562), .ZN(G323));
  XOR2_X1   g203(.A(KEYINPUT81), .B(KEYINPUT11), .Z(new_n629));
  XNOR2_X1  g204(.A(G323), .B(new_n629), .ZN(G282));
  INV_X1    g205(.A(new_n482), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n631), .A2(KEYINPUT82), .A3(G123), .ZN(new_n632));
  INV_X1    g207(.A(new_n485), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G135), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT82), .ZN(new_n635));
  INV_X1    g210(.A(G123), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n482), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  INV_X1    g213(.A(G111), .ZN(new_n639));
  AOI22_X1  g214(.A1(new_n638), .A2(KEYINPUT83), .B1(new_n639), .B2(G2105), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(KEYINPUT83), .B2(new_n638), .ZN(new_n641));
  NAND4_X1  g216(.A1(new_n632), .A2(new_n634), .A3(new_n637), .A4(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n469), .A2(new_n462), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2100), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2435), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2443), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(G2446), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G1341), .B(G1348), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT84), .ZN(new_n662));
  INV_X1    g237(.A(G14), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n659), .B2(new_n660), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G401));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT85), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT17), .ZN(new_n669));
  XOR2_X1   g244(.A(G2067), .B(G2678), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT86), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2084), .B(G2090), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n671), .A2(new_n672), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n674), .B(new_n675), .C1(new_n673), .C2(new_n668), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n670), .A2(new_n672), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n668), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT18), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2096), .B(G2100), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT87), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1981), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n688), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n688), .A2(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n695));
  OAI221_X1 g270(.A(new_n693), .B1(new_n688), .B2(new_n691), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n695), .B2(new_n694), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(G1991), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1996), .ZN(new_n699));
  INV_X1    g274(.A(G1986), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G1996), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n698), .B(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n703), .A2(G1986), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n686), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(G1986), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n699), .A2(new_n700), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n706), .A2(new_n707), .A3(new_n685), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(new_n708), .ZN(G229));
  NOR2_X1   g284(.A1(G4), .A2(G16), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n617), .B2(G16), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1348), .ZN(new_n712));
  INV_X1    g287(.A(G1956), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT23), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G299), .B2(G16), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G20), .ZN(new_n717));
  MUX2_X1   g292(.A(new_n714), .B(new_n715), .S(new_n717), .Z(new_n718));
  AOI21_X1  g293(.A(new_n712), .B1(new_n713), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G35), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G162), .B2(new_n720), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n722), .A2(KEYINPUT29), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(KEYINPUT29), .ZN(new_n724));
  OR3_X1    g299(.A1(new_n723), .A2(new_n724), .A3(G2090), .ZN(new_n725));
  OAI21_X1  g300(.A(G2090), .B1(new_n723), .B2(new_n724), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n716), .A2(G19), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n562), .B2(new_n716), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(G1341), .Z(new_n729));
  AND3_X1   g304(.A1(new_n725), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n720), .A2(G26), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n631), .A2(G128), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n633), .A2(G140), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n470), .A2(G116), .ZN(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n733), .B(new_n734), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  AND3_X1   g312(.A1(new_n737), .A2(KEYINPUT94), .A3(G29), .ZN(new_n738));
  AOI21_X1  g313(.A(KEYINPUT94), .B1(new_n737), .B2(G29), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n732), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G2067), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n718), .A2(new_n713), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n719), .A2(new_n730), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(G168), .A2(G16), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G16), .B2(G21), .ZN(new_n746));
  INV_X1    g321(.A(G1966), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(KEYINPUT97), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n642), .A2(new_n720), .ZN(new_n750));
  AND2_X1   g325(.A1(KEYINPUT24), .A2(G34), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n720), .B1(KEYINPUT24), .B2(G34), .ZN(new_n752));
  OAI22_X1  g327(.A1(G160), .A2(new_n720), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(G2084), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(G2084), .ZN(new_n755));
  INV_X1    g330(.A(G28), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(KEYINPUT30), .ZN(new_n757));
  AOI21_X1  g332(.A(G29), .B1(new_n756), .B2(KEYINPUT30), .ZN(new_n758));
  OR2_X1    g333(.A1(KEYINPUT31), .A2(G11), .ZN(new_n759));
  NAND2_X1  g334(.A1(KEYINPUT31), .A2(G11), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n757), .A2(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n754), .A2(new_n755), .A3(new_n761), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n749), .A2(new_n750), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G1961), .ZN(new_n764));
  NAND2_X1  g339(.A1(G171), .A2(G16), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G5), .B2(G16), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n748), .A2(KEYINPUT97), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G27), .A2(G29), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G164), .B2(G29), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT99), .B(G2078), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(G29), .A2(G32), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT26), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n775), .A2(new_n776), .B1(G105), .B2(new_n462), .ZN(new_n777));
  INV_X1    g352(.A(G129), .ZN(new_n778));
  INV_X1    g353(.A(G141), .ZN(new_n779));
  OAI221_X1 g354(.A(new_n777), .B1(new_n482), .B2(new_n778), .C1(new_n779), .C2(new_n485), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n772), .B1(new_n780), .B2(new_n720), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT27), .B(G1996), .Z(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n781), .A2(new_n783), .ZN(new_n785));
  AOI211_X1 g360(.A(new_n784), .B(new_n785), .C1(new_n747), .C2(new_n746), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n763), .A2(new_n767), .A3(new_n771), .A4(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(G33), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(G29), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n462), .A2(G103), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT25), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n633), .B2(G139), .ZN(new_n792));
  NAND2_X1  g367(.A1(G115), .A2(G2104), .ZN(new_n793));
  INV_X1    g368(.A(G127), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n479), .B2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT95), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(G2105), .B1(new_n795), .B2(new_n796), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n792), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n789), .B1(new_n799), .B2(G29), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n800), .A2(new_n801), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(G2072), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n766), .A2(new_n764), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(KEYINPUT98), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n805), .B2(G2072), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(KEYINPUT98), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n806), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n787), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT100), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT100), .B1(new_n787), .B2(new_n811), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n744), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(KEYINPUT93), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(G95), .A2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n820), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT88), .ZN(new_n822));
  INV_X1    g397(.A(G119), .ZN(new_n823));
  INV_X1    g398(.A(G131), .ZN(new_n824));
  OAI221_X1 g399(.A(new_n822), .B1(new_n482), .B2(new_n823), .C1(new_n824), .C2(new_n485), .ZN(new_n825));
  MUX2_X1   g400(.A(G25), .B(new_n825), .S(G29), .Z(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT35), .B(G1991), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n716), .A2(G24), .ZN(new_n829));
  INV_X1    g404(.A(G290), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n716), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G1986), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(G16), .A2(G22), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G166), .B2(G16), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT91), .B(G1971), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(G305), .A2(G16), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G6), .B2(new_n716), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT32), .B(G1981), .Z(new_n840));
  AOI21_X1  g415(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(G16), .A2(G23), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT89), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(G288), .B2(new_n716), .ZN(new_n844));
  XNOR2_X1  g419(.A(KEYINPUT90), .B(KEYINPUT33), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G1976), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n844), .B(new_n846), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n841), .B(new_n847), .C1(new_n839), .C2(new_n840), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n833), .B1(new_n848), .B2(KEYINPUT34), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT92), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n833), .B(KEYINPUT92), .C1(new_n848), .C2(KEYINPUT34), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n848), .A2(KEYINPUT34), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n819), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n853), .A2(new_n854), .A3(new_n819), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n816), .B1(new_n855), .B2(new_n856), .ZN(G150));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n858));
  NAND2_X1  g433(.A1(G150), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n816), .B(KEYINPUT101), .C1(new_n855), .C2(new_n856), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(G311));
  NAND2_X1  g436(.A1(new_n617), .A2(G559), .ZN(new_n862));
  XOR2_X1   g437(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n863));
  XOR2_X1   g438(.A(new_n862), .B(new_n863), .Z(new_n864));
  AND2_X1   g439(.A1(new_n556), .A2(new_n560), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n526), .A2(G43), .ZN(new_n866));
  INV_X1    g441(.A(G55), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n553), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n543), .A2(G93), .ZN(new_n869));
  NAND2_X1  g444(.A1(G80), .A2(G543), .ZN(new_n870));
  INV_X1    g445(.A(G67), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n542), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(G651), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n865), .B(new_n866), .C1(new_n868), .C2(new_n874), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n869), .A2(new_n873), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n526), .A2(G55), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n876), .B(new_n877), .C1(new_n555), .C2(new_n561), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(KEYINPUT39), .Z(new_n880));
  AOI21_X1  g455(.A(G860), .B1(new_n864), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n864), .B2(new_n880), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n868), .A2(new_n874), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G860), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT37), .Z(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(new_n886), .ZN(G145));
  XNOR2_X1  g462(.A(new_n642), .B(new_n486), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(G160), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n891));
  INV_X1    g466(.A(G118), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n890), .A2(new_n891), .B1(new_n892), .B2(G2105), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n891), .B2(new_n890), .ZN(new_n894));
  INV_X1    g469(.A(G130), .ZN(new_n895));
  INV_X1    g470(.A(G142), .ZN(new_n896));
  OAI221_X1 g471(.A(new_n894), .B1(new_n482), .B2(new_n895), .C1(new_n896), .C2(new_n485), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n825), .B(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n780), .B(new_n645), .Z(new_n900));
  OR2_X1    g475(.A1(new_n900), .A2(new_n799), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n799), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n505), .A2(new_n506), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n737), .B(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n901), .B2(new_n902), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n899), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n908), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n898), .A3(new_n906), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n889), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G37), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n913), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n909), .A2(new_n911), .A3(new_n889), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n914), .A2(new_n915), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT40), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT40), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n917), .A2(new_n915), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n914), .A2(new_n920), .A3(new_n916), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n922), .ZN(G395));
  XNOR2_X1  g498(.A(G290), .B(G305), .ZN(new_n924));
  XNOR2_X1  g499(.A(G288), .B(G166), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n924), .B(new_n925), .Z(new_n926));
  NAND2_X1  g501(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n927));
  OR2_X1    g502(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n924), .B(new_n925), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n930), .A2(KEYINPUT107), .A3(KEYINPUT42), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n879), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n626), .B(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n616), .ZN(new_n935));
  NAND2_X1  g510(.A1(G299), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n574), .A2(new_n616), .A3(new_n578), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n574), .A2(new_n616), .A3(new_n578), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n616), .B1(new_n574), .B2(new_n578), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT105), .B1(new_n942), .B2(KEYINPUT41), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT41), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n938), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n942), .B2(KEYINPUT41), .ZN(new_n948));
  NOR4_X1   g523(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT106), .A4(new_n945), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n943), .B(new_n946), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n939), .B1(new_n951), .B2(new_n934), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n932), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n932), .B2(new_n952), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n953), .B1(new_n932), .B2(new_n952), .ZN(new_n956));
  OAI21_X1  g531(.A(G868), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n884), .A2(new_n620), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT109), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n961), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(G295));
  NAND2_X1  g538(.A1(new_n959), .A2(KEYINPUT110), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n957), .A2(new_n965), .A3(new_n958), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(G331));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  AOI21_X1  g543(.A(G286), .B1(G171), .B2(KEYINPUT111), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n971));
  NAND2_X1  g546(.A1(G301), .A2(new_n971), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n972), .A2(new_n875), .A3(new_n878), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n972), .B1(new_n875), .B2(new_n878), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n972), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n879), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n972), .A2(new_n875), .A3(new_n878), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n969), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n981), .A3(new_n938), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n975), .A2(new_n979), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT112), .B1(new_n950), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(new_n938), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n926), .B(new_n982), .C1(new_n984), .C2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n915), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n944), .B1(new_n938), .B2(new_n945), .ZN(new_n989));
  AOI211_X1 g564(.A(KEYINPUT105), .B(KEYINPUT41), .C1(new_n936), .C2(new_n937), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT106), .B1(new_n938), .B2(new_n945), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n942), .A2(new_n947), .A3(KEYINPUT41), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n980), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n985), .B1(new_n995), .B2(KEYINPUT112), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n926), .B1(new_n996), .B2(new_n982), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n968), .B1(new_n988), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT113), .B1(new_n942), .B2(KEYINPUT41), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n999), .A2(KEYINPUT41), .A3(new_n942), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n983), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n999), .B1(KEYINPUT41), .B2(new_n942), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n985), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(G37), .B1(new_n1003), .B2(new_n930), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(KEYINPUT43), .A3(new_n987), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n998), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT44), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT43), .B1(new_n988), .B2(new_n997), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(new_n968), .A3(new_n987), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1007), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1011), .B1(new_n998), .B2(new_n1005), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT44), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT114), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(new_n1017), .ZN(G397));
  XNOR2_X1  g593(.A(new_n737), .B(G2067), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n1019), .A2(new_n780), .ZN(new_n1020));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n494), .B2(new_n500), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G40), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n472), .A2(new_n474), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT46), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n702), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1020), .A2(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1032));
  XOR2_X1   g607(.A(new_n1032), .B(KEYINPUT47), .Z(new_n1033));
  XNOR2_X1  g608(.A(new_n780), .B(G1996), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n825), .A2(new_n827), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n825), .A2(new_n827), .ZN(new_n1036));
  NOR4_X1   g611(.A1(new_n1019), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1028), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1028), .A2(new_n700), .A3(new_n830), .ZN(new_n1040));
  XOR2_X1   g615(.A(new_n1040), .B(KEYINPUT48), .Z(new_n1041));
  NOR2_X1   g616(.A1(new_n737), .A2(G2067), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1019), .A2(new_n1034), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1042), .B1(new_n1043), .B2(new_n1036), .ZN(new_n1044));
  OAI22_X1  g619(.A1(new_n1039), .A2(new_n1041), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1033), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT63), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n501), .A2(new_n1021), .A3(new_n507), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1027), .B1(new_n1048), .B2(KEYINPUT50), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1384), .B1(new_n505), .B2(new_n506), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI211_X1 g628(.A(KEYINPUT115), .B(G1384), .C1(new_n505), .C2(new_n506), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1050), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1049), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(G2090), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1048), .A2(new_n1023), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n903), .A2(KEYINPUT45), .A3(new_n1021), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1059), .A2(new_n1026), .ZN(new_n1060));
  AOI21_X1  g635(.A(G1971), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT116), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1061), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1063), .B(new_n1064), .C1(G2090), .C2(new_n1056), .ZN(new_n1065));
  NAND2_X1  g640(.A1(G303), .A2(G8), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(KEYINPUT55), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1062), .A2(new_n1065), .A3(G8), .A4(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT118), .B(G1981), .ZN(new_n1070));
  OR2_X1    g645(.A1(G305), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n594), .A2(new_n518), .ZN(new_n1072));
  OAI21_X1  g647(.A(G1981), .B1(new_n1072), .B2(new_n589), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT49), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1026), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1071), .A2(KEYINPUT49), .A3(new_n1073), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1076), .A2(G8), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G288), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G1976), .ZN(new_n1081));
  INV_X1    g656(.A(G1976), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT52), .B1(G288), .B2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1077), .A2(new_n1081), .A3(G8), .A4(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT117), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1079), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1077), .A2(G8), .A3(new_n1081), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT52), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT117), .B1(new_n1088), .B2(new_n1084), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1026), .B1(new_n1048), .B2(KEYINPUT50), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1053), .A2(new_n1054), .A3(new_n1050), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1091), .A2(new_n1092), .A3(G2090), .ZN(new_n1093));
  OAI21_X1  g668(.A(G8), .B1(new_n1093), .B2(new_n1061), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n1067), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1069), .A2(new_n1090), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G8), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1022), .A2(KEYINPUT115), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(new_n1023), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n1021), .A4(new_n507), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1026), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n747), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G2084), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1049), .A2(new_n1055), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1097), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(G168), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1047), .B1(new_n1096), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1062), .A2(G8), .A3(new_n1065), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1067), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1108), .A2(new_n1047), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1111), .A2(new_n1069), .A3(new_n1090), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1077), .A2(G8), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1079), .A2(new_n1082), .A3(new_n1080), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1115), .B1(new_n1116), .B2(new_n1071), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1069), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n1118), .B2(new_n1090), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1114), .A2(new_n1119), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n935), .A2(KEYINPUT60), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1077), .B2(G2067), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1124), .A2(KEYINPUT119), .A3(new_n741), .A4(new_n1026), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1348), .B1(new_n1049), .B2(new_n1055), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1121), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1127), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n616), .B(KEYINPUT60), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1129), .A2(new_n1125), .A3(new_n1123), .A4(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n713), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT56), .B(G2072), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1058), .A2(new_n1060), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(G299), .B(KEYINPUT57), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT61), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1137), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1133), .A2(new_n1135), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT123), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT122), .B1(new_n1145), .B2(KEYINPUT121), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1058), .A2(new_n1060), .A3(new_n702), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT58), .B(G1341), .Z(new_n1148));
  NAND2_X1  g723(.A1(new_n1077), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1146), .B1(new_n1150), .B2(new_n562), .ZN(new_n1151));
  INV_X1    g726(.A(new_n562), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1146), .B1(KEYINPUT122), .B2(new_n1145), .ZN(new_n1153));
  AOI211_X1 g728(.A(new_n1152), .B(new_n1153), .C1(new_n1147), .C2(new_n1149), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1139), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1140), .B(new_n1142), .C1(new_n1156), .C2(KEYINPUT61), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1132), .A2(new_n1144), .A3(new_n1155), .A4(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1159), .A2(new_n616), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n1137), .B(KEYINPUT120), .Z(new_n1161));
  AOI22_X1  g736(.A1(new_n1160), .A2(new_n1140), .B1(new_n1136), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(G2078), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1100), .A2(new_n1164), .A3(new_n1026), .A4(new_n1102), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT125), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1103), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1167), .A2(new_n1168), .A3(new_n1164), .A4(new_n1100), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1166), .A2(new_n1169), .A3(KEYINPUT53), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1058), .A2(new_n1060), .A3(new_n1164), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT53), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1056), .A2(new_n764), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(G301), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1174), .A2(KEYINPUT126), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n1176));
  AOI211_X1 g751(.A(new_n1176), .B(G301), .C1(new_n1170), .C2(new_n1173), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1060), .A2(KEYINPUT53), .A3(new_n1164), .A4(new_n1024), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1173), .A2(G301), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1175), .A2(new_n1177), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1183), .B1(new_n1173), .B2(new_n1178), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1056), .A2(new_n764), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1186));
  AND4_X1   g761(.A1(new_n1183), .A2(new_n1185), .A3(new_n1186), .A4(new_n1178), .ZN(new_n1187));
  OAI21_X1  g762(.A(G171), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1180), .B1(new_n1189), .B2(G301), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1163), .B1(new_n1182), .B2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1174), .B(KEYINPUT126), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT124), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1195), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1104), .A2(new_n1195), .A3(new_n1106), .ZN(new_n1198));
  AOI21_X1  g773(.A(G286), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT51), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1200), .A2(new_n1097), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1201), .ZN(new_n1202));
  OAI22_X1  g777(.A1(new_n1199), .A2(new_n1202), .B1(KEYINPUT51), .B2(new_n1107), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1198), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1201), .B1(new_n1204), .B2(new_n1196), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1205), .A2(G8), .A3(G286), .ZN(new_n1206));
  AOI22_X1  g781(.A1(new_n1193), .A2(new_n1194), .B1(new_n1203), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1192), .A2(new_n1207), .ZN(new_n1208));
  AND2_X1   g783(.A1(new_n1203), .A2(new_n1206), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1193), .A2(KEYINPUT62), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1096), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1120), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g787(.A(G290), .B(new_n700), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1038), .B1(new_n1037), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1046), .B1(new_n1212), .B2(new_n1214), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g790(.A1(G227), .A2(new_n459), .ZN(new_n1217));
  AND4_X1   g791(.A1(new_n665), .A2(new_n705), .A3(new_n708), .A4(new_n1217), .ZN(new_n1218));
  NAND3_X1  g792(.A1(new_n1218), .A2(new_n918), .A3(new_n1010), .ZN(G225));
  INV_X1    g793(.A(G225), .ZN(G308));
endmodule


