//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1250, new_n1251, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1323,
    new_n1324;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND3_X1  g0012(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT65), .B(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n212), .B(new_n222), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G97), .B(G107), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n202), .A2(G68), .ZN(new_n245));
  INV_X1    g0045(.A(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n244), .B(new_n250), .ZN(G351));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  AOI22_X1  g0052(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT8), .A2(G58), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT67), .A2(G58), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT67), .A2(G58), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT8), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n255), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n217), .A2(G33), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n253), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G1), .A2(G13), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT64), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(new_n213), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G13), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n268), .A2(new_n207), .A3(G1), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n262), .A2(new_n267), .B1(new_n202), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n267), .A2(new_n269), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(G1), .B2(new_n207), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n270), .B1(new_n202), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT9), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n263), .B1(G33), .B2(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n277), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n278), .B1(G226), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n279), .B1(new_n214), .B2(new_n215), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G222), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G223), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n286), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n285), .B(new_n290), .C1(G77), .C2(new_n286), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n283), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(G200), .B2(new_n292), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n274), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n283), .A2(new_n291), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n273), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n233), .A2(G1698), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(G226), .B2(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT3), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G33), .ZN(new_n306));
  INV_X1    g0106(.A(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G97), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n304), .A2(new_n309), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n278), .B1(new_n311), .B2(new_n285), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT13), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT68), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n281), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n280), .A2(KEYINPUT68), .A3(new_n277), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(G238), .A3(new_n316), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n312), .A2(new_n313), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n313), .B1(new_n312), .B2(new_n317), .ZN(new_n319));
  OAI21_X1  g0119(.A(G200), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n252), .A2(G50), .B1(G20), .B2(new_n246), .ZN(new_n321));
  INV_X1    g0121(.A(G77), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n321), .B1(new_n261), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n267), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT11), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n271), .B(G68), .C1(G1), .C2(new_n207), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n323), .A2(KEYINPUT11), .A3(new_n267), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n269), .A2(new_n246), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT12), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n320), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n312), .A2(new_n317), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT13), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n312), .A2(new_n313), .A3(new_n317), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(G190), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT69), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n336), .A2(KEYINPUT69), .A3(G190), .A4(new_n337), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n334), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n333), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT70), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n344), .B(G169), .C1(new_n318), .C2(new_n319), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT14), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(G169), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n336), .B2(new_n337), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n336), .A2(G179), .A3(new_n337), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n346), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n342), .B1(new_n343), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT15), .B(G87), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n261), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT8), .B(G58), .ZN(new_n356));
  INV_X1    g0156(.A(new_n252), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n356), .A2(new_n357), .B1(new_n217), .B2(new_n322), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n267), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n269), .A2(new_n322), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n359), .B(new_n360), .C1(new_n322), .C2(new_n272), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n286), .A2(G238), .A3(G1698), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n286), .A2(G232), .A3(new_n288), .ZN(new_n363));
  INV_X1    g0163(.A(G107), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n362), .B(new_n363), .C1(new_n364), .C2(new_n286), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n285), .ZN(new_n366));
  INV_X1    g0166(.A(new_n277), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n367), .A2(new_n280), .A3(G274), .ZN(new_n368));
  INV_X1    g0168(.A(G244), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n281), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n361), .B1(G200), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n370), .B1(new_n365), .B2(new_n285), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G190), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n372), .A2(new_n298), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n300), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(new_n361), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n297), .A2(new_n302), .A3(new_n353), .A4(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n286), .A2(G264), .A3(G1698), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n286), .A2(G257), .A3(new_n288), .ZN(new_n383));
  INV_X1    g0183(.A(G303), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n382), .B(new_n383), .C1(new_n384), .C2(new_n286), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n285), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n206), .A2(G45), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(KEYINPUT5), .B(G41), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n275), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n389), .A2(new_n388), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n275), .A2(new_n276), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n390), .A2(G270), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G200), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n293), .B2(new_n394), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n307), .A2(G1), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n267), .A2(new_n269), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G116), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT78), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G283), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n307), .A2(G97), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n217), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n400), .A2(G20), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n267), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT20), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n404), .A2(KEYINPUT20), .A3(new_n267), .A4(new_n405), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT78), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n398), .A2(new_n411), .A3(G116), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n269), .A2(new_n400), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n401), .A2(new_n410), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n396), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n298), .B1(new_n386), .B2(new_n393), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n416), .A2(KEYINPUT21), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n386), .A2(G179), .A3(new_n393), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n414), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n414), .A2(new_n416), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT21), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT79), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT79), .ZN(new_n424));
  AOI211_X1 g0224(.A(new_n424), .B(KEYINPUT21), .C1(new_n414), .C2(new_n416), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n415), .B(new_n420), .C1(new_n423), .C2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n217), .A2(new_n286), .A3(G87), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT22), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT22), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n217), .A2(new_n286), .A3(new_n429), .A4(G87), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n217), .A2(KEYINPUT23), .A3(G107), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT23), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(new_n364), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G116), .ZN(new_n435));
  AOI21_X1  g0235(.A(G20), .B1(new_n435), .B2(new_n433), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n432), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT24), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n431), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n438), .B1(new_n431), .B2(new_n437), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n267), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n306), .A2(new_n308), .A3(G257), .A4(G1698), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n306), .A2(new_n308), .A3(G250), .A4(new_n288), .ZN(new_n443));
  INV_X1    g0243(.A(G294), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n442), .B(new_n443), .C1(new_n307), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n285), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n391), .A2(new_n392), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n390), .A2(G264), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(G200), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n445), .A2(new_n285), .B1(new_n390), .B2(G264), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(new_n293), .A3(new_n447), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT25), .ZN(new_n455));
  INV_X1    g0255(.A(new_n269), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(G107), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n269), .A2(KEYINPUT25), .A3(new_n364), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n398), .A2(G107), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n441), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT80), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n441), .A2(new_n454), .A3(KEYINPUT80), .A4(new_n459), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n456), .A2(G97), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(new_n398), .B2(G97), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT7), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n286), .B2(G20), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT72), .B1(new_n307), .B2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT72), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(new_n305), .A3(G33), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n470), .A2(new_n472), .A3(new_n308), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n217), .A2(KEYINPUT7), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G107), .ZN(new_n476));
  XNOR2_X1  g0276(.A(G97), .B(G107), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT6), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n478), .A2(new_n310), .A3(G107), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT65), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G20), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n482), .A2(new_n486), .B1(G77), .B2(new_n252), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n476), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n467), .B1(new_n488), .B2(new_n267), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n306), .A2(new_n308), .A3(G244), .A4(new_n288), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n286), .A2(KEYINPUT4), .A3(G244), .A4(new_n288), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n286), .A2(G250), .A3(G1698), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n402), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n285), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n390), .A2(G257), .B1(new_n391), .B2(new_n392), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G200), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n496), .A2(G190), .A3(new_n497), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n489), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n298), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n470), .A2(new_n472), .A3(new_n308), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(KEYINPUT7), .A3(new_n217), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n364), .B1(new_n504), .B2(new_n469), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n480), .B1(new_n478), .B2(new_n477), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n506), .A2(new_n217), .B1(new_n322), .B2(new_n357), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n267), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n466), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n496), .A2(new_n300), .A3(new_n497), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n502), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n501), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n449), .A2(new_n298), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n452), .A2(new_n300), .A3(new_n447), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n515), .B1(new_n441), .B2(new_n459), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n388), .A2(new_n280), .A3(G274), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n280), .A2(G250), .A3(new_n387), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n286), .A2(G238), .A3(new_n288), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n306), .A2(new_n308), .A3(G244), .A4(G1698), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n435), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n520), .B1(new_n523), .B2(new_n285), .ZN(new_n524));
  OR2_X1    g0324(.A1(new_n524), .A2(G169), .ZN(new_n525));
  INV_X1    g0325(.A(new_n267), .ZN(new_n526));
  OR2_X1    g0326(.A1(KEYINPUT75), .A2(G87), .ZN(new_n527));
  NOR2_X1   g0327(.A1(G97), .A2(G107), .ZN(new_n528));
  NAND2_X1  g0328(.A1(KEYINPUT75), .A2(G87), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT19), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n531), .A2(new_n307), .A3(new_n310), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n532), .B2(new_n486), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n483), .A2(new_n485), .A3(G33), .A4(G97), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n531), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n217), .A2(new_n286), .A3(G68), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n526), .B1(new_n537), .B2(KEYINPUT76), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT76), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n533), .A2(new_n535), .A3(new_n539), .A4(new_n536), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n538), .A2(new_n540), .B1(new_n269), .B2(new_n354), .ZN(new_n541));
  INV_X1    g0341(.A(new_n354), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n398), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n543), .B(KEYINPUT77), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n541), .A2(new_n544), .B1(new_n300), .B2(new_n524), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n398), .A2(G87), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n524), .A2(new_n450), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(G190), .B2(new_n524), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n525), .A2(new_n545), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n464), .A2(new_n517), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT73), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n475), .A2(G68), .ZN(new_n553));
  INV_X1    g0353(.A(G159), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n357), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  XNOR2_X1  g0356(.A(KEYINPUT67), .B(G58), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n201), .B1(new_n557), .B2(G68), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n558), .B2(new_n207), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT16), .B1(new_n553), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(KEYINPUT16), .B(new_n556), .C1(new_n558), .C2(new_n207), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT71), .ZN(new_n563));
  AOI21_X1  g0363(.A(G20), .B1(new_n306), .B2(new_n308), .ZN(new_n564));
  OAI21_X1  g0364(.A(G68), .B1(new_n564), .B2(new_n468), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n483), .A2(new_n485), .A3(new_n468), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(new_n286), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n563), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT7), .B1(new_n286), .B2(G20), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n309), .A2(new_n217), .A3(new_n468), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT71), .A4(G68), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n562), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n561), .A2(new_n572), .A3(new_n526), .ZN(new_n573));
  INV_X1    g0373(.A(new_n260), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(new_n456), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n272), .B2(new_n260), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n552), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n562), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n305), .A2(G33), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n207), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n246), .B1(new_n582), .B2(KEYINPUT7), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT71), .B1(new_n583), .B2(new_n570), .ZN(new_n584));
  AND4_X1   g0384(.A1(KEYINPUT71), .A2(new_n569), .A3(new_n570), .A4(G68), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n579), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT16), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n246), .B1(new_n504), .B2(new_n469), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(new_n559), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n267), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n577), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(KEYINPUT73), .A3(new_n591), .ZN(new_n592));
  OR2_X1    g0392(.A1(G223), .A2(G1698), .ZN(new_n593));
  OR2_X1    g0393(.A1(new_n288), .A2(G226), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n286), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G87), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n284), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n368), .B1(new_n281), .B2(new_n233), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G179), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n298), .B2(new_n599), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n578), .A2(new_n592), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT18), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT74), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n568), .A2(new_n571), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n526), .B1(new_n605), .B2(new_n579), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n577), .B1(new_n606), .B2(new_n589), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n599), .A2(new_n293), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(G200), .B2(new_n599), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n604), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n604), .A2(new_n590), .A3(new_n591), .A4(new_n609), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT17), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT17), .B1(new_n607), .B2(new_n609), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT18), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n578), .A2(new_n615), .A3(new_n592), .A4(new_n601), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n603), .A2(new_n612), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  NOR4_X1   g0417(.A1(new_n381), .A2(new_n426), .A3(new_n551), .A4(new_n617), .ZN(G372));
  NOR2_X1   g0418(.A1(new_n381), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n441), .A2(new_n459), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n513), .A2(new_n514), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n420), .B(new_n622), .C1(new_n423), .C2(new_n425), .ZN(new_n623));
  INV_X1    g0423(.A(new_n512), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT81), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n523), .A2(new_n625), .A3(new_n285), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n625), .B1(new_n523), .B2(new_n285), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n518), .B(new_n519), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G200), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n524), .A2(G190), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n541), .A2(new_n546), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n628), .A2(new_n298), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n629), .A2(new_n631), .B1(new_n545), .B2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n623), .A2(new_n464), .A3(new_n624), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n545), .A2(new_n632), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  INV_X1    g0436(.A(new_n511), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n633), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n545), .A2(new_n525), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n547), .A2(new_n549), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(new_n640), .A3(new_n637), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT26), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n634), .A2(new_n635), .A3(new_n638), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n619), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n302), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n590), .A2(new_n591), .A3(new_n609), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT74), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n607), .A2(new_n604), .A3(new_n609), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n613), .B1(new_n649), .B2(KEYINPUT17), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n351), .B1(new_n348), .B2(new_n349), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n345), .A2(KEYINPUT14), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n343), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n379), .A2(KEYINPUT82), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT82), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n377), .A2(new_n655), .A3(new_n378), .A4(new_n361), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n653), .B1(new_n342), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n650), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n601), .B1(new_n573), .B2(new_n577), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(new_n615), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n645), .B1(new_n662), .B2(new_n297), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n644), .A2(new_n663), .ZN(G369));
  NAND3_X1  g0464(.A1(new_n217), .A2(new_n206), .A3(G13), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  OAI21_X1  g0466(.A(G213), .B1(new_n665), .B2(KEYINPUT27), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n414), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n426), .B2(KEYINPUT83), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(KEYINPUT83), .B2(new_n426), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n423), .A2(new_n425), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(new_n420), .A3(new_n671), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n622), .A2(new_n670), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n462), .A2(new_n463), .B1(new_n620), .B2(new_n670), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n516), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n674), .A2(new_n420), .ZN(new_n684));
  INV_X1    g0484(.A(new_n670), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n681), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n678), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n683), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n210), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT84), .ZN(new_n691));
  OR3_X1    g0491(.A1(new_n690), .A2(new_n691), .A3(G41), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n690), .B2(G41), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n530), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n220), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n643), .A2(new_n685), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(KEYINPUT29), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  INV_X1    g0501(.A(new_n633), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT26), .B1(new_n702), .B2(new_n511), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n550), .A2(new_n636), .A3(new_n637), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n703), .A2(new_n634), .A3(new_n635), .A4(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n701), .B1(new_n705), .B2(new_n685), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n700), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G330), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n496), .A2(new_n524), .A3(new_n452), .A4(new_n497), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(new_n418), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT85), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT85), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n713), .B(new_n709), .C1(new_n710), .C2(new_n418), .ZN(new_n714));
  OR3_X1    g0514(.A1(new_n710), .A2(new_n709), .A3(new_n418), .ZN(new_n715));
  AOI21_X1  g0515(.A(G179), .B1(new_n386), .B2(new_n393), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n628), .A2(new_n449), .A3(new_n498), .A4(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n712), .A2(new_n714), .A3(new_n715), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n670), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n715), .A2(new_n711), .A3(new_n717), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n464), .A2(new_n517), .ZN(new_n725));
  INV_X1    g0525(.A(new_n426), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n726), .A3(new_n550), .A4(new_n685), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n708), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n707), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n698), .B1(new_n731), .B2(G1), .ZN(G364));
  INV_X1    g0532(.A(new_n694), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n486), .A2(new_n268), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G45), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT86), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(KEYINPUT86), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(G1), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n677), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n676), .A2(G330), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n676), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n690), .A2(new_n286), .ZN(new_n749));
  INV_X1    g0549(.A(G45), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n221), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n749), .B(new_n751), .C1(new_n750), .C2(new_n250), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n690), .A2(new_n309), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n753), .A2(G355), .B1(new_n400), .B2(new_n690), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n755), .A2(KEYINPUT87), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n216), .B1(G20), .B2(new_n298), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n746), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(new_n755), .B2(KEYINPUT87), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n739), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n217), .A2(G190), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n762), .A2(new_n300), .A3(new_n450), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n217), .B1(G190), .B2(new_n765), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n764), .A2(new_n246), .B1(new_n766), .B2(new_n310), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n527), .A2(new_n529), .ZN(new_n768));
  NOR4_X1   g0568(.A1(new_n207), .A2(new_n293), .A3(new_n450), .A4(G179), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n769), .A2(KEYINPUT90), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(KEYINPUT90), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n309), .B(new_n767), .C1(new_n768), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n217), .A2(new_n300), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G190), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n450), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n776), .A2(G200), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n774), .B1(new_n202), .B2(new_n778), .C1(new_n258), .C2(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n762), .A2(G179), .A3(new_n450), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n782), .A2(KEYINPUT91), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(KEYINPUT91), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G107), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n761), .A2(new_n765), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n554), .ZN(new_n789));
  XNOR2_X1  g0589(.A(KEYINPUT89), .B(KEYINPUT32), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n775), .A2(new_n293), .A3(new_n450), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n793), .A2(KEYINPUT88), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(KEYINPUT88), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n787), .B(new_n791), .C1(new_n322), .C2(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n777), .B(KEYINPUT92), .Z(new_n798));
  INV_X1    g0598(.A(G326), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G311), .ZN(new_n801));
  INV_X1    g0601(.A(G329), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n792), .A2(new_n801), .B1(new_n788), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n772), .A2(new_n384), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT33), .B(G317), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n803), .B(new_n804), .C1(new_n763), .C2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n309), .B1(new_n766), .B2(new_n444), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(new_n779), .B2(G322), .ZN(new_n808));
  INV_X1    g0608(.A(G283), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n806), .B(new_n808), .C1(new_n809), .C2(new_n785), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n781), .A2(new_n797), .B1(new_n800), .B2(new_n810), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT93), .Z(new_n812));
  AOI21_X1  g0612(.A(new_n760), .B1(new_n812), .B2(new_n757), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n743), .B1(new_n748), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NAND4_X1  g0615(.A1(new_n654), .A2(new_n361), .A3(new_n656), .A4(new_n670), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n670), .A2(new_n361), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n376), .A2(new_n379), .A3(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n699), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n819), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n643), .A2(new_n685), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n739), .B1(new_n823), .B2(new_n729), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n729), .B2(new_n823), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n757), .A2(new_n744), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n739), .B1(G77), .B2(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT94), .Z(new_n829));
  OAI221_X1 g0629(.A(new_n309), .B1(new_n766), .B2(new_n310), .C1(new_n780), .C2(new_n444), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G303), .B2(new_n777), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n786), .A2(G87), .ZN(new_n832));
  INV_X1    g0632(.A(new_n796), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G116), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n764), .A2(new_n809), .B1(new_n801), .B2(new_n788), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G107), .B2(new_n773), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n831), .A2(new_n832), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n779), .A2(G143), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  INV_X1    g0639(.A(G150), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n838), .B1(new_n778), .B2(new_n839), .C1(new_n840), .C2(new_n764), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G159), .B2(new_n833), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT34), .ZN(new_n843));
  INV_X1    g0643(.A(new_n788), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n309), .B1(new_n844), .B2(G132), .ZN(new_n845));
  INV_X1    g0645(.A(new_n766), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n773), .A2(G50), .B1(new_n557), .B2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n845), .B(new_n847), .C1(new_n785), .C2(new_n246), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n837), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n829), .B1(new_n849), .B2(new_n757), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n745), .B2(new_n821), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n825), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G384));
  OR2_X1    g0653(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(G116), .A3(new_n218), .A4(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT36), .Z(new_n857));
  OAI211_X1 g0657(.A(new_n221), .B(G77), .C1(new_n246), .C2(new_n258), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n206), .B(G13), .C1(new_n858), .C2(new_n245), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n668), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n661), .A2(new_n861), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n379), .A2(new_n670), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n822), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n340), .A2(new_n341), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(new_n333), .A3(new_n320), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n343), .A2(new_n670), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n653), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n343), .B(new_n670), .C1(new_n342), .C2(new_n352), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n610), .A2(new_n611), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n578), .B(new_n592), .C1(new_n601), .C2(new_n861), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n559), .B1(new_n568), .B2(new_n571), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n606), .B1(KEYINPUT16), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n601), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n878), .A2(new_n591), .B1(new_n879), .B2(new_n668), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT37), .B1(new_n649), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n668), .B1(new_n878), .B2(new_n591), .ZN(new_n882));
  AOI221_X4 g0682(.A(new_n872), .B1(new_n876), .B2(new_n881), .C1(new_n617), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n617), .A2(new_n882), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n876), .A2(new_n881), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n862), .B1(new_n871), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT95), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(KEYINPUT95), .B(new_n862), .C1(new_n871), .C2(new_n887), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT39), .ZN(new_n892));
  INV_X1    g0692(.A(new_n874), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n647), .A2(new_n648), .A3(new_n875), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT96), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT96), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n873), .A2(new_n874), .A3(new_n896), .A4(new_n875), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n578), .A2(new_n592), .A3(new_n861), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(new_n646), .A3(new_n660), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT37), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n895), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n650), .A2(new_n661), .ZN(new_n902));
  INV_X1    g0702(.A(new_n898), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n892), .B1(new_n905), .B2(new_n883), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n352), .A2(new_n343), .A3(new_n685), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n884), .A2(new_n885), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n872), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n884), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(KEYINPUT39), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n906), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n890), .A2(new_n891), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n619), .B1(new_n700), .B2(new_n706), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n663), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n914), .B(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n721), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n727), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n819), .B1(new_n868), .B2(new_n869), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n921), .B(new_n922), .C1(new_n883), .C2(new_n886), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT40), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n876), .A2(KEYINPUT96), .B1(new_n899), .B2(KEYINPUT37), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n925), .A2(new_n897), .B1(new_n903), .B2(new_n902), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n911), .B1(new_n926), .B2(KEYINPUT38), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n551), .A2(new_n426), .A3(new_n670), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n922), .B(KEYINPUT40), .C1(new_n928), .C2(new_n919), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n923), .A2(new_n924), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(new_n619), .A3(new_n921), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(G330), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n931), .B1(new_n619), .B2(new_n921), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n917), .A2(new_n935), .B1(new_n206), .B2(new_n734), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT97), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n917), .A2(new_n935), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n936), .A2(KEYINPUT97), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n860), .B1(new_n939), .B2(new_n940), .ZN(G367));
  INV_X1    g0741(.A(new_n749), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n240), .A2(new_n942), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n746), .B(new_n757), .C1(new_n690), .C2(new_n542), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n740), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT104), .Z(new_n946));
  OAI21_X1  g0746(.A(new_n633), .B1(new_n547), .B2(new_n685), .ZN(new_n947));
  OR3_X1    g0747(.A1(new_n635), .A2(new_n547), .A3(new_n685), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n773), .A2(KEYINPUT46), .A3(G116), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT46), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n772), .B2(new_n400), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n950), .B(new_n952), .C1(new_n384), .C2(new_n780), .ZN(new_n953));
  INV_X1    g0753(.A(G317), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n788), .A2(new_n954), .B1(new_n766), .B2(new_n364), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n286), .B(new_n955), .C1(G294), .C2(new_n763), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n956), .B1(new_n796), .B2(new_n809), .C1(new_n310), .C2(new_n785), .ZN(new_n957));
  INV_X1    g0757(.A(new_n798), .ZN(new_n958));
  XNOR2_X1  g0758(.A(KEYINPUT105), .B(G311), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n953), .B(new_n957), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT106), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n763), .A2(G159), .B1(G137), .B2(new_n844), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n962), .B(new_n286), .C1(new_n258), .C2(new_n772), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n785), .A2(new_n322), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(G50), .C2(new_n833), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n846), .A2(G68), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n780), .B2(new_n840), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(KEYINPUT107), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(KEYINPUT107), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n968), .B(new_n969), .C1(G143), .C2(new_n958), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n961), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n972));
  AND2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n757), .B1(new_n971), .B2(new_n972), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n946), .B1(new_n747), .B2(new_n949), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n624), .B1(new_n489), .B2(new_n685), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n637), .A2(new_n670), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n687), .A2(new_n678), .A3(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT45), .Z(new_n981));
  NOR2_X1   g0781(.A1(new_n688), .A2(new_n978), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(KEYINPUT101), .ZN(new_n983));
  XNOR2_X1  g0783(.A(KEYINPUT100), .B(KEYINPUT44), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n981), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n983), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n982), .A2(KEYINPUT101), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n987), .A2(new_n988), .A3(new_n984), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n682), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n986), .A2(new_n989), .A3(new_n683), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT103), .B1(new_n676), .B2(G330), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT102), .B1(new_n686), .B2(new_n681), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(new_n687), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n687), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n999), .A2(new_n730), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n993), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n731), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n694), .B(KEYINPUT41), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n738), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n687), .A2(new_n978), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(KEYINPUT99), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(KEYINPUT99), .ZN(new_n1010));
  AOI21_X1  g0810(.A(KEYINPUT42), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1009), .A2(KEYINPUT42), .A3(new_n1010), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n511), .B1(new_n976), .B2(new_n622), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1012), .A2(new_n1013), .B1(new_n685), .B2(new_n1014), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n949), .A2(KEYINPUT98), .ZN(new_n1016));
  AOI21_X1  g0816(.A(KEYINPUT43), .B1(new_n949), .B2(KEYINPUT98), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n1016), .A2(new_n1017), .B1(KEYINPUT43), .B2(new_n949), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n683), .A2(new_n979), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1021), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n975), .B1(new_n1005), .B2(new_n1027), .ZN(G387));
  INV_X1    g0828(.A(new_n1000), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n999), .A2(new_n730), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1029), .A2(new_n733), .A3(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n236), .A2(new_n750), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n695), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n1032), .A2(new_n749), .B1(new_n1033), .B2(new_n753), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT50), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n356), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1035), .B1(new_n1036), .B2(new_n202), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n750), .B1(new_n246), .B2(new_n322), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n356), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1039));
  NOR4_X1   g0839(.A1(new_n1033), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1034), .A2(new_n1040), .B1(G107), .B2(new_n210), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n740), .B1(new_n1041), .B2(new_n758), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n309), .B1(new_n773), .B2(G77), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n202), .B2(new_n780), .C1(new_n554), .C2(new_n778), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n785), .A2(new_n310), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n764), .A2(new_n260), .B1(new_n354), .B2(new_n766), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n792), .A2(new_n246), .B1(new_n788), .B2(new_n840), .ZN(new_n1047));
  NOR4_X1   g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n309), .B1(new_n788), .B2(new_n799), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n763), .A2(new_n959), .B1(new_n779), .B2(G317), .ZN(new_n1050));
  INV_X1    g0850(.A(G322), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1050), .B1(new_n796), .B2(new_n384), .C1(new_n798), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT48), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n773), .A2(G294), .B1(G283), .B2(new_n846), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT49), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1049), .B(new_n1059), .C1(G116), .C2(new_n786), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1048), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n757), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1042), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n681), .B2(new_n746), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n999), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1065), .B1(new_n1066), .B2(new_n738), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1031), .A2(new_n1067), .ZN(G393));
  NAND2_X1  g0868(.A1(new_n993), .A2(new_n738), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n758), .B1(new_n310), .B2(new_n210), .C1(new_n942), .C2(new_n244), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT109), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n739), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G150), .A2(new_n777), .B1(new_n779), .B2(G159), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT51), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n309), .B1(new_n844), .B2(G143), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n772), .A2(new_n246), .B1(new_n322), .B2(new_n766), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G50), .B2(new_n763), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n833), .A2(new_n1036), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n832), .A2(new_n1077), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n286), .B1(new_n844), .B2(G322), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n773), .A2(G283), .B1(G303), .B2(new_n763), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n793), .A2(G294), .B1(G116), .B2(new_n846), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n787), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G311), .A2(new_n779), .B1(new_n777), .B2(G317), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT52), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n1076), .A2(new_n1081), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1072), .B(new_n1074), .C1(new_n1088), .C2(new_n757), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n747), .B2(new_n978), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1069), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1001), .A2(new_n733), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n993), .A2(new_n1000), .ZN(new_n1093));
  OAI21_X1  g0893(.A(KEYINPUT110), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1093), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT110), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1095), .A2(new_n1096), .A3(new_n1001), .A4(new_n733), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1091), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(G390));
  AOI21_X1  g0899(.A(new_n708), .B1(new_n920), .B2(new_n727), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n922), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n906), .A2(new_n912), .B1(new_n871), .B2(new_n907), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n705), .A2(new_n685), .A3(new_n821), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n863), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n870), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1106), .A2(new_n927), .A3(new_n907), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1102), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n906), .A2(new_n912), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n871), .A2(new_n907), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1106), .A2(new_n927), .A3(new_n907), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n728), .A2(new_n821), .A3(new_n870), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1108), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1100), .A2(new_n619), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n915), .A2(new_n663), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1100), .A2(new_n821), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n868), .A3(new_n869), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1119), .A2(new_n863), .A3(new_n1104), .A4(new_n1113), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n870), .B1(new_n728), .B2(new_n821), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n864), .B1(new_n1102), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1117), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n694), .B1(new_n1115), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1108), .A2(new_n1114), .A3(new_n1123), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1109), .A2(new_n744), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n286), .B1(new_n773), .B2(G87), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n809), .B2(new_n778), .C1(new_n444), .C2(new_n788), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G68), .B2(new_n786), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n796), .A2(new_n310), .B1(new_n364), .B2(new_n764), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1132), .A2(KEYINPUT111), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(KEYINPUT111), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n779), .A2(G116), .B1(G77), .B2(new_n846), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT112), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1131), .A2(new_n1133), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n786), .A2(G50), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G128), .A2(new_n777), .B1(new_n779), .B2(G132), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n309), .B1(new_n846), .B2(G159), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n763), .A2(G137), .B1(G125), .B2(new_n844), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT54), .B(G143), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n833), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n772), .A2(new_n840), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT53), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1138), .A2(new_n1142), .A3(new_n1145), .A4(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1063), .B1(new_n1137), .B2(new_n1148), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n740), .B(new_n1149), .C1(new_n260), .C2(new_n826), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1128), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n738), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1151), .B1(new_n1115), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1127), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(G378));
  INV_X1    g0955(.A(new_n1117), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1126), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n930), .B1(new_n905), .B2(new_n883), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n922), .B1(new_n928), .B2(new_n919), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n910), .B2(new_n911), .ZN(new_n1160));
  OAI211_X1 g0960(.A(G330), .B(new_n1158), .C1(new_n1160), .C2(KEYINPUT40), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n297), .A2(new_n302), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n273), .A2(new_n861), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1164), .B(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1161), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT114), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1161), .A2(new_n1167), .A3(KEYINPUT114), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n914), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT115), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n1161), .B2(new_n1167), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1164), .B(new_n1165), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n931), .A2(new_n1176), .A3(KEYINPUT115), .A4(G330), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1172), .A2(new_n1173), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1173), .B1(new_n1172), .B2(new_n1178), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1157), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT57), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1182), .B1(new_n1126), .B2(new_n1156), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT116), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(KEYINPUT116), .B(new_n1184), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1183), .A2(new_n1187), .A3(new_n733), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1172), .A2(new_n1178), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n914), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1172), .A2(new_n1173), .A3(new_n1178), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1167), .A2(new_n744), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n739), .B1(G50), .B2(new_n827), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT113), .Z(new_n1196));
  AOI22_X1  g0996(.A1(new_n773), .A2(G77), .B1(G97), .B2(new_n763), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n793), .A2(new_n542), .B1(new_n844), .B2(G283), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n785), .A2(new_n258), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n286), .A2(G41), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n846), .B2(G68), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n778), .B2(new_n400), .C1(new_n364), .C2(new_n780), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1199), .A2(new_n1200), .A3(new_n1204), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1205), .A2(KEYINPUT58), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n773), .A2(new_n1144), .B1(G132), .B2(new_n763), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n793), .A2(G137), .B1(G150), .B2(new_n846), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G125), .A2(new_n777), .B1(new_n779), .B2(G128), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n786), .A2(G159), .ZN(new_n1213));
  AOI211_X1 g1013(.A(G33), .B(G41), .C1(new_n844), .C2(G124), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1205), .A2(KEYINPUT58), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1202), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1206), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1196), .B1(new_n1218), .B2(new_n757), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1193), .A2(new_n738), .B1(new_n1194), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1189), .A2(new_n1220), .ZN(G375));
  AOI21_X1  g1021(.A(new_n740), .B1(new_n246), .B2(new_n826), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n773), .A2(G97), .B1(G303), .B2(new_n844), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n286), .B1(new_n846), .B2(new_n542), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G283), .A2(new_n779), .B1(new_n777), .B2(G294), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n796), .A2(new_n364), .B1(new_n400), .B2(new_n764), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1226), .B(new_n964), .C1(KEYINPUT117), .C2(new_n1227), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1227), .A2(KEYINPUT117), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n309), .B1(new_n844), .B2(G128), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n780), .B2(new_n839), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G132), .B2(new_n777), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n792), .A2(new_n840), .B1(new_n202), .B2(new_n766), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n764), .A2(new_n1143), .B1(new_n554), .B2(new_n772), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1200), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1228), .A2(new_n1229), .B1(new_n1232), .B2(new_n1235), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1222), .B1(new_n1236), .B2(new_n1063), .C1(new_n870), .C2(new_n745), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1237), .B1(new_n1238), .B2(new_n1152), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT118), .Z(new_n1240));
  NAND3_X1  g1040(.A1(new_n1120), .A2(new_n1117), .A3(new_n1122), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1124), .A2(new_n1004), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1240), .A2(new_n1242), .ZN(G381));
  NAND3_X1  g1043(.A1(new_n1031), .A2(new_n814), .A3(new_n1067), .ZN(new_n1244));
  NOR4_X1   g1044(.A1(G387), .A2(G384), .A3(G381), .A4(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(G375), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1245), .A2(new_n1098), .A3(new_n1154), .A4(new_n1246), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT119), .ZN(G407));
  NAND2_X1  g1048(.A1(new_n669), .A2(G213), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1249), .B(KEYINPUT120), .Z(new_n1250));
  NAND3_X1  g1050(.A1(new_n1246), .A2(new_n1154), .A3(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(G407), .A2(G213), .A3(new_n1251), .ZN(G409));
  INV_X1    g1052(.A(KEYINPUT127), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1004), .B(new_n1157), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT122), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1193), .A2(KEYINPUT122), .A3(new_n1004), .A4(new_n1157), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1220), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1154), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1126), .A2(new_n1156), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n733), .B1(new_n1263), .B2(KEYINPUT57), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G378), .B(new_n1220), .C1(new_n1261), .C2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT121), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1189), .A2(KEYINPUT121), .A3(G378), .A4(new_n1220), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1260), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1269), .A2(new_n1250), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1241), .A2(KEYINPUT124), .ZN(new_n1271));
  XOR2_X1   g1071(.A(new_n1271), .B(KEYINPUT60), .Z(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(new_n733), .A3(new_n1124), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1240), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n852), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1273), .A2(G384), .A3(new_n1240), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1270), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1259), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT123), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1250), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT123), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1269), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1277), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1283), .A2(new_n1284), .A3(new_n1286), .A4(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1280), .B1(new_n1288), .B2(new_n1278), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1250), .A2(G2897), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1277), .B(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1270), .A2(new_n1292), .ZN(new_n1293));
  OR2_X1    g1093(.A1(new_n1293), .A2(KEYINPUT61), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1253), .B1(new_n1289), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1270), .A2(new_n1279), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1284), .B1(new_n1269), .B2(new_n1285), .ZN(new_n1297));
  AOI211_X1 g1097(.A(KEYINPUT123), .B(new_n1260), .C1(new_n1267), .C2(new_n1268), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n1277), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1296), .B1(new_n1299), .B2(KEYINPUT62), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1293), .A2(KEYINPUT61), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(KEYINPUT127), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1098), .A2(G387), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1098), .A2(G387), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT126), .B1(new_n1098), .B2(G387), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G393), .A2(G396), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1244), .ZN(new_n1308));
  OAI22_X1  g1108(.A1(new_n1304), .A2(new_n1305), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1309));
  OR2_X1    g1109(.A1(new_n1098), .A2(G387), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1308), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1310), .A2(KEYINPUT126), .A3(new_n1311), .A4(new_n1303), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1309), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1295), .A2(new_n1302), .A3(new_n1313), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1270), .A2(KEYINPUT63), .A3(new_n1287), .ZN(new_n1315));
  NOR3_X1   g1115(.A1(new_n1315), .A2(KEYINPUT61), .A3(new_n1313), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1283), .A2(new_n1284), .A3(new_n1286), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1317), .A2(KEYINPUT125), .A3(new_n1291), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT125), .B1(new_n1317), .B2(new_n1291), .ZN(new_n1320));
  OAI221_X1 g1120(.A(new_n1316), .B1(KEYINPUT63), .B2(new_n1299), .C1(new_n1319), .C2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1314), .A2(new_n1321), .ZN(G405));
  OAI21_X1  g1122(.A(new_n1281), .B1(G378), .B2(new_n1246), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(new_n1323), .B(new_n1287), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1324), .B(new_n1313), .ZN(G402));
endmodule


