//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944;
  INV_X1    g000(.A(KEYINPUT34), .ZN(new_n202));
  INV_X1    g001(.A(G227gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(KEYINPUT72), .A2(G134gat), .ZN(new_n207));
  INV_X1    g006(.A(G120gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G113gat), .ZN(new_n209));
  INV_X1    g008(.A(G113gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G120gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n207), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI211_X1 g013(.A(KEYINPUT1), .B(G134gat), .C1(new_n209), .C2(new_n211), .ZN(new_n215));
  NOR3_X1   g014(.A1(new_n214), .A2(new_n215), .A3(G127gat), .ZN(new_n216));
  INV_X1    g015(.A(G127gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(G113gat), .B(G120gat), .ZN(new_n218));
  OAI211_X1 g017(.A(KEYINPUT72), .B(G134gat), .C1(new_n218), .C2(KEYINPUT1), .ZN(new_n219));
  INV_X1    g018(.A(G134gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n212), .A2(new_n213), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n217), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  OR3_X1    g022(.A1(KEYINPUT71), .A2(G169gat), .A3(G176gat), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n224), .A2(KEYINPUT26), .ZN(new_n225));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n224), .A2(KEYINPUT26), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n225), .A2(new_n230), .B1(G183gat), .B2(G190gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT68), .ZN(new_n232));
  INV_X1    g031(.A(G183gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(G190gat), .B1(new_n236), .B2(KEYINPUT27), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT27), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n233), .B1(KEYINPUT70), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(KEYINPUT70), .B2(new_n238), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT28), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT27), .B(G183gat), .Z(new_n242));
  INV_X1    g041(.A(KEYINPUT28), .ZN(new_n243));
  NOR3_X1   g042(.A1(new_n242), .A2(new_n243), .A3(G190gat), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n231), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G190gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n234), .A2(new_n246), .A3(new_n235), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(KEYINPUT67), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n247), .A2(new_n249), .A3(new_n252), .A4(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT23), .ZN(new_n256));
  INV_X1    g055(.A(G169gat), .ZN(new_n257));
  INV_X1    g056(.A(G176gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n255), .A2(new_n259), .B1(new_n228), .B2(new_n229), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n254), .A2(KEYINPUT25), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n254), .A2(KEYINPUT69), .A3(new_n260), .A4(KEYINPUT25), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n259), .A2(new_n255), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n228), .A2(new_n229), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n250), .A2(KEYINPUT64), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n270), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n248), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n268), .B1(new_n275), .B2(KEYINPUT65), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT65), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n272), .A2(new_n277), .A3(new_n274), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT25), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n223), .B(new_n245), .C1(new_n265), .C2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n272), .A2(new_n277), .A3(new_n274), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n277), .B1(new_n272), .B2(new_n274), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n282), .A2(new_n283), .A3(new_n268), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n263), .B(new_n264), .C1(new_n284), .C2(KEYINPUT25), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n223), .B1(new_n285), .B2(new_n245), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n202), .B(new_n206), .C1(new_n281), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT75), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n281), .A2(new_n286), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT34), .B1(new_n289), .B2(new_n205), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n245), .B1(new_n265), .B2(new_n279), .ZN(new_n291));
  OAI21_X1  g090(.A(G127gat), .B1(new_n214), .B2(new_n215), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n219), .A2(new_n217), .A3(new_n221), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n280), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n296), .A2(new_n297), .A3(new_n202), .A4(new_n206), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n288), .A2(new_n290), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G15gat), .B(G43gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(G71gat), .B(G99gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT33), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(KEYINPUT73), .ZN(new_n305));
  OAI211_X1 g104(.A(KEYINPUT32), .B(new_n305), .C1(new_n296), .C2(new_n206), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n295), .A2(new_n205), .A3(new_n280), .A4(new_n303), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT73), .B1(new_n307), .B2(new_n304), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(new_n289), .B2(new_n205), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n306), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n299), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n299), .A2(new_n311), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT36), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n288), .A2(new_n290), .A3(new_n298), .ZN(new_n319));
  OAI211_X1 g118(.A(KEYINPUT74), .B(new_n306), .C1(new_n308), .C2(new_n310), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(KEYINPUT36), .A3(new_n313), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G228gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(new_n204), .ZN(new_n325));
  OR3_X1    g124(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n326));
  INV_X1    g125(.A(G155gat), .ZN(new_n327));
  INV_X1    g126(.A(G162gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT82), .ZN(new_n330));
  INV_X1    g129(.A(G141gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n330), .B1(new_n331), .B2(G148gat), .ZN(new_n332));
  INV_X1    g131(.A(G148gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n333), .A2(KEYINPUT82), .A3(G141gat), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n332), .B(new_n334), .C1(G141gat), .C2(new_n333), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  OR2_X1    g135(.A1(KEYINPUT80), .A2(KEYINPUT2), .ZN(new_n337));
  NAND2_X1  g136(.A1(KEYINPUT80), .A2(KEYINPUT2), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n331), .A2(G148gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n333), .A2(G141gat), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n337), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT81), .ZN(new_n342));
  XOR2_X1   g141(.A(G155gat), .B(G162gat), .Z(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n342), .B1(new_n341), .B2(new_n343), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n336), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G197gat), .B(G204gat), .ZN(new_n348));
  INV_X1    g147(.A(G218gat), .ZN(new_n349));
  OR2_X1    g148(.A1(KEYINPUT76), .A2(G211gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(KEYINPUT76), .A2(G211gat), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n348), .B1(new_n352), .B2(KEYINPUT22), .ZN(new_n353));
  XNOR2_X1  g152(.A(G211gat), .B(G218gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n348), .B(new_n354), .C1(new_n352), .C2(KEYINPUT22), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT29), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n347), .B1(new_n358), .B2(KEYINPUT3), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n360), .B(new_n336), .C1(new_n345), .C2(new_n346), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT77), .ZN(new_n363));
  INV_X1    g162(.A(new_n357), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT22), .ZN(new_n365));
  AND2_X1   g164(.A1(KEYINPUT76), .A2(G211gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(KEYINPUT76), .A2(G211gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n365), .B1(new_n368), .B2(new_n349), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n354), .B1(new_n369), .B2(new_n348), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n363), .B1(new_n364), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT77), .A3(new_n357), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n361), .A2(new_n362), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT91), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n359), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n361), .A2(new_n362), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n371), .A2(new_n372), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(KEYINPUT91), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n325), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n356), .A2(new_n357), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n325), .B1(new_n383), .B2(KEYINPUT90), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT89), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n347), .B(new_n385), .C1(new_n358), .C2(KEYINPUT3), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n381), .B1(new_n361), .B2(new_n362), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT90), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n387), .A2(new_n388), .B1(new_n359), .B2(KEYINPUT89), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT31), .B(G50gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n380), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n392), .B1(new_n380), .B2(new_n390), .ZN(new_n394));
  XNOR2_X1  g193(.A(G78gat), .B(G106gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(G22gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n325), .ZN(new_n399));
  INV_X1    g198(.A(new_n359), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n400), .B1(new_n378), .B2(KEYINPUT91), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n373), .A2(new_n374), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n359), .A2(KEYINPUT89), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n404), .B(new_n386), .C1(new_n383), .C2(KEYINPUT90), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n399), .B1(new_n387), .B2(new_n388), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n391), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n380), .A2(new_n390), .A3(new_n392), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n396), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n398), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(G226gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n412), .A2(new_n204), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n291), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT78), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n291), .A2(KEYINPUT78), .A3(new_n413), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n413), .B1(new_n291), .B2(new_n362), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n377), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n414), .A3(new_n381), .ZN(new_n423));
  XOR2_X1   g222(.A(G8gat), .B(G36gat), .Z(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(KEYINPUT79), .ZN(new_n425));
  XNOR2_X1  g224(.A(G64gat), .B(G92gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n422), .A2(KEYINPUT30), .A3(new_n423), .A4(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n419), .B1(new_n416), .B2(new_n417), .ZN(new_n430));
  INV_X1    g229(.A(new_n377), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n423), .B(new_n428), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT30), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n423), .B1(new_n430), .B2(new_n431), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n427), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n429), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(G1gat), .B(G29gat), .Z(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G57gat), .B(G85gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  XOR2_X1   g242(.A(KEYINPUT85), .B(KEYINPUT5), .Z(new_n444));
  NAND3_X1  g243(.A1(new_n292), .A2(KEYINPUT83), .A3(new_n293), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT83), .B1(new_n292), .B2(new_n293), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n347), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT84), .B1(new_n223), .B2(new_n347), .ZN(new_n449));
  INV_X1    g248(.A(new_n346), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n450), .A2(new_n344), .B1(new_n329), .B2(new_n335), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT84), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n294), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n448), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(G225gat), .A2(G233gat), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n444), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT4), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n449), .A2(new_n453), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n460), .B1(new_n216), .B2(new_n222), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n445), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n347), .A2(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n361), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n451), .A2(KEYINPUT4), .A3(new_n294), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n459), .A2(new_n455), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n457), .A2(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n464), .A2(new_n455), .A3(new_n444), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT4), .B1(new_n451), .B2(new_n294), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n449), .A2(new_n453), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n469), .B1(new_n470), .B2(KEYINPUT4), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n443), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT88), .B1(new_n473), .B2(KEYINPUT6), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n457), .A2(new_n466), .B1(new_n468), .B2(new_n471), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT88), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477));
  NOR4_X1   g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .A4(new_n443), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n473), .A2(KEYINPUT87), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT6), .B1(new_n475), .B2(new_n443), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT87), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n475), .B2(new_n443), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n437), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n323), .B1(new_n411), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n419), .B1(new_n413), .B2(new_n291), .ZN(new_n487));
  OAI22_X1  g286(.A1(new_n421), .A2(new_n377), .B1(new_n381), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT38), .B1(new_n488), .B2(KEYINPUT37), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n435), .A2(KEYINPUT37), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n427), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n473), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n481), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n491), .A2(new_n479), .A3(new_n432), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n435), .A2(KEYINPUT37), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n490), .A2(new_n495), .A3(new_n427), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT92), .B1(new_n496), .B2(KEYINPUT38), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(KEYINPUT92), .A3(KEYINPUT38), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n411), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n471), .A2(new_n464), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n456), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n503), .A2(KEYINPUT39), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n503), .B(KEYINPUT39), .C1(new_n456), .C2(new_n454), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(new_n443), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT40), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n473), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT40), .A4(new_n443), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n501), .B1(new_n510), .B2(new_n437), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n486), .B1(new_n500), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT93), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n397), .B1(new_n393), .B2(new_n394), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n408), .A2(new_n396), .A3(new_n409), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n313), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n513), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n411), .A2(new_n321), .A3(KEYINPUT93), .A4(new_n313), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n485), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT35), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT94), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(KEYINPUT94), .A3(KEYINPUT35), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n501), .A2(new_n314), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT35), .B1(new_n479), .B2(new_n493), .ZN(new_n527));
  INV_X1    g326(.A(new_n437), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n512), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(G197gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT11), .B(G169gat), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n532), .B(new_n533), .Z(new_n534));
  XOR2_X1   g333(.A(new_n534), .B(KEYINPUT12), .Z(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT99), .ZN(new_n537));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT16), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT98), .B1(new_n539), .B2(G1gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n539), .A2(KEYINPUT98), .A3(G1gat), .ZN(new_n542));
  OAI221_X1 g341(.A(new_n537), .B1(G1gat), .B2(new_n538), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n543), .B(G8gat), .Z(new_n544));
  XNOR2_X1  g343(.A(G43gat), .B(G50gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT15), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT14), .ZN(new_n547));
  OR3_X1    g346(.A1(new_n547), .A2(G29gat), .A3(G36gat), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(G29gat), .B2(G36gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT95), .B(G29gat), .ZN(new_n550));
  INV_X1    g349(.A(G36gat), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n548), .B(new_n549), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  OR3_X1    g351(.A1(new_n546), .A2(KEYINPUT96), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(KEYINPUT15), .A3(new_n545), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n554), .B(KEYINPUT96), .C1(new_n552), .C2(new_n546), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n544), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n553), .A2(new_n555), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT97), .B(KEYINPUT17), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n544), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n556), .A2(KEYINPUT17), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n557), .B1(new_n563), .B2(KEYINPUT100), .ZN(new_n564));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT100), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n561), .B2(new_n562), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT18), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n544), .B(new_n556), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n565), .B(KEYINPUT13), .Z(new_n572));
  AOI22_X1  g371(.A1(new_n568), .A2(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n536), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n570), .A2(new_n573), .A3(new_n536), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n530), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G57gat), .B(G64gat), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G71gat), .B(G78gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(G127gat), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n544), .B1(new_n585), .B2(new_n584), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(new_n327), .ZN(new_n593));
  XOR2_X1   g392(.A(G183gat), .B(G211gat), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n591), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AND2_X1   g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT41), .ZN(new_n602));
  NAND2_X1  g401(.A1(G99gat), .A2(G106gat), .ZN(new_n603));
  INV_X1    g402(.A(G85gat), .ZN(new_n604));
  INV_X1    g403(.A(G92gat), .ZN(new_n605));
  AOI22_X1  g404(.A1(KEYINPUT8), .A2(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT103), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G85gat), .A2(G92gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G99gat), .B(G106gat), .Z(new_n613));
  OR2_X1    g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n560), .A2(new_n616), .ZN(new_n617));
  OAI221_X1 g416(.A(new_n602), .B1(new_n556), .B2(new_n616), .C1(new_n617), .C2(new_n562), .ZN(new_n618));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n618), .B(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n601), .A2(KEYINPUT41), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT101), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n622), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n600), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT106), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n584), .B1(new_n614), .B2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(new_n616), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G120gat), .B(G148gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT108), .ZN(new_n638));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n616), .A2(new_n642), .A3(new_n584), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT107), .B(KEYINPUT10), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n634), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n635), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n636), .B(new_n641), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT109), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n645), .A2(new_n646), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n636), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n640), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n631), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n579), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n479), .A2(new_n484), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT110), .B(G1gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(G1324gat));
  NAND3_X1  g461(.A1(new_n579), .A2(new_n437), .A3(new_n657), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n663), .A2(G8gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT16), .B(G8gat), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT42), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(KEYINPUT42), .B2(new_n666), .ZN(G1325gat));
  OAI21_X1  g467(.A(G15gat), .B1(new_n658), .B2(new_n323), .ZN(new_n669));
  INV_X1    g468(.A(new_n579), .ZN(new_n670));
  OR3_X1    g469(.A1(new_n656), .A2(G15gat), .A3(new_n314), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(G1326gat));
  NOR2_X1   g471(.A1(new_n658), .A2(new_n411), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT43), .B(G22gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  INV_X1    g474(.A(new_n630), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n676), .A2(new_n654), .A3(new_n599), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n579), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n659), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n550), .ZN(new_n680));
  OR3_X1    g479(.A1(new_n678), .A2(KEYINPUT111), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT111), .B1(new_n678), .B2(new_n680), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n681), .A2(KEYINPUT45), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT45), .B1(new_n681), .B2(new_n682), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n599), .B(KEYINPUT112), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(new_n577), .A3(new_n655), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT113), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n520), .A2(KEYINPUT94), .A3(KEYINPUT35), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT94), .B1(new_n520), .B2(KEYINPUT35), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n529), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n500), .A2(new_n511), .ZN(new_n692));
  INV_X1    g491(.A(new_n486), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n676), .B1(new_n691), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n688), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI211_X1 g496(.A(KEYINPUT113), .B(KEYINPUT44), .C1(new_n530), .C2(new_n676), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT114), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n525), .B2(new_n529), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n700), .B(new_n529), .C1(new_n689), .C2(new_n690), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n694), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n696), .A3(new_n630), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n687), .B1(new_n699), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n659), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n685), .B1(new_n550), .B2(new_n708), .ZN(G1328gat));
  OAI21_X1  g508(.A(G36gat), .B1(new_n707), .B2(new_n528), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n528), .A2(G36gat), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT46), .B1(new_n678), .B2(new_n712), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n678), .A2(KEYINPUT46), .A3(new_n712), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n710), .A2(new_n713), .A3(new_n714), .ZN(G1329gat));
  INV_X1    g514(.A(G43gat), .ZN(new_n716));
  INV_X1    g515(.A(new_n323), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n716), .B1(new_n706), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n678), .A2(G43gat), .A3(new_n314), .ZN(new_n720));
  OR3_X1    g519(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n718), .B2(new_n720), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1330gat));
  INV_X1    g522(.A(G50gat), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n724), .B1(new_n706), .B2(new_n501), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n678), .A2(G50gat), .A3(new_n411), .ZN(new_n727));
  OR3_X1    g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n725), .B2(new_n727), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(G1331gat));
  NAND2_X1  g529(.A1(new_n691), .A2(KEYINPUT114), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n512), .B1(new_n731), .B2(new_n702), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n578), .A2(new_n631), .A3(new_n654), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n679), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g535(.A(new_n528), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT115), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1333gat));
  INV_X1    g540(.A(G71gat), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n323), .A2(new_n742), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n734), .A2(KEYINPUT116), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT116), .B1(new_n734), .B2(new_n743), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n732), .A2(new_n314), .A3(new_n733), .ZN(new_n746));
  OAI22_X1  g545(.A1(new_n744), .A2(new_n745), .B1(G71gat), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n734), .A2(new_n501), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g549(.A1(new_n577), .A2(new_n599), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n655), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n754), .B1(new_n699), .B2(new_n705), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n755), .A2(new_n679), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n704), .A2(new_n630), .A3(new_n751), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n731), .A2(new_n702), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n676), .B1(new_n760), .B2(new_n694), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(KEYINPUT51), .A3(new_n751), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n654), .A2(new_n679), .A3(new_n604), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n756), .A2(new_n604), .B1(new_n764), .B2(new_n765), .ZN(G1336gat));
  NOR3_X1   g565(.A1(new_n655), .A2(G92gat), .A3(new_n528), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT51), .B1(new_n761), .B2(new_n751), .ZN(new_n768));
  NOR4_X1   g567(.A1(new_n732), .A2(new_n758), .A3(new_n676), .A4(new_n752), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n605), .B1(new_n755), .B2(new_n437), .ZN(new_n776));
  NOR2_X1   g575(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n777), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n773), .B1(new_n763), .B2(new_n767), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n697), .A2(new_n698), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n732), .A2(KEYINPUT44), .A3(new_n676), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n437), .B(new_n753), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G92gat), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n779), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n778), .A2(new_n785), .ZN(G1337gat));
  NAND2_X1  g585(.A1(new_n755), .A2(new_n717), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT118), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G99gat), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n787), .A2(KEYINPUT118), .ZN(new_n790));
  OR3_X1    g589(.A1(new_n655), .A2(G99gat), .A3(new_n314), .ZN(new_n791));
  OAI22_X1  g590(.A1(new_n789), .A2(new_n790), .B1(new_n764), .B2(new_n791), .ZN(G1338gat));
  INV_X1    g591(.A(G106gat), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n755), .B2(new_n501), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n655), .A2(G106gat), .A3(new_n411), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT119), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n759), .B2(new_n762), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT53), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  INV_X1    g598(.A(new_n795), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n764), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n798), .B1(new_n801), .B2(new_n794), .ZN(G1339gat));
  INV_X1    g601(.A(KEYINPUT120), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n645), .A2(new_n646), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n651), .A2(KEYINPUT54), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n641), .B1(new_n650), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(KEYINPUT55), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n649), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT55), .B1(new_n805), .B2(new_n807), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n803), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n810), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n812), .A2(KEYINPUT120), .A3(new_n649), .A4(new_n808), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(new_n813), .A3(new_n577), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n565), .B1(new_n564), .B2(new_n567), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n571), .A2(new_n572), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n534), .ZN(new_n818));
  OR3_X1    g617(.A1(new_n817), .A2(KEYINPUT121), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT121), .B1(new_n817), .B2(new_n818), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n654), .A2(new_n576), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n630), .B1(new_n814), .B2(new_n821), .ZN(new_n822));
  AND4_X1   g621(.A1(new_n576), .A2(new_n819), .A3(new_n630), .A4(new_n820), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n823), .A2(new_n811), .A3(new_n813), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n686), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n656), .A2(new_n577), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n828), .A2(new_n679), .A3(new_n528), .A4(new_n526), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n829), .A2(new_n210), .A3(new_n578), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n659), .B1(new_n825), .B2(new_n827), .ZN(new_n831));
  AND4_X1   g630(.A1(new_n528), .A2(new_n831), .A3(new_n518), .A4(new_n519), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n577), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n830), .B1(new_n833), .B2(new_n210), .ZN(G1340gat));
  NOR3_X1   g633(.A1(new_n829), .A2(new_n208), .A3(new_n655), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n654), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(new_n208), .ZN(G1341gat));
  XOR2_X1   g636(.A(KEYINPUT72), .B(G127gat), .Z(new_n838));
  NOR3_X1   g637(.A1(new_n829), .A2(new_n686), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n832), .A2(new_n599), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(new_n838), .ZN(G1342gat));
  NAND3_X1  g640(.A1(new_n832), .A2(new_n220), .A3(new_n630), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n843));
  OAI21_X1  g642(.A(G134gat), .B1(new_n829), .B2(new_n676), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(G1343gat));
  NOR3_X1   g645(.A1(new_n717), .A2(new_n659), .A3(new_n437), .ZN(new_n847));
  INV_X1    g646(.A(new_n576), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n649), .B(new_n808), .C1(new_n848), .C2(new_n574), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n805), .A2(KEYINPUT122), .A3(new_n807), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT122), .B1(new_n805), .B2(new_n807), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT55), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n821), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n676), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n600), .B1(new_n855), .B2(new_n824), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n411), .B1(new_n856), .B2(new_n827), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n847), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n411), .B1(new_n825), .B2(new_n827), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n860), .A2(new_n858), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(G141gat), .B1(new_n862), .B2(new_n578), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n323), .A2(new_n501), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(new_n437), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n831), .A2(new_n866), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n867), .A2(G141gat), .A3(new_n578), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n863), .A2(new_n864), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n859), .A2(new_n861), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n331), .B1(new_n871), .B2(new_n577), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT58), .B1(new_n872), .B2(new_n868), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n870), .A2(new_n873), .ZN(G1344gat));
  INV_X1    g673(.A(new_n867), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n333), .A3(new_n654), .ZN(new_n876));
  AOI211_X1 g675(.A(KEYINPUT59), .B(new_n333), .C1(new_n871), .C2(new_n654), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n860), .A2(new_n879), .A3(KEYINPUT57), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n823), .A2(new_n649), .A3(new_n808), .A4(new_n812), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n599), .B1(new_n854), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n501), .B1(new_n882), .B2(new_n826), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT123), .B1(new_n883), .B2(new_n858), .ZN(new_n884));
  AOI211_X1 g683(.A(new_n858), .B(new_n411), .C1(new_n825), .C2(new_n827), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n654), .A3(new_n847), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n878), .B1(new_n887), .B2(G148gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n876), .B1(new_n877), .B2(new_n888), .ZN(G1345gat));
  OAI21_X1  g688(.A(G155gat), .B1(new_n862), .B2(new_n686), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n327), .A3(new_n599), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1346gat));
  AOI21_X1  g691(.A(G162gat), .B1(new_n875), .B2(new_n630), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n676), .A2(new_n328), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(new_n871), .B2(new_n894), .ZN(G1347gat));
  NOR2_X1   g694(.A1(new_n679), .A2(new_n528), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n828), .A2(new_n526), .A3(new_n896), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n897), .A2(new_n257), .A3(new_n578), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n679), .B1(new_n825), .B2(new_n827), .ZN(new_n899));
  AND4_X1   g698(.A1(new_n437), .A2(new_n899), .A3(new_n518), .A4(new_n519), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n577), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n898), .B1(new_n901), .B2(new_n257), .ZN(G1348gat));
  NAND3_X1  g701(.A1(new_n900), .A2(new_n258), .A3(new_n654), .ZN(new_n903));
  OAI21_X1  g702(.A(G176gat), .B1(new_n897), .B2(new_n655), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1349gat));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(KEYINPUT60), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n600), .A2(new_n242), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n900), .A2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n236), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n897), .B2(new_n686), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n907), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n906), .A2(KEYINPUT60), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n912), .B(new_n913), .ZN(G1350gat));
  OAI21_X1  g713(.A(G190gat), .B1(new_n897), .B2(new_n676), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT61), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n246), .A3(new_n630), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1351gat));
  NOR2_X1   g717(.A1(new_n865), .A2(new_n528), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n899), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(G197gat), .B1(new_n920), .B2(new_n577), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n896), .A2(new_n323), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n886), .A2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n577), .A2(G197gat), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(G1352gat));
  NOR2_X1   g725(.A1(new_n655), .A2(G204gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n899), .A2(new_n919), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT125), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n929), .A2(KEYINPUT62), .ZN(new_n930));
  OAI21_X1  g729(.A(G204gat), .B1(new_n923), .B2(new_n655), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n929), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n932));
  AOI21_X1  g731(.A(KEYINPUT126), .B1(new_n929), .B2(KEYINPUT62), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n930), .B(new_n931), .C1(new_n932), .C2(new_n933), .ZN(G1353gat));
  NAND3_X1  g733(.A1(new_n920), .A2(new_n368), .A3(new_n599), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n886), .A2(new_n599), .A3(new_n922), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(G1354gat));
  NAND3_X1  g738(.A1(new_n886), .A2(KEYINPUT127), .A3(new_n922), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n630), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT127), .B1(new_n886), .B2(new_n922), .ZN(new_n942));
  OAI21_X1  g741(.A(G218gat), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n920), .A2(new_n349), .A3(new_n630), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1355gat));
endmodule


