

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589;

  XNOR2_X1 U322 ( .A(n341), .B(n291), .ZN(n342) );
  INV_X1 U323 ( .A(KEYINPUT101), .ZN(n470) );
  XOR2_X1 U324 ( .A(n420), .B(n419), .Z(n503) );
  XOR2_X1 U325 ( .A(KEYINPUT36), .B(KEYINPUT100), .Z(n290) );
  XOR2_X1 U326 ( .A(n340), .B(n339), .Z(n291) );
  NAND2_X1 U327 ( .A1(n455), .A2(n538), .ZN(n456) );
  XNOR2_X1 U328 ( .A(n458), .B(KEYINPUT25), .ZN(n459) );
  INV_X1 U329 ( .A(KEYINPUT30), .ZN(n346) );
  XNOR2_X1 U330 ( .A(n460), .B(n459), .ZN(n466) );
  XNOR2_X1 U331 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U332 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n421) );
  XNOR2_X1 U333 ( .A(n349), .B(n348), .ZN(n353) );
  XNOR2_X1 U334 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U335 ( .A(n422), .B(n421), .ZN(n444) );
  XNOR2_X1 U336 ( .A(n412), .B(n411), .ZN(n414) );
  XNOR2_X1 U337 ( .A(n479), .B(n290), .ZN(n587) );
  XNOR2_X1 U338 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U339 ( .A(n358), .B(n357), .Z(n508) );
  XOR2_X1 U340 ( .A(n309), .B(n419), .Z(n538) );
  XOR2_X1 U341 ( .A(KEYINPUT38), .B(n474), .Z(n505) );
  XNOR2_X1 U342 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U343 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(G99GAT), .B(G71GAT), .ZN(n292) );
  XNOR2_X1 U345 ( .A(n292), .B(G120GAT), .ZN(n363) );
  XOR2_X1 U346 ( .A(n363), .B(KEYINPUT81), .Z(n294) );
  XOR2_X1 U347 ( .A(G190GAT), .B(G134GAT), .Z(n338) );
  XNOR2_X1 U348 ( .A(n338), .B(KEYINPUT79), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n304) );
  XOR2_X1 U350 ( .A(KEYINPUT80), .B(KEYINPUT20), .Z(n296) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U352 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U353 ( .A(n297), .B(KEYINPUT78), .Z(n302) );
  XOR2_X1 U354 ( .A(G15GAT), .B(G113GAT), .Z(n299) );
  XNOR2_X1 U355 ( .A(G169GAT), .B(G43GAT), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n349) );
  XNOR2_X1 U357 ( .A(G127GAT), .B(KEYINPUT77), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n300), .B(KEYINPUT0), .ZN(n431) );
  XNOR2_X1 U359 ( .A(n349), .B(n431), .ZN(n301) );
  XNOR2_X1 U360 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n304), .B(n303), .ZN(n309) );
  XOR2_X1 U362 ( .A(G176GAT), .B(KEYINPUT82), .Z(n306) );
  XNOR2_X1 U363 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n308) );
  XOR2_X1 U365 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n419) );
  INV_X1 U367 ( .A(n538), .ZN(n475) );
  XNOR2_X1 U368 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n310), .B(KEYINPUT2), .ZN(n439) );
  XOR2_X1 U370 ( .A(G218GAT), .B(G162GAT), .Z(n335) );
  XOR2_X1 U371 ( .A(n439), .B(n335), .Z(n312) );
  NAND2_X1 U372 ( .A1(G228GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U373 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U374 ( .A(n313), .B(KEYINPUT84), .Z(n315) );
  XOR2_X1 U375 ( .A(G141GAT), .B(G22GAT), .Z(n354) );
  XNOR2_X1 U376 ( .A(G50GAT), .B(n354), .ZN(n314) );
  XNOR2_X1 U377 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U378 ( .A(G204GAT), .B(KEYINPUT24), .Z(n317) );
  XNOR2_X1 U379 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n316) );
  XOR2_X1 U380 ( .A(n317), .B(n316), .Z(n318) );
  XNOR2_X1 U381 ( .A(n319), .B(n318), .ZN(n328) );
  XNOR2_X1 U382 ( .A(G106GAT), .B(G78GAT), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n320), .B(G148GAT), .ZN(n369) );
  INV_X1 U384 ( .A(KEYINPUT21), .ZN(n321) );
  NAND2_X1 U385 ( .A1(G211GAT), .A2(n321), .ZN(n324) );
  INV_X1 U386 ( .A(G211GAT), .ZN(n322) );
  NAND2_X1 U387 ( .A1(n322), .A2(KEYINPUT21), .ZN(n323) );
  NAND2_X1 U388 ( .A1(n324), .A2(n323), .ZN(n326) );
  XNOR2_X1 U389 ( .A(G197GAT), .B(KEYINPUT85), .ZN(n325) );
  XNOR2_X1 U390 ( .A(n326), .B(n325), .ZN(n408) );
  XNOR2_X1 U391 ( .A(n369), .B(n408), .ZN(n327) );
  XNOR2_X1 U392 ( .A(n328), .B(n327), .ZN(n461) );
  XOR2_X1 U393 ( .A(KEYINPUT7), .B(G50GAT), .Z(n330) );
  XNOR2_X1 U394 ( .A(G36GAT), .B(G29GAT), .ZN(n329) );
  XNOR2_X1 U395 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U396 ( .A(KEYINPUT8), .B(n331), .Z(n358) );
  XOR2_X1 U397 ( .A(KEYINPUT71), .B(G106GAT), .Z(n333) );
  XNOR2_X1 U398 ( .A(G43GAT), .B(G99GAT), .ZN(n332) );
  XNOR2_X1 U399 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U400 ( .A(n358), .B(n334), .ZN(n345) );
  XOR2_X1 U401 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n337) );
  XOR2_X1 U402 ( .A(G92GAT), .B(G85GAT), .Z(n359) );
  XNOR2_X1 U403 ( .A(n335), .B(n359), .ZN(n336) );
  XNOR2_X1 U404 ( .A(n337), .B(n336), .ZN(n343) );
  XNOR2_X1 U405 ( .A(n338), .B(KEYINPUT65), .ZN(n341) );
  XOR2_X1 U406 ( .A(KEYINPUT10), .B(KEYINPUT64), .Z(n340) );
  NAND2_X1 U407 ( .A1(G232GAT), .A2(G233GAT), .ZN(n339) );
  XOR2_X1 U408 ( .A(n345), .B(n344), .Z(n558) );
  INV_X1 U409 ( .A(n558), .ZN(n479) );
  NAND2_X1 U410 ( .A1(G229GAT), .A2(G233GAT), .ZN(n347) );
  XOR2_X1 U411 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n351) );
  XNOR2_X1 U412 ( .A(G197GAT), .B(KEYINPUT67), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U414 ( .A(n353), .B(n352), .Z(n356) );
  XOR2_X1 U415 ( .A(G8GAT), .B(G1GAT), .Z(n376) );
  XNOR2_X1 U416 ( .A(n354), .B(n376), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n357) );
  INV_X1 U418 ( .A(n508), .ZN(n574) );
  XOR2_X1 U419 ( .A(G204GAT), .B(G64GAT), .Z(n410) );
  XOR2_X1 U420 ( .A(n359), .B(n410), .Z(n373) );
  XOR2_X1 U421 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n361) );
  XNOR2_X1 U422 ( .A(G176GAT), .B(KEYINPUT70), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n361), .B(n360), .ZN(n367) );
  INV_X1 U424 ( .A(KEYINPUT33), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n365) );
  NAND2_X1 U426 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U428 ( .A(n367), .B(n366), .Z(n371) );
  XNOR2_X1 U429 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n368) );
  XNOR2_X1 U430 ( .A(n368), .B(KEYINPUT69), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n369), .B(n377), .ZN(n370) );
  XNOR2_X1 U432 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U433 ( .A(n373), .B(n372), .ZN(n577) );
  XNOR2_X1 U434 ( .A(KEYINPUT41), .B(n577), .ZN(n507) );
  AND2_X1 U435 ( .A1(n574), .A2(n507), .ZN(n375) );
  XNOR2_X1 U436 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n396) );
  XOR2_X1 U438 ( .A(n377), .B(n376), .Z(n379) );
  NAND2_X1 U439 ( .A1(G231GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U440 ( .A(n379), .B(n378), .ZN(n395) );
  XOR2_X1 U441 ( .A(KEYINPUT75), .B(KEYINPUT12), .Z(n381) );
  XNOR2_X1 U442 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n381), .B(n380), .ZN(n393) );
  XOR2_X1 U444 ( .A(G71GAT), .B(G127GAT), .Z(n383) );
  XNOR2_X1 U445 ( .A(G15GAT), .B(G183GAT), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n391) );
  XOR2_X1 U447 ( .A(KEYINPUT15), .B(KEYINPUT73), .Z(n385) );
  XNOR2_X1 U448 ( .A(KEYINPUT72), .B(KEYINPUT74), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U450 ( .A(G155GAT), .B(G211GAT), .Z(n387) );
  XNOR2_X1 U451 ( .A(G22GAT), .B(G78GAT), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U453 ( .A(n389), .B(n388), .Z(n390) );
  XNOR2_X1 U454 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U455 ( .A(n393), .B(n392), .Z(n394) );
  XNOR2_X1 U456 ( .A(n395), .B(n394), .ZN(n582) );
  NOR2_X1 U457 ( .A1(n396), .A2(n582), .ZN(n397) );
  NAND2_X1 U458 ( .A1(n479), .A2(n397), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n398), .B(KEYINPUT47), .ZN(n399) );
  XNOR2_X1 U460 ( .A(KEYINPUT111), .B(n399), .ZN(n406) );
  XOR2_X1 U461 ( .A(KEYINPUT68), .B(n508), .Z(n561) );
  XOR2_X1 U462 ( .A(KEYINPUT45), .B(KEYINPUT112), .Z(n401) );
  NAND2_X1 U463 ( .A1(n582), .A2(n587), .ZN(n400) );
  XNOR2_X1 U464 ( .A(n401), .B(n400), .ZN(n402) );
  NAND2_X1 U465 ( .A1(n402), .A2(n577), .ZN(n403) );
  NOR2_X1 U466 ( .A1(n561), .A2(n403), .ZN(n404) );
  XNOR2_X1 U467 ( .A(KEYINPUT113), .B(n404), .ZN(n405) );
  NAND2_X1 U468 ( .A1(n406), .A2(n405), .ZN(n407) );
  XNOR2_X1 U469 ( .A(n407), .B(KEYINPUT48), .ZN(n534) );
  XNOR2_X1 U470 ( .A(KEYINPUT88), .B(n408), .ZN(n412) );
  AND2_X1 U471 ( .A1(G226GAT), .A2(G233GAT), .ZN(n409) );
  XOR2_X1 U472 ( .A(G36GAT), .B(G218GAT), .Z(n413) );
  XNOR2_X1 U473 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U474 ( .A(G92GAT), .B(G190GAT), .Z(n416) );
  XNOR2_X1 U475 ( .A(G169GAT), .B(G8GAT), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U477 ( .A(n418), .B(n417), .ZN(n420) );
  INV_X1 U478 ( .A(n503), .ZN(n455) );
  NAND2_X1 U479 ( .A1(n534), .A2(n455), .ZN(n422) );
  XOR2_X1 U480 ( .A(KEYINPUT86), .B(G57GAT), .Z(n424) );
  XNOR2_X1 U481 ( .A(G141GAT), .B(G1GAT), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U483 ( .A(G162GAT), .B(G148GAT), .Z(n426) );
  XNOR2_X1 U484 ( .A(G113GAT), .B(G120GAT), .ZN(n425) );
  XNOR2_X1 U485 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n443) );
  XOR2_X1 U487 ( .A(G85GAT), .B(KEYINPUT71), .Z(n430) );
  XNOR2_X1 U488 ( .A(G29GAT), .B(G134GAT), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n435) );
  XOR2_X1 U490 ( .A(KEYINPUT4), .B(n431), .Z(n433) );
  NAND2_X1 U491 ( .A1(G225GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U493 ( .A(n435), .B(n434), .Z(n441) );
  XOR2_X1 U494 ( .A(KEYINPUT87), .B(KEYINPUT6), .Z(n437) );
  XNOR2_X1 U495 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U497 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U499 ( .A(n443), .B(n442), .Z(n523) );
  INV_X1 U500 ( .A(n523), .ZN(n498) );
  NAND2_X1 U501 ( .A1(n444), .A2(n498), .ZN(n571) );
  NOR2_X1 U502 ( .A1(n461), .A2(n571), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n445), .B(KEYINPUT55), .ZN(n446) );
  NOR2_X1 U504 ( .A1(n475), .A2(n446), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n447), .B(KEYINPUT120), .ZN(n567) );
  NAND2_X1 U506 ( .A1(n567), .A2(n558), .ZN(n451) );
  XOR2_X1 U507 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n449) );
  INV_X1 U508 ( .A(G190GAT), .ZN(n448) );
  INV_X1 U509 ( .A(G43GAT), .ZN(n478) );
  XNOR2_X1 U510 ( .A(KEYINPUT27), .B(n503), .ZN(n463) );
  NOR2_X1 U511 ( .A1(n498), .A2(n463), .ZN(n535) );
  XOR2_X1 U512 ( .A(n461), .B(KEYINPUT28), .Z(n537) );
  INV_X1 U513 ( .A(n537), .ZN(n531) );
  XOR2_X1 U514 ( .A(KEYINPUT83), .B(n538), .Z(n452) );
  NOR2_X1 U515 ( .A1(n531), .A2(n452), .ZN(n453) );
  NAND2_X1 U516 ( .A1(n535), .A2(n453), .ZN(n454) );
  XNOR2_X1 U517 ( .A(n454), .B(KEYINPUT89), .ZN(n469) );
  XNOR2_X1 U518 ( .A(n456), .B(KEYINPUT91), .ZN(n457) );
  NOR2_X1 U519 ( .A1(n461), .A2(n457), .ZN(n460) );
  XNOR2_X1 U520 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n458) );
  NAND2_X1 U521 ( .A1(n475), .A2(n461), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n462), .B(KEYINPUT26), .ZN(n572) );
  NOR2_X1 U523 ( .A1(n572), .A2(n463), .ZN(n464) );
  XNOR2_X1 U524 ( .A(KEYINPUT90), .B(n464), .ZN(n465) );
  NOR2_X1 U525 ( .A1(n466), .A2(n465), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n467), .A2(n523), .ZN(n468) );
  NOR2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n482) );
  NOR2_X1 U528 ( .A1(n582), .A2(n482), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n471), .B(n470), .ZN(n472) );
  NAND2_X1 U530 ( .A1(n472), .A2(n587), .ZN(n473) );
  XOR2_X1 U531 ( .A(KEYINPUT37), .B(n473), .Z(n522) );
  NAND2_X1 U532 ( .A1(n561), .A2(n577), .ZN(n485) );
  NOR2_X1 U533 ( .A1(n522), .A2(n485), .ZN(n474) );
  NOR2_X1 U534 ( .A1(n505), .A2(n475), .ZN(n476) );
  XNOR2_X1 U535 ( .A(KEYINPUT40), .B(n476), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n478), .B(n477), .ZN(G1330GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(KEYINPUT76), .Z(n481) );
  NAND2_X1 U538 ( .A1(n582), .A2(n479), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(n484) );
  INV_X1 U540 ( .A(n482), .ZN(n483) );
  NAND2_X1 U541 ( .A1(n484), .A2(n483), .ZN(n509) );
  NOR2_X1 U542 ( .A1(n485), .A2(n509), .ZN(n486) );
  XNOR2_X1 U543 ( .A(KEYINPUT94), .B(n486), .ZN(n496) );
  NAND2_X1 U544 ( .A1(n496), .A2(n523), .ZN(n489) );
  XOR2_X1 U545 ( .A(G1GAT), .B(KEYINPUT34), .Z(n487) );
  XNOR2_X1 U546 ( .A(KEYINPUT95), .B(n487), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(G1324GAT) );
  NAND2_X1 U548 ( .A1(n496), .A2(n455), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n490), .B(KEYINPUT96), .ZN(n491) );
  XNOR2_X1 U550 ( .A(G8GAT), .B(n491), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT35), .B(KEYINPUT98), .Z(n493) );
  NAND2_X1 U552 ( .A1(n538), .A2(n496), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(n495) );
  XOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT97), .Z(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NAND2_X1 U556 ( .A1(n496), .A2(n531), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n497), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U558 ( .A1(n505), .A2(n498), .ZN(n502) );
  XOR2_X1 U559 ( .A(KEYINPUT99), .B(KEYINPUT102), .Z(n500) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NOR2_X1 U563 ( .A1(n503), .A2(n505), .ZN(n504) );
  XOR2_X1 U564 ( .A(G36GAT), .B(n504), .Z(G1329GAT) );
  NOR2_X1 U565 ( .A1(n537), .A2(n505), .ZN(n506) );
  XOR2_X1 U566 ( .A(G50GAT), .B(n506), .Z(G1331GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n511) );
  NAND2_X1 U568 ( .A1(n508), .A2(n507), .ZN(n521) );
  NOR2_X1 U569 ( .A1(n521), .A2(n509), .ZN(n517) );
  NAND2_X1 U570 ( .A1(n517), .A2(n523), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n514) );
  NAND2_X1 U574 ( .A1(n517), .A2(n455), .ZN(n513) );
  XNOR2_X1 U575 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n517), .A2(n538), .ZN(n516) );
  XNOR2_X1 U578 ( .A(n516), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U580 ( .A1(n517), .A2(n531), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(n520), .ZN(G1335GAT) );
  NOR2_X1 U583 ( .A1(n522), .A2(n521), .ZN(n530) );
  NAND2_X1 U584 ( .A1(n530), .A2(n523), .ZN(n524) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  XOR2_X1 U586 ( .A(G92GAT), .B(KEYINPUT107), .Z(n526) );
  NAND2_X1 U587 ( .A1(n530), .A2(n455), .ZN(n525) );
  XNOR2_X1 U588 ( .A(n526), .B(n525), .ZN(G1337GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n528) );
  NAND2_X1 U590 ( .A1(n530), .A2(n538), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U592 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  NAND2_X1 U593 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U594 ( .A(n532), .B(KEYINPUT44), .ZN(n533) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NAND2_X1 U596 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U597 ( .A(n536), .B(KEYINPUT114), .ZN(n550) );
  NAND2_X1 U598 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U599 ( .A1(n550), .A2(n539), .ZN(n546) );
  NAND2_X1 U600 ( .A1(n546), .A2(n561), .ZN(n540) );
  XNOR2_X1 U601 ( .A(n540), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U603 ( .A1(n546), .A2(n507), .ZN(n541) );
  XNOR2_X1 U604 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n544) );
  NAND2_X1 U606 ( .A1(n546), .A2(n582), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n548) );
  NAND2_X1 U610 ( .A1(n546), .A2(n558), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U612 ( .A(G134GAT), .B(n549), .ZN(G1343GAT) );
  NOR2_X1 U613 ( .A1(n572), .A2(n550), .ZN(n551) );
  XOR2_X1 U614 ( .A(KEYINPUT117), .B(n551), .Z(n557) );
  NAND2_X1 U615 ( .A1(n574), .A2(n557), .ZN(n552) );
  XNOR2_X1 U616 ( .A(n552), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  NAND2_X1 U618 ( .A1(n557), .A2(n507), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n557), .A2(n582), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(KEYINPUT118), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n560), .ZN(G1347GAT) );
  NAND2_X1 U626 ( .A1(n567), .A2(n561), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n567), .A2(n507), .ZN(n564) );
  XOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT121), .Z(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n566) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  NAND2_X1 U633 ( .A1(n567), .A2(n582), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(KEYINPUT124), .ZN(n570) );
  XOR2_X1 U637 ( .A(KEYINPUT59), .B(n570), .Z(n576) );
  OR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(KEYINPUT123), .B(n573), .ZN(n586) );
  NAND2_X1 U640 ( .A1(n586), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n580) );
  INV_X1 U643 ( .A(n577), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n586), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n581), .Z(G1353GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n584) );
  NAND2_X1 U648 ( .A1(n586), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(n585), .ZN(G1354GAT) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

