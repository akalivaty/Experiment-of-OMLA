

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782;

  INV_X1 U376 ( .A(G953), .ZN(n667) );
  XNOR2_X2 U377 ( .A(n373), .B(KEYINPUT80), .ZN(n621) );
  NAND2_X2 U378 ( .A1(n400), .A2(n577), .ZN(n554) );
  XNOR2_X2 U379 ( .A(n562), .B(KEYINPUT38), .ZN(n727) );
  NOR2_X2 U380 ( .A1(n700), .A2(n640), .ZN(n703) );
  XNOR2_X2 U381 ( .A(n501), .B(n500), .ZN(n769) );
  XNOR2_X2 U382 ( .A(n510), .B(G134), .ZN(n501) );
  XNOR2_X2 U383 ( .A(n540), .B(n535), .ZN(n605) );
  NAND2_X1 U384 ( .A1(n417), .A2(n443), .ZN(n416) );
  AND2_X1 U385 ( .A1(n413), .A2(n620), .ZN(n412) );
  XNOR2_X1 U386 ( .A(n600), .B(KEYINPUT32), .ZN(n682) );
  NAND2_X1 U387 ( .A1(n375), .A2(n374), .ZN(n782) );
  AND2_X1 U388 ( .A1(n377), .A2(n376), .ZN(n375) );
  NOR2_X1 U389 ( .A1(n557), .A2(n583), .ZN(n570) );
  NAND2_X2 U390 ( .A1(n438), .A2(n434), .ZN(n713) );
  XNOR2_X1 U391 ( .A(n382), .B(KEYINPUT103), .ZN(n557) );
  XNOR2_X1 U392 ( .A(n456), .B(n455), .ZN(n561) );
  XOR2_X1 U393 ( .A(n651), .B(KEYINPUT59), .Z(n652) );
  XNOR2_X1 U394 ( .A(n769), .B(G146), .ZN(n533) );
  XNOR2_X1 U395 ( .A(KEYINPUT4), .B(G131), .ZN(n500) );
  XNOR2_X1 U396 ( .A(KEYINPUT94), .B(KEYINPUT4), .ZN(n506) );
  INV_X1 U397 ( .A(KEYINPUT60), .ZN(n354) );
  XNOR2_X1 U398 ( .A(n355), .B(n354), .ZN(G60) );
  NAND2_X1 U399 ( .A1(n654), .A2(n691), .ZN(n355) );
  INV_X1 U400 ( .A(KEYINPUT89), .ZN(n386) );
  NOR2_X1 U401 ( .A1(n416), .A2(n409), .ZN(n405) );
  XNOR2_X1 U402 ( .A(G137), .B(KEYINPUT70), .ZN(n527) );
  NOR2_X1 U403 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U404 ( .A(n384), .B(n567), .ZN(n383) );
  OR2_X1 U405 ( .A1(n380), .A2(n422), .ZN(n417) );
  NOR2_X1 U406 ( .A1(n619), .A2(KEYINPUT65), .ZN(n415) );
  OR2_X1 U407 ( .A1(n644), .A2(G902), .ZN(n488) );
  XNOR2_X1 U408 ( .A(n462), .B(n461), .ZN(n558) );
  XNOR2_X1 U409 ( .A(n427), .B(n426), .ZN(n674) );
  INV_X1 U410 ( .A(G104), .ZN(n426) );
  XNOR2_X1 U411 ( .A(G107), .B(G110), .ZN(n427) );
  XNOR2_X1 U412 ( .A(n431), .B(KEYINPUT7), .ZN(n430) );
  INV_X1 U413 ( .A(KEYINPUT9), .ZN(n431) );
  NAND2_X1 U414 ( .A1(n390), .A2(n387), .ZN(n496) );
  AND2_X1 U415 ( .A1(n389), .A2(n388), .ZN(n387) );
  NAND2_X1 U416 ( .A1(n392), .A2(n391), .ZN(n390) );
  NAND2_X1 U417 ( .A1(G237), .A2(KEYINPUT83), .ZN(n389) );
  XNOR2_X1 U418 ( .A(G140), .B(KEYINPUT10), .ZN(n453) );
  XNOR2_X1 U419 ( .A(G104), .B(G113), .ZN(n444) );
  XNOR2_X1 U420 ( .A(n674), .B(KEYINPUT74), .ZN(n531) );
  XNOR2_X1 U421 ( .A(G101), .B(G140), .ZN(n526) );
  XNOR2_X1 U422 ( .A(n539), .B(n359), .ZN(n542) );
  XNOR2_X1 U423 ( .A(n554), .B(n358), .ZN(n588) );
  AND2_X1 U424 ( .A1(n440), .A2(n439), .ZN(n438) );
  NAND2_X1 U425 ( .A1(n503), .A2(G902), .ZN(n439) );
  XNOR2_X1 U426 ( .A(n593), .B(KEYINPUT22), .ZN(n594) );
  INV_X1 U427 ( .A(KEYINPUT82), .ZN(n409) );
  INV_X1 U428 ( .A(KEYINPUT77), .ZN(n423) );
  NOR2_X1 U429 ( .A1(n575), .A2(n574), .ZN(n576) );
  INV_X1 U430 ( .A(G237), .ZN(n518) );
  INV_X1 U431 ( .A(KEYINPUT92), .ZN(n636) );
  NOR2_X1 U432 ( .A1(KEYINPUT83), .A2(G237), .ZN(n392) );
  NAND2_X1 U433 ( .A1(G953), .A2(KEYINPUT83), .ZN(n388) );
  XNOR2_X1 U434 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n446) );
  NAND2_X1 U435 ( .A1(n406), .A2(n405), .ZN(n404) );
  XNOR2_X1 U436 ( .A(KEYINPUT15), .B(G902), .ZN(n641) );
  XOR2_X1 U437 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n508) );
  NAND2_X1 U438 ( .A1(G237), .A2(G234), .ZN(n467) );
  NAND2_X1 U439 ( .A1(n727), .A2(n577), .ZN(n424) );
  NAND2_X1 U440 ( .A1(n437), .A2(n436), .ZN(n435) );
  INV_X1 U441 ( .A(KEYINPUT0), .ZN(n589) );
  XNOR2_X1 U442 ( .A(G137), .B(KEYINPUT81), .ZN(n495) );
  XNOR2_X1 U443 ( .A(KEYINPUT16), .B(G122), .ZN(n515) );
  XNOR2_X1 U444 ( .A(n770), .B(n482), .ZN(n644) );
  BUF_X1 U445 ( .A(n771), .Z(n401) );
  INV_X1 U446 ( .A(KEYINPUT42), .ZN(n378) );
  XNOR2_X1 U447 ( .A(n381), .B(KEYINPUT104), .ZN(n583) );
  NOR2_X1 U448 ( .A1(n561), .A2(n558), .ZN(n381) );
  BUF_X1 U449 ( .A(n540), .Z(n627) );
  XNOR2_X1 U450 ( .A(n460), .B(n428), .ZN(n690) );
  XNOR2_X1 U451 ( .A(n501), .B(n429), .ZN(n428) );
  XNOR2_X1 U452 ( .A(n459), .B(n430), .ZN(n429) );
  XNOR2_X1 U453 ( .A(n363), .B(n451), .ZN(n651) );
  XNOR2_X1 U454 ( .A(n533), .B(n410), .ZN(n695) );
  XNOR2_X1 U455 ( .A(n531), .B(n532), .ZN(n410) );
  AND2_X1 U456 ( .A1(n599), .A2(n596), .ZN(n369) );
  XNOR2_X1 U457 ( .A(n566), .B(KEYINPUT108), .ZN(n779) );
  NAND2_X1 U458 ( .A1(n370), .A2(n588), .ZN(n758) );
  OR2_X1 U459 ( .A1(n604), .A2(n603), .ZN(n666) );
  XNOR2_X1 U460 ( .A(n394), .B(n635), .ZN(n681) );
  AND2_X1 U461 ( .A1(n634), .A2(n596), .ZN(n393) );
  AND2_X1 U462 ( .A1(n408), .A2(n407), .ZN(n356) );
  INV_X1 U463 ( .A(G902), .ZN(n436) );
  OR2_X1 U464 ( .A1(n555), .A2(n378), .ZN(n357) );
  XOR2_X1 U465 ( .A(KEYINPUT67), .B(KEYINPUT19), .Z(n358) );
  XOR2_X1 U466 ( .A(KEYINPUT28), .B(KEYINPUT110), .Z(n359) );
  AND2_X1 U467 ( .A1(n620), .A2(n618), .ZN(n360) );
  NAND2_X1 U468 ( .A1(n638), .A2(n639), .ZN(n361) );
  NAND2_X1 U469 ( .A1(n639), .A2(KEYINPUT90), .ZN(n362) );
  INV_X1 U470 ( .A(G953), .ZN(n391) );
  NAND2_X1 U471 ( .A1(n683), .A2(KEYINPUT44), .ZN(n402) );
  NAND2_X1 U472 ( .A1(n369), .A2(n601), .ZN(n600) );
  AND2_X1 U473 ( .A1(n681), .A2(n372), .ZN(n403) );
  XNOR2_X1 U474 ( .A(n452), .B(n475), .ZN(n363) );
  NOR2_X1 U475 ( .A1(n572), .A2(n758), .ZN(n573) );
  XNOR2_X2 U476 ( .A(n364), .B(KEYINPUT45), .ZN(n668) );
  NAND2_X1 U477 ( .A1(n367), .A2(n365), .ZN(n364) );
  NAND2_X1 U478 ( .A1(n366), .A2(n414), .ZN(n365) );
  NAND2_X1 U479 ( .A1(n412), .A2(n415), .ZN(n366) );
  XNOR2_X1 U480 ( .A(n368), .B(n636), .ZN(n367) );
  NAND2_X1 U481 ( .A1(n403), .A2(n402), .ZN(n368) );
  INV_X1 U482 ( .A(n555), .ZN(n370) );
  NAND2_X2 U483 ( .A1(n371), .A2(n420), .ZN(n418) );
  NAND2_X1 U484 ( .A1(n419), .A2(n379), .ZN(n371) );
  NAND2_X1 U485 ( .A1(n632), .A2(n724), .ZN(n372) );
  OR2_X2 U486 ( .A1(n718), .A2(n631), .ZN(n626) );
  NAND2_X1 U487 ( .A1(n416), .A2(n409), .ZN(n407) );
  NOR2_X2 U488 ( .A1(n605), .A2(n706), .ZN(n373) );
  XNOR2_X1 U489 ( .A(n607), .B(KEYINPUT33), .ZN(n723) );
  XNOR2_X2 U490 ( .A(n595), .B(n594), .ZN(n601) );
  OR2_X1 U491 ( .A1(n743), .A2(n357), .ZN(n374) );
  XNOR2_X2 U492 ( .A(n544), .B(n543), .ZN(n743) );
  NOR2_X2 U493 ( .A1(n781), .A2(n782), .ZN(n552) );
  NAND2_X1 U494 ( .A1(n555), .A2(n378), .ZN(n376) );
  NAND2_X1 U495 ( .A1(n743), .A2(n378), .ZN(n377) );
  INV_X1 U496 ( .A(n421), .ZN(n379) );
  NAND2_X1 U497 ( .A1(n553), .A2(n767), .ZN(n421) );
  AND2_X1 U498 ( .A1(n380), .A2(n422), .ZN(n419) );
  XNOR2_X1 U499 ( .A(n576), .B(n423), .ZN(n380) );
  NAND2_X1 U500 ( .A1(n561), .A2(n558), .ZN(n382) );
  NAND2_X1 U501 ( .A1(n568), .A2(n383), .ZN(n575) );
  NAND2_X1 U502 ( .A1(n779), .A2(n385), .ZN(n384) );
  XNOR2_X1 U503 ( .A(n559), .B(n386), .ZN(n385) );
  NAND2_X1 U504 ( .A1(n496), .A2(G214), .ZN(n450) );
  NAND2_X1 U505 ( .A1(n601), .A2(n393), .ZN(n394) );
  XNOR2_X2 U506 ( .A(n395), .B(n643), .ZN(n693) );
  NAND2_X1 U507 ( .A1(n399), .A2(n396), .ZN(n395) );
  NAND2_X1 U508 ( .A1(n398), .A2(n397), .ZN(n396) );
  NAND2_X1 U509 ( .A1(n433), .A2(n362), .ZN(n397) );
  NAND2_X1 U510 ( .A1(n432), .A2(n361), .ZN(n398) );
  NOR2_X1 U511 ( .A1(n703), .A2(n642), .ZN(n399) );
  NAND2_X1 U512 ( .A1(n421), .A2(KEYINPUT48), .ZN(n420) );
  NAND2_X1 U513 ( .A1(n682), .A2(n666), .ZN(n619) );
  NAND2_X1 U514 ( .A1(n588), .A2(n442), .ZN(n590) );
  INV_X1 U515 ( .A(n562), .ZN(n400) );
  XNOR2_X2 U516 ( .A(n522), .B(n521), .ZN(n562) );
  NAND2_X1 U517 ( .A1(n356), .A2(n404), .ZN(n637) );
  XNOR2_X2 U518 ( .A(n488), .B(n487), .ZN(n710) );
  NAND2_X1 U519 ( .A1(n619), .A2(n360), .ZN(n414) );
  XNOR2_X2 U520 ( .A(n614), .B(n613), .ZN(n683) );
  INV_X1 U521 ( .A(n418), .ZN(n406) );
  NAND2_X1 U522 ( .A1(n418), .A2(n409), .ZN(n408) );
  NOR2_X1 U523 ( .A1(n418), .A2(n416), .ZN(n771) );
  NAND2_X1 U524 ( .A1(n411), .A2(n736), .ZN(n744) );
  INV_X1 U525 ( .A(n743), .ZN(n411) );
  NAND2_X1 U526 ( .A1(n616), .A2(n615), .ZN(n413) );
  INV_X1 U527 ( .A(KEYINPUT48), .ZN(n422) );
  NAND2_X1 U528 ( .A1(n725), .A2(n731), .ZN(n544) );
  XNOR2_X2 U529 ( .A(n424), .B(KEYINPUT111), .ZN(n725) );
  XNOR2_X2 U530 ( .A(n425), .B(n534), .ZN(n540) );
  OR2_X2 U531 ( .A1(n695), .A2(G902), .ZN(n425) );
  INV_X1 U532 ( .A(n583), .ZN(n764) );
  INV_X1 U533 ( .A(n557), .ZN(n760) );
  INV_X1 U534 ( .A(n570), .ZN(n724) );
  NAND2_X1 U535 ( .A1(n570), .A2(KEYINPUT47), .ZN(n559) );
  XNOR2_X2 U536 ( .A(G143), .B(G128), .ZN(n510) );
  INV_X1 U537 ( .A(n433), .ZN(n432) );
  NAND2_X1 U538 ( .A1(n637), .A2(n668), .ZN(n433) );
  OR2_X1 U539 ( .A1(n684), .A2(n435), .ZN(n434) );
  INV_X1 U540 ( .A(n503), .ZN(n437) );
  NAND2_X1 U541 ( .A1(n684), .A2(n503), .ZN(n440) );
  XNOR2_X1 U542 ( .A(n441), .B(n545), .ZN(n549) );
  NAND2_X1 U543 ( .A1(n713), .A2(n577), .ZN(n441) );
  NAND2_X1 U544 ( .A1(n648), .A2(n691), .ZN(n650) );
  XNOR2_X1 U545 ( .A(n646), .B(n645), .ZN(n648) );
  BUF_X1 U546 ( .A(n562), .Z(n581) );
  OR2_X1 U547 ( .A1(n587), .A2(n586), .ZN(n442) );
  AND2_X1 U548 ( .A1(n664), .A2(n768), .ZN(n443) );
  INV_X1 U549 ( .A(KEYINPUT86), .ZN(n567) );
  INV_X1 U550 ( .A(KEYINPUT124), .ZN(n649) );
  XOR2_X1 U551 ( .A(KEYINPUT101), .B(G122), .Z(n445) );
  XNOR2_X1 U552 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U553 ( .A(G131), .B(G143), .Z(n447) );
  XNOR2_X1 U554 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U555 ( .A(n449), .B(n448), .ZN(n452) );
  XNOR2_X1 U556 ( .A(n450), .B(KEYINPUT100), .ZN(n451) );
  XNOR2_X1 U557 ( .A(n453), .B(KEYINPUT69), .ZN(n454) );
  XNOR2_X1 U558 ( .A(G146), .B(G125), .ZN(n511) );
  XNOR2_X2 U559 ( .A(n454), .B(n511), .ZN(n475) );
  NAND2_X1 U560 ( .A1(n651), .A2(n436), .ZN(n456) );
  XOR2_X1 U561 ( .A(KEYINPUT13), .B(G475), .Z(n455) );
  AND2_X1 U562 ( .A1(G234), .A2(n667), .ZN(n457) );
  XNOR2_X1 U563 ( .A(n457), .B(KEYINPUT8), .ZN(n479) );
  NAND2_X1 U564 ( .A1(n479), .A2(G217), .ZN(n458) );
  XNOR2_X1 U565 ( .A(n458), .B(G122), .ZN(n460) );
  XNOR2_X1 U566 ( .A(G107), .B(G116), .ZN(n459) );
  NAND2_X1 U567 ( .A1(n690), .A2(n436), .ZN(n462) );
  XOR2_X1 U568 ( .A(KEYINPUT102), .B(G478), .Z(n461) );
  NAND2_X1 U569 ( .A1(n641), .A2(G234), .ZN(n464) );
  INV_X1 U570 ( .A(KEYINPUT20), .ZN(n463) );
  XNOR2_X1 U571 ( .A(n464), .B(n463), .ZN(n483) );
  INV_X1 U572 ( .A(G221), .ZN(n465) );
  OR2_X1 U573 ( .A1(n483), .A2(n465), .ZN(n466) );
  XNOR2_X1 U574 ( .A(n466), .B(KEYINPUT21), .ZN(n709) );
  XNOR2_X1 U575 ( .A(n467), .B(KEYINPUT14), .ZN(n468) );
  NAND2_X1 U576 ( .A1(G952), .A2(n468), .ZN(n742) );
  NOR2_X1 U577 ( .A1(n742), .A2(G953), .ZN(n586) );
  NAND2_X1 U578 ( .A1(G902), .A2(n468), .ZN(n469) );
  XOR2_X1 U579 ( .A(KEYINPUT96), .B(n469), .Z(n470) );
  NAND2_X1 U580 ( .A1(G953), .A2(n470), .ZN(n585) );
  NOR2_X1 U581 ( .A1(n585), .A2(G900), .ZN(n471) );
  NOR2_X1 U582 ( .A1(n586), .A2(n471), .ZN(n472) );
  NOR2_X1 U583 ( .A1(n709), .A2(n472), .ZN(n546) );
  XNOR2_X1 U584 ( .A(KEYINPUT71), .B(n546), .ZN(n537) );
  INV_X1 U585 ( .A(n537), .ZN(n473) );
  NAND2_X1 U586 ( .A1(n557), .A2(n473), .ZN(n489) );
  INV_X1 U587 ( .A(n527), .ZN(n474) );
  XNOR2_X2 U588 ( .A(n475), .B(n474), .ZN(n770) );
  XNOR2_X1 U589 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n478) );
  XNOR2_X1 U590 ( .A(G119), .B(G110), .ZN(n476) );
  XNOR2_X1 U591 ( .A(G128), .B(n476), .ZN(n477) );
  XNOR2_X1 U592 ( .A(n478), .B(n477), .ZN(n481) );
  NAND2_X1 U593 ( .A1(n479), .A2(G221), .ZN(n480) );
  XNOR2_X1 U594 ( .A(n481), .B(n480), .ZN(n482) );
  INV_X1 U595 ( .A(n483), .ZN(n484) );
  AND2_X1 U596 ( .A1(n484), .A2(G217), .ZN(n486) );
  XNOR2_X1 U597 ( .A(KEYINPUT97), .B(KEYINPUT25), .ZN(n485) );
  XNOR2_X1 U598 ( .A(n486), .B(n485), .ZN(n487) );
  INV_X1 U599 ( .A(n710), .ZN(n633) );
  NOR2_X1 U600 ( .A1(n489), .A2(n633), .ZN(n505) );
  XNOR2_X1 U601 ( .A(G119), .B(G116), .ZN(n491) );
  XNOR2_X1 U602 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n490) );
  XNOR2_X1 U603 ( .A(n491), .B(n490), .ZN(n494) );
  XNOR2_X1 U604 ( .A(G113), .B(G101), .ZN(n492) );
  XNOR2_X1 U605 ( .A(n492), .B(KEYINPUT3), .ZN(n493) );
  XNOR2_X1 U606 ( .A(n494), .B(n493), .ZN(n516) );
  XNOR2_X1 U607 ( .A(n495), .B(KEYINPUT5), .ZN(n498) );
  NAND2_X1 U608 ( .A1(n496), .A2(G210), .ZN(n497) );
  XNOR2_X1 U609 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U610 ( .A(n516), .B(n499), .ZN(n502) );
  XNOR2_X1 U611 ( .A(n533), .B(n502), .ZN(n684) );
  XNOR2_X1 U612 ( .A(G472), .B(KEYINPUT98), .ZN(n503) );
  INV_X1 U613 ( .A(n713), .ZN(n504) );
  XNOR2_X1 U614 ( .A(n504), .B(KEYINPUT6), .ZN(n606) );
  NAND2_X1 U615 ( .A1(n505), .A2(n606), .ZN(n579) );
  XOR2_X1 U616 ( .A(n579), .B(KEYINPUT113), .Z(n524) );
  NAND2_X1 U617 ( .A1(G224), .A2(n667), .ZN(n507) );
  XNOR2_X1 U618 ( .A(n507), .B(n506), .ZN(n509) );
  XNOR2_X1 U619 ( .A(n509), .B(n508), .ZN(n513) );
  XNOR2_X1 U620 ( .A(n510), .B(n511), .ZN(n512) );
  XNOR2_X1 U621 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U622 ( .A(n514), .B(n531), .ZN(n517) );
  XNOR2_X1 U623 ( .A(n516), .B(n515), .ZN(n675) );
  XNOR2_X1 U624 ( .A(n517), .B(n675), .ZN(n655) );
  NAND2_X1 U625 ( .A1(n655), .A2(n641), .ZN(n522) );
  NAND2_X1 U626 ( .A1(n436), .A2(n518), .ZN(n523) );
  NAND2_X1 U627 ( .A1(n523), .A2(G210), .ZN(n520) );
  INV_X1 U628 ( .A(KEYINPUT95), .ZN(n519) );
  XNOR2_X1 U629 ( .A(n520), .B(n519), .ZN(n521) );
  AND2_X1 U630 ( .A1(n523), .A2(G214), .ZN(n728) );
  NOR2_X1 U631 ( .A1(n524), .A2(n554), .ZN(n525) );
  XNOR2_X1 U632 ( .A(n525), .B(KEYINPUT36), .ZN(n536) );
  XNOR2_X1 U633 ( .A(n527), .B(n526), .ZN(n530) );
  NAND2_X1 U634 ( .A1(n667), .A2(G227), .ZN(n528) );
  XNOR2_X1 U635 ( .A(n528), .B(KEYINPUT84), .ZN(n529) );
  XNOR2_X1 U636 ( .A(n530), .B(n529), .ZN(n532) );
  INV_X1 U637 ( .A(G469), .ZN(n534) );
  XNOR2_X1 U638 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n535) );
  BUF_X2 U639 ( .A(n605), .Z(n707) );
  XNOR2_X1 U640 ( .A(n707), .B(KEYINPUT93), .ZN(n597) );
  NAND2_X1 U641 ( .A1(n536), .A2(n597), .ZN(n767) );
  NOR2_X1 U642 ( .A1(n537), .A2(n633), .ZN(n538) );
  NAND2_X1 U643 ( .A1(n538), .A2(n713), .ZN(n539) );
  XNOR2_X1 U644 ( .A(n627), .B(KEYINPUT109), .ZN(n541) );
  NAND2_X1 U645 ( .A1(n542), .A2(n541), .ZN(n555) );
  INV_X1 U646 ( .A(n728), .ZN(n577) );
  INV_X1 U647 ( .A(n558), .ZN(n560) );
  OR2_X1 U648 ( .A1(n561), .A2(n560), .ZN(n591) );
  INV_X1 U649 ( .A(n591), .ZN(n731) );
  XOR2_X1 U650 ( .A(KEYINPUT41), .B(KEYINPUT112), .Z(n543) );
  XNOR2_X1 U651 ( .A(KEYINPUT30), .B(KEYINPUT107), .ZN(n545) );
  NAND2_X1 U652 ( .A1(n633), .A2(n546), .ZN(n547) );
  NOR2_X1 U653 ( .A1(n627), .A2(n547), .ZN(n548) );
  AND2_X1 U654 ( .A1(n549), .A2(n548), .ZN(n565) );
  NAND2_X1 U655 ( .A1(n565), .A2(n727), .ZN(n550) );
  XNOR2_X1 U656 ( .A(n550), .B(KEYINPUT39), .ZN(n584) );
  AND2_X1 U657 ( .A1(n557), .A2(n584), .ZN(n551) );
  XNOR2_X1 U658 ( .A(n551), .B(KEYINPUT40), .ZN(n781) );
  XNOR2_X1 U659 ( .A(n552), .B(KEYINPUT46), .ZN(n553) );
  NAND2_X1 U660 ( .A1(n758), .A2(KEYINPUT47), .ZN(n556) );
  XNOR2_X1 U661 ( .A(n556), .B(KEYINPUT88), .ZN(n568) );
  AND2_X1 U662 ( .A1(n561), .A2(n560), .ZN(n610) );
  INV_X1 U663 ( .A(n610), .ZN(n563) );
  NOR2_X1 U664 ( .A1(n563), .A2(n581), .ZN(n564) );
  NAND2_X1 U665 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U666 ( .A(KEYINPUT68), .B(KEYINPUT47), .ZN(n569) );
  XNOR2_X1 U667 ( .A(n571), .B(KEYINPUT79), .ZN(n572) );
  XNOR2_X1 U668 ( .A(n573), .B(KEYINPUT78), .ZN(n574) );
  NAND2_X1 U669 ( .A1(n707), .A2(n577), .ZN(n578) );
  OR2_X1 U670 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U671 ( .A(n580), .B(KEYINPUT43), .ZN(n582) );
  NAND2_X1 U672 ( .A1(n582), .A2(n581), .ZN(n664) );
  NAND2_X1 U673 ( .A1(n584), .A2(n583), .ZN(n768) );
  NOR2_X1 U674 ( .A1(n585), .A2(G898), .ZN(n587) );
  XNOR2_X2 U675 ( .A(n590), .B(n589), .ZN(n624) );
  NOR2_X1 U676 ( .A1(n591), .A2(n709), .ZN(n592) );
  NAND2_X1 U677 ( .A1(n624), .A2(n592), .ZN(n595) );
  INV_X1 U678 ( .A(KEYINPUT76), .ZN(n593) );
  INV_X1 U679 ( .A(n606), .ZN(n596) );
  AND2_X1 U680 ( .A1(n597), .A2(n710), .ZN(n598) );
  XNOR2_X1 U681 ( .A(n598), .B(KEYINPUT106), .ZN(n599) );
  INV_X1 U682 ( .A(n601), .ZN(n604) );
  NOR2_X1 U683 ( .A1(n713), .A2(n633), .ZN(n602) );
  NAND2_X1 U684 ( .A1(n707), .A2(n602), .ZN(n603) );
  OR2_X2 U685 ( .A1(n710), .A2(n709), .ZN(n706) );
  NAND2_X1 U686 ( .A1(n621), .A2(n606), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n723), .A2(n624), .ZN(n609) );
  XNOR2_X1 U688 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n608) );
  XNOR2_X1 U689 ( .A(n609), .B(n608), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n611), .A2(n610), .ZN(n614) );
  INV_X1 U691 ( .A(KEYINPUT85), .ZN(n612) );
  XNOR2_X1 U692 ( .A(n612), .B(KEYINPUT35), .ZN(n613) );
  INV_X1 U693 ( .A(n683), .ZN(n616) );
  INV_X1 U694 ( .A(KEYINPUT44), .ZN(n615) );
  INV_X1 U695 ( .A(KEYINPUT65), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n617), .A2(KEYINPUT44), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n615), .A2(KEYINPUT65), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n713), .ZN(n623) );
  INV_X1 U699 ( .A(KEYINPUT99), .ZN(n622) );
  XNOR2_X1 U700 ( .A(n623), .B(n622), .ZN(n718) );
  INV_X1 U701 ( .A(n624), .ZN(n631) );
  INV_X1 U702 ( .A(KEYINPUT31), .ZN(n625) );
  XNOR2_X2 U703 ( .A(n626), .B(n625), .ZN(n763) );
  NOR2_X1 U704 ( .A1(n713), .A2(n706), .ZN(n629) );
  INV_X1 U705 ( .A(n627), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n630) );
  OR2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n753) );
  NAND2_X1 U708 ( .A1(n763), .A2(n753), .ZN(n632) );
  AND2_X1 U709 ( .A1(n707), .A2(n633), .ZN(n634) );
  INV_X1 U710 ( .A(KEYINPUT105), .ZN(n635) );
  NOR2_X1 U711 ( .A1(n641), .A2(KEYINPUT90), .ZN(n638) );
  INV_X1 U712 ( .A(KEYINPUT2), .ZN(n639) );
  NAND2_X1 U713 ( .A1(n771), .A2(KEYINPUT2), .ZN(n640) );
  INV_X1 U714 ( .A(n668), .ZN(n700) );
  AND2_X1 U715 ( .A1(n641), .A2(KEYINPUT90), .ZN(n642) );
  INV_X1 U716 ( .A(KEYINPUT64), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n693), .A2(G217), .ZN(n646) );
  INV_X1 U718 ( .A(n644), .ZN(n645) );
  INV_X1 U719 ( .A(G952), .ZN(n647) );
  NAND2_X1 U720 ( .A1(n647), .A2(G953), .ZN(n691) );
  XNOR2_X1 U721 ( .A(n650), .B(n649), .ZN(G66) );
  NAND2_X1 U722 ( .A1(n693), .A2(G475), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n653), .B(n652), .ZN(n654) );
  NAND2_X1 U724 ( .A1(n693), .A2(G210), .ZN(n660) );
  BUF_X1 U725 ( .A(n655), .Z(n656) );
  XNOR2_X1 U726 ( .A(KEYINPUT87), .B(KEYINPUT54), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n657), .B(KEYINPUT55), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n656), .B(n658), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U730 ( .A1(n661), .A2(n691), .ZN(n663) );
  INV_X1 U731 ( .A(KEYINPUT56), .ZN(n662) );
  XNOR2_X1 U732 ( .A(n663), .B(n662), .ZN(G51) );
  XNOR2_X1 U733 ( .A(n664), .B(G140), .ZN(G42) );
  XOR2_X1 U734 ( .A(G110), .B(KEYINPUT115), .Z(n665) );
  XNOR2_X1 U735 ( .A(n666), .B(n665), .ZN(G12) );
  NAND2_X1 U736 ( .A1(n668), .A2(n391), .ZN(n673) );
  NAND2_X1 U737 ( .A1(G953), .A2(G224), .ZN(n669) );
  XNOR2_X1 U738 ( .A(KEYINPUT61), .B(n669), .ZN(n670) );
  NAND2_X1 U739 ( .A1(n670), .A2(G898), .ZN(n671) );
  XOR2_X1 U740 ( .A(KEYINPUT125), .B(n671), .Z(n672) );
  NAND2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n680) );
  XNOR2_X1 U742 ( .A(n675), .B(n674), .ZN(n677) );
  NOR2_X1 U743 ( .A1(n391), .A2(G898), .ZN(n676) );
  NOR2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U745 ( .A(n678), .B(KEYINPUT126), .ZN(n679) );
  XNOR2_X1 U746 ( .A(n680), .B(n679), .ZN(G69) );
  XNOR2_X1 U747 ( .A(n681), .B(G101), .ZN(G3) );
  XNOR2_X1 U748 ( .A(n682), .B(G119), .ZN(G21) );
  XOR2_X1 U749 ( .A(n683), .B(G122), .Z(G24) );
  NAND2_X1 U750 ( .A1(n693), .A2(G472), .ZN(n686) );
  XOR2_X1 U751 ( .A(KEYINPUT62), .B(n684), .Z(n685) );
  XNOR2_X1 U752 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U753 ( .A1(n687), .A2(n691), .ZN(n688) );
  XNOR2_X1 U754 ( .A(n688), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U755 ( .A1(n693), .A2(G478), .ZN(n689) );
  XOR2_X1 U756 ( .A(n690), .B(n689), .Z(n692) );
  INV_X1 U757 ( .A(n691), .ZN(n698) );
  NOR2_X1 U758 ( .A1(n692), .A2(n698), .ZN(G63) );
  NAND2_X1 U759 ( .A1(n693), .A2(G469), .ZN(n697) );
  XOR2_X1 U760 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n694) );
  XNOR2_X1 U761 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U762 ( .A(n697), .B(n696), .ZN(n699) );
  NOR2_X1 U763 ( .A1(n699), .A2(n698), .ZN(G54) );
  INV_X1 U764 ( .A(n401), .ZN(n701) );
  NOR2_X1 U765 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U766 ( .A1(n702), .A2(KEYINPUT2), .ZN(n704) );
  NOR2_X1 U767 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U768 ( .A(n705), .B(KEYINPUT91), .ZN(n748) );
  NAND2_X1 U769 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U770 ( .A(n708), .B(KEYINPUT50), .ZN(n716) );
  XOR2_X1 U771 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n712) );
  NAND2_X1 U772 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U773 ( .A(n712), .B(n711), .Z(n714) );
  NOR2_X1 U774 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U775 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U776 ( .A(KEYINPUT119), .B(n717), .Z(n719) );
  NAND2_X1 U777 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U778 ( .A(KEYINPUT51), .B(n720), .ZN(n721) );
  NOR2_X1 U779 ( .A1(n743), .A2(n721), .ZN(n722) );
  XOR2_X1 U780 ( .A(KEYINPUT120), .B(n722), .Z(n738) );
  BUF_X1 U781 ( .A(n723), .Z(n736) );
  NAND2_X1 U782 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U783 ( .A(KEYINPUT122), .B(n726), .ZN(n734) );
  INV_X1 U784 ( .A(n727), .ZN(n729) );
  NAND2_X1 U785 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U786 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U787 ( .A(KEYINPUT121), .B(n732), .Z(n733) );
  NAND2_X1 U788 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U789 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U790 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U791 ( .A(n739), .B(KEYINPUT123), .ZN(n740) );
  XNOR2_X1 U792 ( .A(n740), .B(KEYINPUT52), .ZN(n741) );
  NOR2_X1 U793 ( .A1(n742), .A2(n741), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n744), .A2(n391), .ZN(n745) );
  NOR2_X1 U795 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U796 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U797 ( .A(KEYINPUT53), .B(n749), .Z(G75) );
  NOR2_X1 U798 ( .A1(n753), .A2(n760), .ZN(n750) );
  XOR2_X1 U799 ( .A(G104), .B(n750), .Z(G6) );
  XOR2_X1 U800 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n752) );
  XNOR2_X1 U801 ( .A(G107), .B(KEYINPUT114), .ZN(n751) );
  XNOR2_X1 U802 ( .A(n752), .B(n751), .ZN(n755) );
  NOR2_X1 U803 ( .A1(n753), .A2(n764), .ZN(n754) );
  XOR2_X1 U804 ( .A(n755), .B(n754), .Z(G9) );
  NOR2_X1 U805 ( .A1(n758), .A2(n764), .ZN(n757) );
  XNOR2_X1 U806 ( .A(G128), .B(KEYINPUT29), .ZN(n756) );
  XNOR2_X1 U807 ( .A(n757), .B(n756), .ZN(G30) );
  NOR2_X1 U808 ( .A1(n758), .A2(n760), .ZN(n759) );
  XOR2_X1 U809 ( .A(G146), .B(n759), .Z(G48) );
  NOR2_X1 U810 ( .A1(n760), .A2(n763), .ZN(n762) );
  XNOR2_X1 U811 ( .A(G113), .B(KEYINPUT117), .ZN(n761) );
  XNOR2_X1 U812 ( .A(n762), .B(n761), .ZN(G15) );
  NOR2_X1 U813 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U814 ( .A(G116), .B(n765), .Z(G18) );
  XOR2_X1 U815 ( .A(G125), .B(KEYINPUT37), .Z(n766) );
  XNOR2_X1 U816 ( .A(n767), .B(n766), .ZN(G27) );
  XNOR2_X1 U817 ( .A(G134), .B(n768), .ZN(G36) );
  XNOR2_X1 U818 ( .A(n769), .B(n770), .ZN(n773) );
  XNOR2_X1 U819 ( .A(n401), .B(n773), .ZN(n772) );
  NAND2_X1 U820 ( .A1(n772), .A2(n391), .ZN(n778) );
  XOR2_X1 U821 ( .A(G227), .B(n773), .Z(n774) );
  NAND2_X1 U822 ( .A1(n774), .A2(G900), .ZN(n775) );
  NAND2_X1 U823 ( .A1(G953), .A2(n775), .ZN(n776) );
  XOR2_X1 U824 ( .A(KEYINPUT127), .B(n776), .Z(n777) );
  NAND2_X1 U825 ( .A1(n778), .A2(n777), .ZN(G72) );
  XNOR2_X1 U826 ( .A(G143), .B(n779), .ZN(n780) );
  XNOR2_X1 U827 ( .A(n780), .B(KEYINPUT116), .ZN(G45) );
  XOR2_X1 U828 ( .A(G131), .B(n781), .Z(G33) );
  XOR2_X1 U829 ( .A(n782), .B(G137), .Z(G39) );
endmodule

