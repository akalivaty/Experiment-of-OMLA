//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n543, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n469), .C1(new_n462), .C2(new_n463), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n469), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n473));
  AND3_X1   g048(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n470), .B2(new_n472), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n464), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n464), .A2(new_n469), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G138), .B(new_n469), .C1(new_n462), .C2(new_n463), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT3), .B(G2104), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .A3(G138), .A4(new_n469), .ZN(new_n490));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(new_n494), .A3(G2104), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n488), .A2(new_n490), .A3(new_n491), .A4(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  NAND2_X1  g072(.A1(G75), .A2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G62), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(KEYINPUT67), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT67), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT6), .A3(G651), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n499), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n505), .A2(G651), .B1(G50), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n503), .B1(new_n508), .B2(new_n510), .ZN(new_n513));
  XOR2_X1   g088(.A(KEYINPUT68), .B(G88), .Z(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n519));
  INV_X1    g094(.A(new_n511), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT69), .B(G51), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(KEYINPUT70), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(KEYINPUT70), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n523), .A2(new_n524), .B1(G89), .B2(new_n513), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  AOI22_X1  g104(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(new_n507), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n513), .A2(G90), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n511), .A2(G52), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G56), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n503), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n538), .A2(G651), .B1(G43), .B2(new_n511), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n513), .A2(G81), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G188));
  NAND2_X1  g122(.A1(new_n511), .A2(G53), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT9), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n509), .A2(KEYINPUT6), .A3(G651), .ZN(new_n550));
  AOI21_X1  g125(.A(KEYINPUT6), .B1(new_n509), .B2(G651), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n518), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n508), .A2(new_n510), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n555), .A2(KEYINPUT71), .A3(new_n518), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G91), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT72), .B1(new_n559), .B2(new_n507), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n503), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n563), .A2(new_n564), .A3(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n549), .A2(new_n558), .A3(new_n566), .ZN(G299));
  NAND2_X1  g142(.A1(new_n557), .A2(G87), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n518), .A2(G74), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(G49), .B2(new_n511), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(G288));
  NAND2_X1  g146(.A1(new_n511), .A2(G48), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n557), .B2(G86), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n518), .B2(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n575), .B1(new_n578), .B2(new_n507), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n576), .B1(new_n503), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n581), .A2(KEYINPUT73), .A3(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n574), .A2(new_n583), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(KEYINPUT74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(KEYINPUT74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(G47), .B2(new_n511), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n513), .A2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n557), .A2(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n557), .A2(KEYINPUT10), .A3(G92), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n503), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n596), .A2(new_n597), .B1(G651), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n511), .A2(G54), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n593), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n593), .B1(new_n604), .B2(G868), .ZN(G321));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G299), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G168), .B2(new_n607), .ZN(G280));
  XNOR2_X1  g184(.A(G280), .B(KEYINPUT75), .ZN(G297));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n539), .A2(new_n540), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(new_n607), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n603), .A2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n607), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n489), .A2(new_n471), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT13), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n480), .A2(G123), .ZN(new_n622));
  OR2_X1    g197(.A1(G99), .A2(G2105), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n623), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(G135), .B2(new_n478), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2096), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n621), .A2(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(G2451), .B(G2454), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n632), .B(new_n633), .Z(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2435), .ZN(new_n636));
  XOR2_X1   g211(.A(G2427), .B(G2438), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n634), .B(new_n639), .ZN(new_n640));
  AND2_X1   g215(.A1(new_n640), .A2(G14), .ZN(G401));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  XNOR2_X1  g217(.A(G2072), .B(G2078), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT17), .ZN(new_n644));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n642), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n643), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT76), .Z(new_n649));
  NAND3_X1  g224(.A1(new_n646), .A2(new_n642), .A3(new_n643), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT18), .Z(new_n651));
  INV_X1    g226(.A(new_n644), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n652), .A2(new_n642), .A3(new_n645), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n649), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(G227));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n658), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  AOI22_X1  g239(.A1(new_n662), .A2(KEYINPUT20), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n666), .A2(new_n658), .A3(new_n661), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n665), .B(new_n667), .C1(KEYINPUT20), .C2(new_n662), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT77), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(G229));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n676), .A2(G20), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(KEYINPUT23), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT23), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(G299), .B2(G16), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n678), .B1(new_n680), .B2(new_n677), .ZN(new_n681));
  INV_X1    g256(.A(G1956), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(G2090), .ZN(new_n684));
  AND2_X1   g259(.A1(KEYINPUT78), .A2(G29), .ZN(new_n685));
  NOR2_X1   g260(.A1(KEYINPUT78), .A2(G29), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G35), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G162), .B2(new_n688), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n690), .A2(KEYINPUT87), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(KEYINPUT87), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT86), .B(KEYINPUT29), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(new_n691), .B2(new_n692), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n683), .B1(new_n684), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT89), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G33), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n489), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n702), .A2(new_n469), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT82), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n478), .A2(G139), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n471), .A2(G103), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT25), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n704), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n701), .B1(new_n710), .B2(new_n700), .ZN(new_n711));
  INV_X1    g286(.A(G2072), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n478), .A2(G140), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n480), .A2(G128), .ZN(new_n715));
  NOR2_X1   g290(.A1(G104), .A2(G2105), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(new_n469), .B2(G116), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n714), .B(new_n715), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G29), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n688), .A2(KEYINPUT28), .A3(G26), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(KEYINPUT28), .B1(new_n688), .B2(G26), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(G2067), .Z(new_n724));
  OR2_X1    g299(.A1(G29), .A2(G32), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n478), .A2(G141), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n480), .A2(G129), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n471), .A2(G105), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT26), .Z(new_n730));
  NAND4_X1  g305(.A1(new_n726), .A2(new_n727), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n725), .B1(new_n731), .B2(new_n700), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT27), .B(G1996), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G28), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n626), .A2(new_n687), .B1(new_n700), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n734), .A2(new_n735), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G5), .A2(G16), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G171), .B2(G16), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(G1961), .ZN(new_n742));
  NOR3_X1   g317(.A1(new_n724), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n676), .A2(G19), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n541), .B2(new_n676), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(G1341), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(G1341), .ZN(new_n747));
  INV_X1    g322(.A(G2084), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT83), .B(KEYINPUT24), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G34), .ZN(new_n750));
  OAI22_X1  g325(.A1(new_n476), .A2(new_n700), .B1(new_n687), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n747), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n746), .B(new_n752), .C1(new_n748), .C2(new_n751), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n713), .A2(new_n743), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(G2090), .B1(new_n695), .B2(new_n696), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(KEYINPUT88), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(KEYINPUT88), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT31), .B(G11), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n741), .A2(G1961), .ZN(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  NOR2_X1   g336(.A1(G164), .A2(new_n688), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G27), .B2(new_n688), .ZN(new_n763));
  NAND2_X1  g338(.A1(G168), .A2(G16), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G16), .B2(G21), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT84), .B(G1966), .Z(new_n766));
  OAI221_X1 g341(.A(new_n760), .B1(new_n761), .B2(new_n763), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n676), .A2(G4), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n604), .B2(new_n676), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1348), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n765), .A2(new_n766), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n767), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  AND4_X1   g347(.A1(new_n699), .A2(new_n758), .A3(new_n759), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n676), .A2(G24), .ZN(new_n774));
  INV_X1    g349(.A(G290), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n676), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1986), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT80), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G16), .B2(G23), .ZN(new_n779));
  OR3_X1    g354(.A1(new_n778), .A2(G16), .A3(G23), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n779), .B(new_n780), .C1(G288), .C2(new_n676), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT33), .B(G1976), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n676), .A2(G22), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G166), .B2(new_n676), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G1971), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n783), .A2(new_n784), .A3(new_n787), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n676), .A2(G6), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G305), .B2(G16), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT32), .B(G1981), .Z(new_n791));
  AOI21_X1  g366(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n786), .A2(G1971), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n777), .B1(new_n795), .B2(KEYINPUT34), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT34), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n792), .A2(new_n793), .A3(new_n797), .A4(new_n794), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n688), .A2(G25), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n478), .A2(G131), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n480), .A2(G119), .ZN(new_n801));
  OR2_X1    g376(.A1(G95), .A2(G2105), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n802), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT79), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n799), .B1(new_n805), .B2(new_n688), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT35), .B(G1991), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n806), .B(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n796), .A2(new_n798), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT81), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n811), .A2(new_n812), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n810), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n763), .A2(new_n761), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n796), .A2(new_n813), .A3(new_n798), .A4(new_n809), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n773), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(G150));
  INV_X1    g394(.A(KEYINPUT90), .ZN(new_n820));
  XNOR2_X1  g395(.A(G150), .B(new_n820), .ZN(G311));
  INV_X1    g396(.A(KEYINPUT95), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n603), .A2(new_n611), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT38), .ZN(new_n824));
  OAI21_X1  g399(.A(KEYINPUT94), .B1(new_n541), .B2(KEYINPUT93), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT93), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n613), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n513), .A2(G93), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT91), .B(G55), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n511), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT92), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT92), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n830), .A2(new_n835), .A3(new_n832), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(G80), .A2(G543), .ZN(new_n838));
  INV_X1    g413(.A(G67), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n503), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G651), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n539), .A2(KEYINPUT93), .A3(new_n540), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n837), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n829), .A2(new_n843), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n834), .A2(new_n836), .B1(G651), .B2(new_n840), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n845), .A2(new_n825), .A3(new_n842), .A4(new_n828), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n824), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n822), .B1(new_n849), .B2(KEYINPUT39), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(KEYINPUT95), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT96), .B(G860), .Z(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n850), .A2(new_n852), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n845), .A2(new_n855), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT37), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(G145));
  XNOR2_X1  g436(.A(new_n484), .B(KEYINPUT98), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G160), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n626), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n488), .A2(new_n490), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n491), .A2(new_n495), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n491), .A2(KEYINPUT99), .A3(new_n495), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n718), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n871), .A2(new_n731), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n731), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n710), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(KEYINPUT100), .A3(new_n710), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n874), .B2(new_n710), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n872), .A2(KEYINPUT101), .A3(new_n709), .A4(new_n873), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n619), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT79), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n804), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n804), .A2(new_n886), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n478), .A2(G142), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n480), .A2(G130), .ZN(new_n891));
  OR2_X1    g466(.A1(G106), .A2(G2105), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n892), .B(G2104), .C1(G118), .C2(new_n469), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n805), .A2(new_n894), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n898), .B1(new_n896), .B2(new_n897), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n885), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n889), .A2(new_n895), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n805), .A2(new_n894), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT102), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(new_n619), .A3(new_n899), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n884), .A2(KEYINPUT104), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n900), .A2(new_n885), .A3(new_n901), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n619), .B1(new_n905), .B2(new_n899), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n902), .A2(KEYINPUT103), .A3(new_n906), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n877), .A2(new_n878), .B1(new_n881), .B2(new_n882), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n909), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n879), .A2(new_n883), .B1(new_n906), .B2(new_n902), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n864), .B(new_n908), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n864), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n915), .A2(new_n916), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n915), .A2(new_n916), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n927));
  XNOR2_X1  g502(.A(G288), .B(G303), .ZN(new_n928));
  NAND2_X1  g503(.A1(G305), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(G288), .B(G166), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n930), .A2(new_n586), .A3(new_n585), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n775), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n775), .B1(new_n929), .B2(new_n931), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n927), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n929), .A2(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(G290), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(KEYINPUT106), .A3(new_n932), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(KEYINPUT42), .A3(new_n938), .ZN(new_n939));
  OR3_X1    g514(.A1(new_n933), .A2(KEYINPUT42), .A3(new_n934), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n603), .A2(G299), .ZN(new_n943));
  INV_X1    g518(.A(G299), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n601), .A2(new_n944), .A3(new_n602), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT41), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT41), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n943), .A2(new_n948), .A3(new_n945), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(KEYINPUT105), .A3(new_n949), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n949), .A2(KEYINPUT105), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n847), .B1(G559), .B2(new_n603), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n615), .A2(new_n846), .A3(new_n844), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n946), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n942), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n950), .A2(new_n951), .B1(new_n954), .B2(new_n953), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n961), .A2(KEYINPUT107), .A3(new_n958), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n941), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n956), .A2(new_n942), .A3(new_n959), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT107), .B1(new_n961), .B2(new_n958), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n939), .A2(new_n940), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n963), .A2(G868), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n845), .A2(G868), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(new_n972), .B2(new_n969), .ZN(G295));
  OAI21_X1  g548(.A(new_n970), .B1(new_n972), .B2(new_n969), .ZN(G331));
  XNOR2_X1  g549(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n847), .A2(G171), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n844), .A2(G301), .A3(new_n846), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(G286), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(G168), .A3(new_n977), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(new_n951), .A3(new_n950), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n979), .A2(new_n957), .A3(new_n980), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(new_n938), .A3(new_n935), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n924), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n982), .A2(new_n983), .B1(new_n938), .B2(new_n935), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n975), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n947), .A2(new_n949), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n981), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(KEYINPUT111), .A3(new_n983), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n935), .A2(new_n938), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n983), .A2(KEYINPUT111), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n975), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n993), .A2(new_n924), .A3(new_n984), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n987), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n993), .A2(new_n924), .A3(new_n984), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1000));
  INV_X1    g575(.A(new_n986), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1001), .A2(new_n924), .A3(new_n984), .A4(new_n994), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(KEYINPUT44), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n998), .A2(new_n1003), .ZN(G397));
  NAND2_X1  g579(.A1(new_n868), .A2(new_n869), .ZN(new_n1005));
  INV_X1    g580(.A(new_n865), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1384), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(KEYINPUT45), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT112), .B(G40), .Z(new_n1009));
  OAI211_X1 g584(.A(new_n468), .B(new_n1009), .C1(new_n474), .C2(new_n475), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n718), .B(G2067), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT114), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(G1996), .A3(new_n731), .ZN(new_n1017));
  XOR2_X1   g592(.A(new_n1017), .B(KEYINPUT113), .Z(new_n1018));
  NOR2_X1   g593(.A1(new_n1012), .A2(G1996), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1016), .B(new_n1018), .C1(new_n731), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1022), .A2(new_n808), .A3(new_n805), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n718), .A2(G2067), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1012), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n805), .B(new_n808), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n1013), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1012), .A2(G1986), .A3(G290), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1028), .B(KEYINPUT48), .Z(new_n1029));
  AND3_X1   g604(.A1(new_n1022), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1019), .A2(KEYINPUT46), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1013), .B1(new_n731), .B2(new_n1014), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1019), .A2(KEYINPUT46), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  XOR2_X1   g609(.A(new_n1034), .B(KEYINPUT47), .Z(new_n1035));
  NOR3_X1   g610(.A1(new_n1025), .A2(new_n1030), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1011), .A2(new_n1007), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT116), .B(G8), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G288), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n1040), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT52), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n555), .A2(KEYINPUT71), .A3(new_n518), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT71), .B1(new_n555), .B2(new_n518), .ZN(new_n1048));
  OAI21_X1  g623(.A(G86), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G1981), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n583), .A2(new_n1049), .A3(new_n1050), .A4(new_n572), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT117), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n574), .A2(new_n1053), .A3(new_n1050), .A4(new_n583), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n573), .B1(G86), .B2(new_n513), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n507), .B2(new_n578), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G1981), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(KEYINPUT49), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT118), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1052), .A2(new_n1054), .B1(G1981), .B2(new_n1057), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(KEYINPUT49), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT49), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1039), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1046), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(G303), .A2(G8), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1069), .B(new_n1070), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n491), .A2(KEYINPUT99), .A3(new_n495), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT99), .B1(new_n491), .B2(new_n495), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n488), .B(new_n490), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT50), .ZN(new_n1075));
  INV_X1    g650(.A(G1384), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n496), .A2(new_n1076), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT50), .ZN(new_n1079));
  AND4_X1   g654(.A1(new_n684), .A2(new_n1077), .A3(new_n1011), .A4(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT115), .B(G1971), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT45), .B1(new_n496), .B2(new_n1076), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(new_n1010), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1074), .A2(KEYINPUT45), .A3(new_n1076), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1071), .B(G8), .C1(new_n1080), .C2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1068), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1055), .ZN(new_n1089));
  AOI21_X1  g664(.A(G1976), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1090));
  INV_X1    g665(.A(G288), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1088), .B1(new_n1092), .B2(new_n1039), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1086), .A2(KEYINPUT119), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1075), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n496), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NOR4_X1   g672(.A1(new_n1095), .A2(new_n1097), .A3(G2090), .A4(new_n1010), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1038), .B1(new_n1098), .B2(new_n1085), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1071), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1094), .A2(new_n1101), .ZN(new_n1102));
  AND4_X1   g677(.A1(new_n1062), .A2(new_n1055), .A3(KEYINPUT49), .A4(new_n1058), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1062), .B1(new_n1061), .B2(KEYINPUT49), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1067), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1046), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1099), .A2(KEYINPUT119), .A3(new_n1100), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1102), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n1076), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1011), .B(new_n1109), .C1(new_n1007), .C2(KEYINPUT45), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n766), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1010), .B1(KEYINPUT50), .B2(new_n1078), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(new_n748), .A3(new_n1077), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1038), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(G286), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT120), .B1(new_n1108), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT63), .ZN(new_n1119));
  AOI22_X1  g694(.A1(KEYINPUT119), .A2(new_n1086), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1107), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1122), .A2(new_n1123), .A3(new_n1068), .A4(new_n1116), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1118), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(G8), .B1(new_n1080), .B2(new_n1085), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1117), .B1(new_n1100), .B2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1127), .A2(KEYINPUT63), .A3(new_n1068), .A4(new_n1086), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1093), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1129), .A2(KEYINPUT121), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  AOI211_X1 g706(.A(new_n1131), .B(new_n1093), .C1(new_n1125), .C2(new_n1128), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n1133));
  NAND2_X1  g708(.A1(G299), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(G299), .A2(new_n1133), .A3(KEYINPUT57), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1095), .A2(new_n1010), .ZN(new_n1139));
  AOI21_X1  g714(.A(G1956), .B1(new_n1139), .B2(new_n1096), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT123), .B(KEYINPUT56), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(new_n712), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1083), .A2(new_n1084), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1138), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1011), .B1(new_n1007), .B2(new_n1075), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n682), .B1(new_n1146), .B2(new_n1097), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1147), .A2(new_n1137), .A3(new_n1136), .A4(new_n1143), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT61), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1077), .A2(new_n1011), .A3(new_n1079), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1112), .A2(KEYINPUT124), .A3(new_n1077), .ZN(new_n1153));
  AOI21_X1  g728(.A(G1348), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1037), .A2(G2067), .ZN(new_n1155));
  NOR4_X1   g730(.A1(new_n1154), .A2(KEYINPUT60), .A3(new_n603), .A4(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1149), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(G1348), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT124), .B1(new_n1112), .B2(new_n1077), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1155), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n603), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1154), .A2(new_n604), .A3(new_n1155), .ZN(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT60), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(KEYINPUT125), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1147), .A2(new_n1167), .A3(new_n1143), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1166), .A2(new_n1168), .A3(new_n1138), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1169), .A2(KEYINPUT61), .A3(new_n1148), .ZN(new_n1170));
  XOR2_X1   g745(.A(KEYINPUT58), .B(G1341), .Z(new_n1171));
  NAND2_X1  g746(.A1(new_n1037), .A2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(KEYINPUT126), .B(G1996), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1083), .A2(new_n1084), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n613), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1175), .B(KEYINPUT59), .Z(new_n1176));
  NAND4_X1  g751(.A1(new_n1157), .A2(new_n1165), .A3(new_n1170), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1169), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1148), .B1(new_n1178), .B2(new_n1163), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1181));
  NAND2_X1  g756(.A1(G286), .A2(new_n1038), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(G8), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1182), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(KEYINPUT51), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT51), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1115), .A2(new_n1187), .A3(new_n1182), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1183), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g764(.A(G301), .B(KEYINPUT54), .ZN(new_n1190));
  INV_X1    g765(.A(G1961), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1191), .B1(new_n1160), .B2(new_n1159), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1083), .A2(new_n761), .A3(new_n1084), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT53), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n761), .A2(KEYINPUT53), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1192), .B(new_n1195), .C1(new_n1196), .C2(new_n1110), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1189), .B1(new_n1190), .B2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1122), .A2(KEYINPUT127), .A3(new_n1068), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1108), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(G40), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1008), .A2(new_n1203), .ZN(new_n1204));
  AOI211_X1 g779(.A(new_n476), .B(new_n1196), .C1(new_n1007), .C2(KEYINPUT45), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1190), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1192), .A2(new_n1195), .A3(new_n1206), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n1180), .A2(new_n1198), .A3(new_n1202), .A4(new_n1207), .ZN(new_n1208));
  AOI22_X1  g783(.A1(new_n1114), .A2(G8), .B1(G286), .B2(new_n1038), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1188), .B1(new_n1209), .B2(new_n1187), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1210), .B1(new_n1182), .B2(new_n1181), .ZN(new_n1211));
  AOI21_X1  g786(.A(G301), .B1(new_n1211), .B2(KEYINPUT62), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT62), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1189), .A2(new_n1213), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1212), .A2(new_n1202), .A3(new_n1197), .A4(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1208), .A2(new_n1215), .ZN(new_n1216));
  NOR3_X1   g791(.A1(new_n1130), .A2(new_n1132), .A3(new_n1216), .ZN(new_n1217));
  XOR2_X1   g792(.A(G290), .B(G1986), .Z(new_n1218));
  OAI211_X1 g793(.A(new_n1022), .B(new_n1027), .C1(new_n1012), .C2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1036), .B1(new_n1217), .B2(new_n1219), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g795(.A1(G227), .A2(G401), .ZN(new_n1222));
  AND2_X1   g796(.A1(new_n925), .A2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g797(.A1(G229), .A2(new_n460), .ZN(new_n1224));
  AND3_X1   g798(.A1(new_n1223), .A2(new_n996), .A3(new_n1224), .ZN(G308));
  NAND3_X1  g799(.A1(new_n1223), .A2(new_n996), .A3(new_n1224), .ZN(G225));
endmodule


