//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G183gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT27), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT27), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT28), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT28), .A4(new_n207), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT66), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT27), .B(G183gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT28), .A4(new_n207), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n208), .A2(KEYINPUT65), .A3(new_n209), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n212), .A2(new_n214), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n221), .B1(new_n223), .B2(KEYINPUT26), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT26), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G169gat), .ZN(new_n231));
  INV_X1    g030(.A(G176gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT23), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n233), .A2(new_n235), .A3(new_n236), .A4(new_n220), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT25), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n233), .A2(new_n235), .A3(new_n220), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT24), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n203), .ZN(new_n241));
  NAND2_X1  g040(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(G190gat), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n207), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n238), .B1(new_n239), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n239), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n242), .A2(G190gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n207), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n248), .B1(new_n249), .B2(new_n241), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n247), .A2(new_n250), .A3(KEYINPUT64), .A4(KEYINPUT25), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n219), .A2(new_n230), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n202), .B1(new_n252), .B2(KEYINPUT29), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT22), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT73), .B(G211gat), .ZN(new_n255));
  INV_X1    g054(.A(G218gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G197gat), .B(G204gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(G211gat), .B(G218gat), .Z(new_n260));
  AND2_X1   g059(.A1(new_n260), .A2(KEYINPUT74), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n259), .B(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n251), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n214), .A2(new_n217), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n208), .A2(KEYINPUT65), .A3(new_n209), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT65), .B1(new_n208), .B2(new_n209), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n263), .B1(new_n267), .B2(new_n229), .ZN(new_n268));
  INV_X1    g067(.A(new_n202), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n253), .A2(new_n262), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n262), .B1(new_n253), .B2(new_n270), .ZN(new_n272));
  XNOR2_X1  g071(.A(G8gat), .B(G36gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT75), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT76), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT75), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n273), .B(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT76), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n275), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n280), .B1(new_n275), .B2(new_n279), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NOR3_X1   g083(.A1(new_n271), .A2(new_n272), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT77), .ZN(new_n286));
  NOR3_X1   g085(.A1(new_n281), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n280), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n277), .A2(new_n278), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n274), .A2(KEYINPUT76), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n279), .A3(new_n280), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT77), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n262), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT29), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n269), .B1(new_n268), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n252), .A2(new_n202), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n253), .A2(new_n270), .A3(new_n262), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n294), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT30), .B1(new_n285), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n299), .A2(new_n283), .A3(new_n300), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT30), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT40), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT39), .ZN(new_n308));
  XOR2_X1   g107(.A(G141gat), .B(G148gat), .Z(new_n309));
  INV_X1    g108(.A(G155gat), .ZN(new_n310));
  INV_X1    g109(.A(G162gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(KEYINPUT2), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n309), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G141gat), .B(G148gat), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n313), .B(new_n312), .C1(new_n317), .C2(KEYINPUT2), .ZN(new_n318));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320));
  INV_X1    g119(.A(G113gat), .ZN(new_n321));
  INV_X1    g120(.A(G120gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G113gat), .A2(G120gat), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n319), .A2(new_n320), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n316), .A2(new_n318), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT67), .ZN(new_n327));
  AND2_X1   g126(.A1(G113gat), .A2(G120gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(G113gat), .A2(G120gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n323), .A2(KEYINPUT67), .A3(new_n324), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(new_n331), .A3(new_n320), .ZN(new_n332));
  INV_X1    g131(.A(new_n319), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n332), .A2(KEYINPUT68), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT68), .B1(new_n332), .B2(new_n333), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n326), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n325), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n332), .A2(new_n333), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT68), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n332), .A2(KEYINPUT68), .A3(new_n333), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n338), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n316), .A2(new_n318), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT79), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n325), .B1(new_n334), .B2(new_n335), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT79), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n344), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n337), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G225gat), .A2(G233gat), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n308), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n336), .A2(KEYINPUT4), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n326), .B(new_n354), .C1(new_n334), .C2(new_n335), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(KEYINPUT80), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n344), .B(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n347), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n336), .A2(new_n360), .A3(KEYINPUT4), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n356), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n351), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n352), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n308), .A3(new_n363), .ZN(new_n366));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT0), .ZN(new_n368));
  XNOR2_X1  g167(.A(G57gat), .B(G85gat), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n368), .B(new_n369), .Z(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n307), .B1(new_n365), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n353), .A2(KEYINPUT78), .A3(new_n355), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n363), .B1(new_n358), .B2(new_n347), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n337), .A2(new_n375), .A3(new_n354), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n377), .B(KEYINPUT5), .C1(new_n351), .C2(new_n350), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT5), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n356), .A2(new_n379), .A3(new_n374), .A4(new_n361), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n370), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n352), .A2(new_n364), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n384), .A2(KEYINPUT40), .A3(new_n370), .A4(new_n366), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n306), .A2(new_n372), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G78gat), .B(G106gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT31), .B(G50gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n387), .B(new_n388), .Z(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G228gat), .A2(G233gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n391), .B(KEYINPUT81), .Z(new_n392));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n393), .B1(new_n257), .B2(new_n258), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n394), .A2(new_n260), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n257), .A2(new_n393), .A3(new_n258), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n394), .B2(new_n260), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n296), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n345), .B1(new_n398), .B2(new_n357), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT29), .B1(new_n345), .B2(new_n357), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(new_n262), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n392), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n391), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT3), .B1(new_n262), .B2(new_n296), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n403), .B1(new_n345), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n390), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT83), .B(G22gat), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n402), .A2(new_n405), .A3(new_n390), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n408), .ZN(new_n411));
  INV_X1    g210(.A(new_n409), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n411), .B1(new_n412), .B2(new_n406), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n386), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n378), .A2(new_n370), .A3(new_n380), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n383), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n294), .A2(KEYINPUT38), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n271), .A2(new_n272), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT37), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT37), .B1(new_n271), .B2(new_n272), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n285), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n420), .A2(new_n421), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(new_n284), .A3(new_n423), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT38), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n381), .A2(KEYINPUT6), .A3(new_n382), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n418), .A2(new_n424), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n306), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n417), .A2(new_n416), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n370), .B1(new_n378), .B2(new_n380), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n428), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n410), .A2(new_n413), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n415), .A2(new_n429), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n265), .A2(new_n266), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n214), .A2(new_n217), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n229), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT25), .ZN(new_n441));
  NOR4_X1   g240(.A1(new_n245), .A2(new_n239), .A3(new_n236), .A4(new_n441), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n247), .A2(new_n250), .B1(new_n237), .B2(KEYINPUT25), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT69), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT69), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n446), .B(new_n263), .C1(new_n267), .C2(new_n229), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n347), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(G227gat), .ZN(new_n449));
  INV_X1    g248(.A(G233gat), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n268), .A2(KEYINPUT69), .A3(new_n343), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n448), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT32), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(G15gat), .B(G43gat), .Z(new_n457));
  XNOR2_X1  g256(.A(G71gat), .B(G99gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n454), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n459), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n453), .B(KEYINPUT32), .C1(new_n455), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n452), .ZN(new_n464));
  INV_X1    g263(.A(new_n451), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT34), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(KEYINPUT71), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n463), .A2(new_n472), .ZN(new_n473));
  AOI211_X1 g272(.A(new_n451), .B(new_n471), .C1(new_n448), .C2(new_n452), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n466), .B2(new_n468), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(new_n460), .A3(new_n462), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(KEYINPUT72), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT36), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT72), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n475), .A2(new_n479), .A3(new_n460), .A4(new_n462), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n473), .A2(KEYINPUT36), .A3(new_n476), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n414), .A2(new_n476), .A3(new_n473), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT35), .B1(new_n435), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n477), .A2(new_n480), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n436), .A2(KEYINPUT35), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n306), .B1(new_n418), .B2(new_n428), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n437), .A2(new_n483), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT88), .ZN(new_n491));
  XNOR2_X1  g290(.A(G15gat), .B(G22gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G1gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n492), .A2(new_n493), .A3(G1gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT16), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(G8gat), .ZN(new_n501));
  XOR2_X1   g300(.A(G43gat), .B(G50gat), .Z(new_n502));
  INV_X1    g301(.A(G36gat), .ZN(new_n503));
  AND2_X1   g302(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G29gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n507), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n502), .B1(new_n509), .B2(KEYINPUT15), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(KEYINPUT15), .B2(new_n509), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(KEYINPUT15), .A3(new_n502), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n491), .B1(new_n501), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G8gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n500), .B(new_n515), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n511), .A2(new_n512), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT88), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n513), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n514), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT89), .ZN(new_n521));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n522), .B(KEYINPUT13), .Z(new_n523));
  AND3_X1   g322(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n521), .B1(new_n520), .B2(new_n523), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n513), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n511), .A2(KEYINPUT17), .A3(new_n512), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n516), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(new_n522), .A3(new_n519), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT18), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT86), .B1(new_n526), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G113gat), .B(G141gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT85), .ZN(new_n536));
  XNOR2_X1  g335(.A(G169gat), .B(G197gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT12), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n534), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g342(.A(KEYINPUT86), .B(new_n541), .C1(new_n526), .C2(new_n533), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n490), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G64gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(G57gat), .ZN(new_n548));
  XOR2_X1   g347(.A(KEYINPUT92), .B(G57gat), .Z(new_n549));
  OAI21_X1  g348(.A(new_n548), .B1(new_n549), .B2(new_n547), .ZN(new_n550));
  XNOR2_X1  g349(.A(G71gat), .B(G78gat), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT90), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G57gat), .B(G64gat), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n551), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT91), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT91), .ZN(new_n559));
  AOI211_X1 g358(.A(new_n559), .B(new_n551), .C1(new_n553), .C2(new_n555), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n554), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT21), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G127gat), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n566), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n516), .B1(new_n561), .B2(new_n562), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(G155gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n572), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n577), .B1(new_n572), .B2(new_n573), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n581), .A2(KEYINPUT41), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G134gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(new_n311), .ZN(new_n584));
  NAND2_X1  g383(.A1(G85gat), .A2(G92gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT7), .ZN(new_n586));
  NAND2_X1  g385(.A1(G99gat), .A2(G106gat), .ZN(new_n587));
  INV_X1    g386(.A(G85gat), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  AOI22_X1  g388(.A1(KEYINPUT8), .A2(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(G99gat), .B(G106gat), .Z(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n592), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(new_n586), .A3(new_n590), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n513), .A2(new_n597), .B1(KEYINPUT41), .B2(new_n581), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT93), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n528), .A2(new_n529), .A3(new_n596), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n584), .B1(new_n603), .B2(KEYINPUT94), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n601), .A2(new_n602), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n602), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n605), .A2(KEYINPUT94), .A3(new_n606), .A4(new_n584), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n580), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n558), .ZN(new_n612));
  INV_X1    g411(.A(new_n560), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n593), .A2(new_n615), .A3(new_n595), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n596), .A2(KEYINPUT95), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n614), .A2(new_n554), .A3(new_n616), .A4(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n561), .A2(new_n615), .A3(new_n597), .ZN(new_n619));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  AND2_X1   g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT96), .B(KEYINPUT10), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n627), .B1(new_n618), .B2(new_n619), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n561), .A2(new_n629), .A3(new_n596), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT97), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n620), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n628), .A2(KEYINPUT97), .A3(new_n630), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n626), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n620), .B1(new_n628), .B2(new_n630), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n622), .ZN(new_n636));
  INV_X1    g435(.A(new_n625), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n634), .A2(KEYINPUT98), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT98), .B1(new_n634), .B2(new_n638), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n611), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n546), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n433), .A2(new_n434), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT99), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(new_n495), .ZN(G1324gat));
  INV_X1    g446(.A(new_n643), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n515), .B1(new_n648), .B2(new_n306), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT16), .B(G8gat), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n643), .A2(new_n430), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT42), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(KEYINPUT42), .B2(new_n651), .ZN(G1325gat));
  AOI21_X1  g452(.A(G15gat), .B1(new_n648), .B2(new_n486), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT100), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n481), .A2(G15gat), .A3(new_n482), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n655), .B1(new_n648), .B2(new_n656), .ZN(G1326gat));
  NOR2_X1   g456(.A1(new_n643), .A2(new_n414), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT43), .B(G22gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(G1327gat));
  NOR2_X1   g461(.A1(new_n580), .A2(new_n641), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n608), .A2(new_n609), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT103), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n546), .ZN(new_n667));
  INV_X1    g466(.A(new_n645), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n507), .ZN(new_n669));
  OR3_X1    g468(.A1(new_n667), .A2(KEYINPUT104), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT104), .B1(new_n667), .B2(new_n669), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(KEYINPUT45), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT44), .B1(new_n490), .B2(new_n610), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n664), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n429), .A2(new_n414), .A3(new_n386), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(new_n488), .B2(new_n414), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n435), .A2(KEYINPUT105), .A3(new_n436), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n483), .A2(new_n676), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n489), .A2(new_n485), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n675), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n673), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n543), .A2(new_n544), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(new_n685), .A3(new_n663), .ZN(new_n686));
  OAI21_X1  g485(.A(G29gat), .B1(new_n686), .B2(new_n645), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT45), .B1(new_n670), .B2(new_n671), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n688), .A2(new_n689), .ZN(G1328gat));
  NOR3_X1   g489(.A1(new_n667), .A2(G36gat), .A3(new_n430), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT46), .ZN(new_n692));
  OAI21_X1  g491(.A(G36gat), .B1(new_n686), .B2(new_n430), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(G1329gat));
  INV_X1    g493(.A(new_n486), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n667), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n481), .A2(G43gat), .A3(new_n482), .ZN(new_n697));
  OAI22_X1  g496(.A1(new_n696), .A2(G43gat), .B1(new_n686), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g498(.A(G50gat), .B1(new_n686), .B2(new_n414), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n414), .A2(G50gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n666), .A2(new_n546), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT106), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT48), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1331gat));
  AND2_X1   g504(.A1(new_n679), .A2(new_n678), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n429), .A2(new_n415), .B1(new_n481), .B2(new_n482), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n706), .A2(new_n707), .B1(new_n485), .B2(new_n489), .ZN(new_n708));
  INV_X1    g507(.A(new_n641), .ZN(new_n709));
  NOR4_X1   g508(.A1(new_n708), .A2(new_n685), .A3(new_n611), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n668), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(new_n549), .ZN(G1332gat));
  XOR2_X1   g511(.A(new_n306), .B(KEYINPUT107), .Z(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT49), .B(G64gat), .Z(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(new_n714), .B2(new_n716), .ZN(G1333gat));
  XNOR2_X1  g516(.A(new_n486), .B(KEYINPUT108), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(G71gat), .B1(new_n710), .B2(new_n719), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n481), .A2(G71gat), .A3(new_n482), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n710), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1334gat));
  NAND2_X1  g523(.A1(new_n710), .A2(new_n436), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g525(.A1(new_n709), .A2(new_n685), .A3(new_n580), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n673), .B2(new_n683), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G85gat), .B1(new_n730), .B2(new_n645), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n578), .A2(new_n579), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n664), .A2(new_n733), .A3(new_n545), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n708), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n680), .A2(new_n681), .ZN(new_n736));
  INV_X1    g535(.A(new_n734), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n736), .A2(KEYINPUT51), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n709), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n739), .A2(new_n588), .A3(new_n668), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n731), .A2(new_n740), .ZN(G1336gat));
  INV_X1    g540(.A(KEYINPUT114), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n589), .B1(new_n729), .B2(new_n713), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n641), .A2(new_n713), .A3(new_n589), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT111), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT51), .B1(new_n736), .B2(new_n737), .ZN(new_n747));
  AOI211_X1 g546(.A(new_n732), .B(new_n734), .C1(new_n680), .C2(new_n681), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n743), .A2(new_n752), .A3(KEYINPUT113), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n735), .A2(new_n738), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n750), .B1(new_n755), .B2(new_n746), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n435), .A2(new_n436), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n483), .A2(new_n757), .A3(new_n676), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n681), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n674), .B1(new_n759), .B2(new_n664), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n713), .B(new_n727), .C1(new_n760), .C2(new_n682), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G92gat), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n754), .B1(new_n756), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n753), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765));
  INV_X1    g564(.A(new_n749), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n306), .B(new_n727), .C1(new_n760), .C2(new_n682), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G92gat), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n767), .A2(KEYINPUT110), .A3(G92gat), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n765), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n742), .B1(new_n764), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n768), .A2(new_n769), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(new_n749), .A3(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT52), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT113), .B1(new_n743), .B2(new_n752), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n756), .A2(new_n754), .A3(new_n762), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(KEYINPUT114), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n773), .A2(new_n780), .ZN(G1337gat));
  INV_X1    g580(.A(G99gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n729), .A2(new_n481), .A3(new_n482), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n784), .B2(new_n783), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n739), .A2(new_n782), .A3(new_n486), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(G1338gat));
  INV_X1    g587(.A(G106gat), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n789), .B1(new_n729), .B2(new_n436), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n791), .B2(KEYINPUT53), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n739), .A2(new_n789), .A3(new_n436), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n794), .B(new_n795), .ZN(G1339gat));
  NOR3_X1   g595(.A1(new_n611), .A2(new_n685), .A3(new_n641), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n526), .A2(new_n533), .A3(new_n542), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n520), .A2(new_n523), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n522), .B1(new_n530), .B2(new_n519), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n540), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g602(.A(KEYINPUT117), .B(new_n540), .C1(new_n799), .C2(new_n800), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n798), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n639), .B2(new_n640), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n637), .B1(new_n635), .B2(KEYINPUT54), .ZN(new_n808));
  OR3_X1    g607(.A1(new_n628), .A2(KEYINPUT97), .A3(new_n630), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(new_n620), .A3(new_n631), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n628), .A2(new_n630), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n812), .B2(new_n621), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n808), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n543), .B(new_n544), .C1(KEYINPUT55), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n810), .A2(new_n813), .ZN(new_n816));
  INV_X1    g615(.A(new_n808), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n634), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n807), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n610), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n814), .A2(KEYINPUT55), .B1(new_n810), .B2(new_n626), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n818), .A2(new_n819), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n664), .A2(new_n806), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n797), .B1(new_n826), .B2(new_n733), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n827), .A2(new_n484), .A3(new_n645), .ZN(new_n828));
  INV_X1    g627(.A(new_n713), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830), .B2(new_n685), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n827), .A2(new_n436), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n832), .A2(new_n486), .A3(new_n668), .A4(new_n829), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n833), .A2(new_n321), .A3(new_n545), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n831), .A2(new_n834), .ZN(G1340gat));
  NAND3_X1  g634(.A1(new_n830), .A2(new_n322), .A3(new_n641), .ZN(new_n836));
  OAI21_X1  g635(.A(G120gat), .B1(new_n833), .B2(new_n709), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(KEYINPUT118), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n837), .A2(KEYINPUT118), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(G1341gat));
  NAND3_X1  g639(.A1(new_n830), .A2(new_n566), .A3(new_n580), .ZN(new_n841));
  OAI21_X1  g640(.A(G127gat), .B1(new_n833), .B2(new_n733), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(G1342gat));
  NAND2_X1  g642(.A1(new_n664), .A2(new_n430), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(G134gat), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n846), .A2(KEYINPUT56), .ZN(new_n847));
  OAI21_X1  g646(.A(G134gat), .B1(new_n833), .B2(new_n610), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(KEYINPUT56), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(G1343gat));
  AND3_X1   g649(.A1(new_n668), .A2(new_n483), .A3(new_n829), .ZN(new_n851));
  INV_X1    g650(.A(G141gat), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n545), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n414), .A2(new_n855), .ZN(new_n856));
  AND4_X1   g655(.A1(new_n664), .A2(new_n806), .A3(new_n823), .A4(new_n824), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n822), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n685), .A2(new_n823), .A3(new_n824), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n664), .B1(new_n860), .B2(new_n807), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT120), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n580), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n854), .B(new_n856), .C1(new_n863), .C2(new_n797), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n733), .B1(new_n861), .B2(new_n857), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n642), .A2(new_n545), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n414), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT119), .B1(new_n867), .B2(KEYINPUT57), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n869), .B(new_n855), .C1(new_n827), .C2(new_n414), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n864), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n825), .B1(new_n861), .B2(KEYINPUT120), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n822), .A2(new_n858), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n733), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n866), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n854), .B1(new_n875), .B2(new_n856), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n851), .B(new_n853), .C1(new_n871), .C2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n827), .A2(new_n645), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n414), .B1(new_n481), .B2(new_n482), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n829), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n852), .B1(new_n880), .B2(new_n545), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT58), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n877), .A2(KEYINPUT58), .A3(new_n881), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1344gat));
  OAI211_X1 g685(.A(new_n641), .B(new_n851), .C1(new_n871), .C2(new_n876), .ZN(new_n887));
  INV_X1    g686(.A(G148gat), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(KEYINPUT59), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n867), .A2(KEYINPUT57), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n827), .A2(new_n855), .A3(new_n414), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n851), .A2(new_n641), .ZN(new_n894));
  OAI21_X1  g693(.A(G148gat), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT59), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n880), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n888), .A3(new_n641), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1345gat));
  OAI21_X1  g699(.A(new_n851), .B1(new_n871), .B2(new_n876), .ZN(new_n901));
  OAI21_X1  g700(.A(G155gat), .B1(new_n901), .B2(new_n733), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n898), .A2(new_n310), .A3(new_n580), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1346gat));
  OAI21_X1  g703(.A(G162gat), .B1(new_n901), .B2(new_n610), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n844), .A2(G162gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n878), .A2(new_n879), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1347gat));
  NOR2_X1   g707(.A1(new_n827), .A2(new_n668), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n829), .A2(new_n484), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n231), .B1(new_n911), .B2(new_n545), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n645), .A2(new_n306), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT122), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n914), .A2(new_n719), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n832), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n685), .A2(G169gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n912), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  XOR2_X1   g717(.A(new_n918), .B(KEYINPUT123), .Z(G1348gat));
  OAI21_X1  g718(.A(G176gat), .B1(new_n916), .B2(new_n709), .ZN(new_n920));
  INV_X1    g719(.A(new_n911), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n232), .A3(new_n641), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1349gat));
  OAI21_X1  g722(.A(G183gat), .B1(new_n916), .B2(new_n733), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n580), .A2(new_n215), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n910), .A3(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n924), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g730(.A1(new_n921), .A2(new_n207), .A3(new_n664), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT125), .ZN(new_n933));
  OAI21_X1  g732(.A(G190gat), .B1(new_n916), .B2(new_n610), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n933), .A2(new_n936), .A3(new_n937), .ZN(G1351gat));
  NAND2_X1  g737(.A1(new_n879), .A2(new_n713), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT126), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n909), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n685), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n914), .A2(new_n483), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT127), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n914), .A2(new_n946), .A3(new_n483), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n893), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n685), .A2(G197gat), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n943), .B1(new_n948), .B2(new_n949), .ZN(G1352gat));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n641), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G204gat), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n941), .A2(G204gat), .A3(new_n709), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT62), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n942), .A2(new_n255), .A3(new_n580), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n945), .A2(new_n947), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n957), .B(new_n580), .C1(new_n891), .C2(new_n892), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(G1354gat));
  NAND3_X1  g760(.A1(new_n942), .A2(new_n256), .A3(new_n664), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n948), .A2(new_n664), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n963), .B2(new_n256), .ZN(G1355gat));
endmodule


