//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G140), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  AND2_X1   g003(.A1(new_n189), .A2(G227), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n193), .A2(G143), .ZN(new_n199));
  AOI22_X1  g013(.A1(new_n197), .A2(new_n198), .B1(KEYINPUT1), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n194), .A2(new_n196), .A3(new_n201), .A4(G128), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT79), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(G143), .B(G146), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n205), .A2(KEYINPUT79), .A3(new_n201), .A4(G128), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n200), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n208));
  INV_X1    g022(.A(G104), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G107), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n208), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT77), .B1(new_n213), .B2(G104), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT77), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n209), .A3(G107), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G101), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(G104), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n212), .A2(new_n217), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n209), .A2(G107), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n222), .A3(KEYINPUT78), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n223), .B(G101), .C1(KEYINPUT78), .C2(new_n222), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n207), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n200), .A2(new_n202), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n221), .A2(new_n224), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n228), .A3(KEYINPUT81), .ZN(new_n229));
  INV_X1    g043(.A(G134), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G137), .ZN(new_n231));
  INV_X1    g045(.A(G137), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT65), .B1(new_n232), .B2(G134), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n231), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n236), .B(new_n234), .C1(new_n230), .C2(G137), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(G131), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n236), .B1(new_n230), .B2(G137), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT11), .ZN(new_n241));
  INV_X1    g055(.A(G131), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n241), .A2(new_n242), .A3(new_n237), .A4(new_n231), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT81), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n226), .A2(new_n227), .A3(new_n245), .ZN(new_n246));
  XOR2_X1   g060(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n247));
  NAND4_X1  g061(.A1(new_n229), .A2(new_n244), .A3(new_n246), .A4(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n249));
  INV_X1    g063(.A(new_n243), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n232), .A2(G134), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n251), .B1(new_n240), .B2(KEYINPUT11), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n242), .B1(new_n252), .B2(new_n237), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n249), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n239), .A2(KEYINPUT69), .A3(new_n243), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n229), .A2(new_n256), .A3(new_n246), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT82), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT12), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n258), .B1(new_n257), .B2(new_n259), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n248), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n256), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n212), .A2(new_n217), .A3(new_n220), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G101), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n205), .A2(KEYINPUT0), .A3(G128), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT0), .B(G128), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n267), .B1(new_n205), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n264), .A2(new_n271), .A3(G101), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n266), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT10), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n225), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n227), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n200), .A2(new_n202), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(KEYINPUT10), .A3(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n263), .A2(new_n273), .A3(new_n275), .A4(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n192), .B1(new_n262), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n273), .A2(new_n275), .A3(new_n278), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n256), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(new_n192), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT83), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n284), .B2(new_n283), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n187), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G469), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT84), .ZN(new_n289));
  INV_X1    g103(.A(new_n283), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n262), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n192), .B1(new_n282), .B2(new_n279), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(G902), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G469), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n289), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n292), .B1(new_n262), .B2(new_n290), .ZN(new_n297));
  NOR4_X1   g111(.A1(new_n297), .A2(KEYINPUT84), .A3(G469), .A4(G902), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n288), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT91), .B(G475), .Z(new_n300));
  INV_X1    g114(.A(G237), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(new_n189), .A3(G214), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(G143), .ZN(new_n303));
  NAND2_X1  g117(.A1(KEYINPUT18), .A2(G131), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n303), .B(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(G125), .B(G140), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n306), .A2(new_n193), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G125), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(KEYINPUT75), .A3(G140), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n307), .B1(new_n313), .B2(G146), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n305), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n309), .A2(KEYINPUT16), .A3(new_n311), .ZN(new_n316));
  OR2_X1    g130(.A1(new_n310), .A2(G140), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT16), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n193), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n316), .A2(new_n193), .A3(new_n319), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n302), .B(new_n195), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT17), .A3(G131), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT88), .B1(new_n323), .B2(G131), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT88), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n303), .A2(new_n327), .A3(new_n242), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT17), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n323), .A2(G131), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n326), .A2(new_n328), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n315), .B1(new_n325), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G113), .B(G122), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(new_n209), .ZN(new_n334));
  XOR2_X1   g148(.A(new_n334), .B(KEYINPUT90), .Z(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n332), .B2(new_n334), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n300), .B1(new_n337), .B2(new_n187), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT89), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n312), .A2(KEYINPUT19), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(KEYINPUT19), .B2(new_n306), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n320), .B1(new_n342), .B2(new_n193), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n326), .A2(new_n328), .A3(new_n330), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n315), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n340), .B1(new_n345), .B2(new_n334), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n193), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(new_n344), .A3(new_n321), .ZN(new_n348));
  INV_X1    g162(.A(new_n315), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n334), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(KEYINPUT89), .A3(new_n351), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n346), .A2(new_n352), .B1(new_n332), .B2(new_n335), .ZN(new_n353));
  NOR2_X1   g167(.A1(G475), .A2(G902), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n353), .A2(KEYINPUT20), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT20), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT89), .B1(new_n350), .B2(new_n351), .ZN(new_n358));
  AOI211_X1 g172(.A(new_n340), .B(new_n334), .C1(new_n348), .C2(new_n349), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n336), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n357), .B1(new_n360), .B2(new_n354), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n339), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G478), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(KEYINPUT15), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT9), .B(G234), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(G217), .A3(new_n189), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  OR2_X1    g182(.A1(KEYINPUT67), .A2(G116), .ZN(new_n369));
  NAND2_X1  g183(.A1(KEYINPUT67), .A2(G116), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G122), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G116), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(G122), .ZN(new_n375));
  OAI21_X1  g189(.A(G107), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(KEYINPUT67), .B(G116), .Z(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G122), .ZN(new_n378));
  INV_X1    g192(.A(new_n375), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n213), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT92), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n376), .A2(new_n380), .A3(KEYINPUT92), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT13), .B1(new_n195), .B2(G128), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n198), .B2(G143), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n386), .A2(KEYINPUT93), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT93), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n198), .A2(G143), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n388), .B1(new_n389), .B2(KEYINPUT13), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n230), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G128), .B(G143), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n387), .A2(new_n391), .B1(new_n230), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n383), .A2(new_n384), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n392), .B(G134), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n395), .A2(KEYINPUT94), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n213), .B1(new_n373), .B2(KEYINPUT14), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n378), .A2(new_n379), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n397), .B1(new_n398), .B2(KEYINPUT14), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(KEYINPUT94), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n396), .A2(new_n399), .A3(new_n380), .A4(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n368), .B1(new_n394), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n394), .A2(new_n401), .A3(new_n368), .ZN(new_n404));
  AOI21_X1  g218(.A(G902), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(KEYINPUT95), .ZN(new_n406));
  INV_X1    g220(.A(new_n404), .ZN(new_n407));
  OAI211_X1 g221(.A(KEYINPUT95), .B(new_n187), .C1(new_n407), .C2(new_n402), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n364), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  OAI22_X1  g224(.A1(new_n405), .A2(KEYINPUT95), .B1(KEYINPUT15), .B2(new_n363), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n189), .A2(G952), .ZN(new_n413));
  INV_X1    g227(.A(G234), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n413), .B1(new_n414), .B2(new_n301), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AOI211_X1 g230(.A(new_n187), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT21), .B(G898), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n362), .A2(new_n412), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G221), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n366), .B2(new_n187), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(G214), .B1(G237), .B2(G902), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G210), .B1(G237), .B2(G902), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n277), .A2(new_n310), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n310), .B2(new_n269), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n189), .A2(G224), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n428), .B1(KEYINPUT7), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT7), .B1(new_n429), .B2(KEYINPUT86), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(KEYINPUT86), .B2(new_n429), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n428), .A2(KEYINPUT87), .A3(new_n432), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n430), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT5), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n377), .A2(G119), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n374), .A2(G119), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT68), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n369), .A2(new_n441), .A3(G119), .A4(new_n370), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n438), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n438), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G113), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n443), .A2(new_n444), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT2), .B(G113), .ZN(new_n450));
  OAI221_X1 g264(.A(new_n227), .B1(new_n445), .B2(new_n447), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G110), .B(G122), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT8), .ZN(new_n453));
  INV_X1    g267(.A(new_n445), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n447), .B(KEYINPUT85), .Z(new_n455));
  INV_X1    g269(.A(new_n450), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n454), .A2(new_n455), .B1(new_n448), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n451), .B(new_n453), .C1(new_n227), .C2(new_n457), .ZN(new_n458));
  OAI221_X1 g272(.A(new_n276), .B1(new_n445), .B2(new_n447), .C1(new_n449), .C2(new_n450), .ZN(new_n459));
  INV_X1    g273(.A(G119), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n371), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n442), .ZN(new_n462));
  OAI211_X1 g276(.A(KEYINPUT66), .B(new_n444), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n456), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n443), .A2(KEYINPUT66), .A3(new_n444), .A4(new_n450), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n266), .A3(new_n272), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n459), .A2(new_n467), .A3(new_n452), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n437), .A2(new_n458), .A3(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n469), .A2(new_n187), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n459), .A2(new_n467), .ZN(new_n471));
  INV_X1    g285(.A(new_n452), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(KEYINPUT6), .A3(new_n468), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT6), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n471), .A2(new_n475), .A3(new_n472), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n428), .B(new_n429), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n426), .B1(new_n470), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n470), .A2(new_n478), .A3(new_n426), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n425), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n299), .A2(new_n420), .A3(new_n423), .A4(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT96), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n460), .A2(G128), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n198), .A2(G119), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT24), .B(G110), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G110), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n486), .A2(KEYINPUT23), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n487), .A2(KEYINPUT74), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n492), .B(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n322), .ZN(new_n495));
  OAI221_X1 g309(.A(new_n490), .B1(new_n491), .B2(new_n494), .C1(new_n495), .C2(new_n320), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n491), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n488), .A2(new_n489), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n307), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n321), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT22), .B(G137), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n421), .A2(new_n414), .A3(G953), .ZN(new_n503));
  XOR2_X1   g317(.A(new_n502), .B(new_n503), .Z(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n496), .A2(new_n500), .A3(new_n504), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n187), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT25), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G217), .B1(new_n414), .B2(G902), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT73), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(G902), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n506), .A2(new_n507), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(G472), .A2(G902), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n239), .A2(KEYINPUT69), .A3(new_n243), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT69), .B1(new_n239), .B2(new_n243), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n270), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n230), .A2(G137), .ZN(new_n521));
  OAI21_X1  g335(.A(G131), .B1(new_n521), .B2(new_n251), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT70), .B1(new_n243), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n243), .A2(KEYINPUT70), .A3(new_n522), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n277), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n520), .A2(KEYINPUT30), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n243), .A2(new_n522), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n226), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n269), .B1(new_n239), .B2(new_n243), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n527), .A2(new_n466), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n466), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n520), .A3(new_n526), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n301), .A2(new_n189), .A3(G210), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT27), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT26), .B(G101), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n533), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT31), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n533), .A2(KEYINPUT31), .A3(new_n535), .A4(new_n539), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n269), .B1(new_n254), .B2(new_n255), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n243), .A2(KEYINPUT70), .A3(new_n522), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n546), .A2(new_n523), .A3(new_n226), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n545), .A2(new_n547), .A3(new_n466), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n530), .A2(new_n531), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n534), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT28), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT71), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n548), .B2(KEYINPUT28), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT28), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n535), .A2(KEYINPUT71), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n551), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n539), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT72), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n544), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n559), .B1(new_n544), .B2(new_n558), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n517), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT32), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT32), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n564), .B(new_n517), .C1(new_n560), .C2(new_n561), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT29), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n533), .A2(new_n535), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n557), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n567), .B(new_n569), .C1(new_n556), .C2(new_n557), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n553), .A2(new_n555), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n466), .B1(new_n545), .B2(new_n547), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n535), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n571), .B1(KEYINPUT28), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n557), .A2(new_n567), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n570), .A2(new_n187), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(G472), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n516), .B1(new_n566), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n257), .A2(new_n259), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT82), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n283), .B1(new_n583), .B2(new_n248), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n295), .B(new_n187), .C1(new_n584), .C2(new_n292), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT84), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n294), .A2(new_n289), .A3(new_n295), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n422), .B1(new_n588), .B2(new_n288), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n589), .A2(KEYINPUT96), .A3(new_n482), .A4(new_n420), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n485), .A2(new_n579), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  OAI21_X1  g406(.A(new_n187), .B1(new_n560), .B2(new_n561), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G472), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n562), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n299), .A2(new_n423), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n595), .A2(new_n596), .A3(new_n516), .ZN(new_n597));
  INV_X1    g411(.A(new_n419), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n482), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n363), .A2(new_n187), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n405), .B2(new_n363), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n403), .A2(new_n404), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT98), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n403), .A2(new_n606), .A3(KEYINPUT33), .A4(new_n404), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n604), .B1(new_n407), .B2(new_n402), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT97), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n603), .A2(new_n611), .A3(new_n604), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n602), .B1(new_n614), .B2(G478), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n362), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n599), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n597), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT34), .B(G104), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  OAI21_X1  g434(.A(KEYINPUT20), .B1(new_n353), .B2(new_n355), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n360), .A2(new_n357), .A3(new_n354), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n361), .A2(KEYINPUT99), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n339), .A3(new_n412), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(new_n599), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n597), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NOR2_X1   g446(.A1(new_n505), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n501), .B(new_n633), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n510), .A2(new_n512), .B1(new_n514), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n594), .A2(new_n562), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n485), .A2(new_n590), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT37), .B(G110), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT100), .B(KEYINPUT101), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G12));
  AOI22_X1  g457(.A1(new_n563), .A2(new_n565), .B1(G472), .B2(new_n577), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n299), .A2(new_n423), .A3(new_n482), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n412), .A2(new_n339), .ZN(new_n647));
  INV_X1    g461(.A(G900), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n417), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n415), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR4_X1   g465(.A1(new_n647), .A2(new_n626), .A3(new_n635), .A4(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n646), .A2(KEYINPUT102), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n544), .A2(new_n558), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT72), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n544), .A2(new_n558), .A3(new_n559), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n564), .B1(new_n657), .B2(new_n517), .ZN(new_n658));
  INV_X1    g472(.A(new_n565), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n578), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n586), .A2(new_n587), .B1(G469), .B2(new_n287), .ZN(new_n661));
  INV_X1    g475(.A(new_n481), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n424), .B1(new_n662), .B2(new_n479), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n661), .A2(new_n663), .A3(new_n422), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n660), .A2(new_n664), .A3(new_n652), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n653), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  INV_X1    g483(.A(new_n566), .ZN(new_n670));
  INV_X1    g484(.A(G472), .ZN(new_n671));
  INV_X1    g485(.A(new_n573), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n540), .B1(new_n672), .B2(new_n539), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n671), .B1(new_n673), .B2(new_n187), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n480), .A2(new_n481), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n676), .B(KEYINPUT38), .Z(new_n677));
  AOI21_X1  g491(.A(new_n425), .B1(new_n410), .B2(new_n411), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n362), .ZN(new_n679));
  NOR4_X1   g493(.A1(new_n675), .A2(new_n636), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n680), .A2(KEYINPUT103), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(KEYINPUT103), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n650), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n589), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(KEYINPUT40), .Z(new_n686));
  NAND3_X1  g500(.A1(new_n681), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G143), .ZN(G45));
  NAND4_X1  g502(.A1(new_n636), .A2(new_n615), .A3(new_n362), .A4(new_n650), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n660), .A2(new_n664), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT105), .B(G146), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G48));
  OAI21_X1  g507(.A(G469), .B1(new_n297), .B2(G902), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n423), .B(new_n694), .C1(new_n296), .C2(new_n298), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n588), .A2(KEYINPUT106), .A3(new_n423), .A4(new_n694), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n579), .A3(new_n617), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  INV_X1    g516(.A(new_n516), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n660), .A2(new_n703), .A3(new_n697), .A4(new_n698), .ZN(new_n704));
  INV_X1    g518(.A(new_n629), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT107), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n699), .A2(new_n579), .A3(new_n707), .A4(new_n629), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  AND3_X1   g524(.A1(new_n697), .A2(new_n482), .A3(new_n698), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n420), .A2(new_n636), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n644), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  OAI21_X1  g529(.A(new_n544), .B1(new_n574), .B2(new_n539), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n517), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(G902), .B1(new_n655), .B2(new_n656), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT108), .B1(new_n719), .B2(new_n671), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n593), .A2(new_n721), .A3(G472), .ZN(new_n722));
  AOI211_X1 g536(.A(new_n516), .B(new_n718), .C1(new_n720), .C2(new_n722), .ZN(new_n723));
  AND4_X1   g537(.A1(new_n676), .A2(new_n362), .A3(new_n598), .A4(new_n678), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n697), .A2(new_n698), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  NAND2_X1  g541(.A1(new_n720), .A2(new_n722), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n690), .A3(new_n717), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n697), .A2(new_n482), .A3(new_n698), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT109), .B(G125), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G27));
  NAND2_X1  g547(.A1(new_n566), .A2(KEYINPUT110), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n563), .A2(new_n735), .A3(new_n565), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n734), .A2(new_n578), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n703), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n676), .A2(new_n425), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n589), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n615), .A2(new_n362), .A3(new_n650), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT42), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n740), .A2(new_n644), .A3(new_n516), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT42), .ZN(new_n746));
  INV_X1    g560(.A(new_n741), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  NOR2_X1   g564(.A1(new_n628), .A2(new_n651), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n745), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  NOR2_X1   g567(.A1(new_n280), .A2(new_n286), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n754), .A2(KEYINPUT45), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(KEYINPUT45), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(G469), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(G469), .A2(G902), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n757), .A2(KEYINPUT46), .A3(new_n758), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n588), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n423), .A3(new_n684), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n338), .B1(new_n621), .B2(new_n622), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n615), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n767), .B1(KEYINPUT111), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n769), .A2(KEYINPUT112), .A3(new_n771), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n635), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT44), .B1(new_n776), .B2(new_n595), .ZN(new_n777));
  INV_X1    g591(.A(new_n739), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n776), .A2(KEYINPUT44), .A3(new_n595), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(KEYINPUT113), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(KEYINPUT113), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n765), .B(new_n779), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  NAND2_X1  g598(.A1(new_n763), .A2(new_n423), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n763), .A2(KEYINPUT47), .A3(new_n423), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n644), .A2(new_n516), .A3(new_n747), .A4(new_n739), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT114), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n793));
  AOI211_X1 g607(.A(new_n793), .B(new_n790), .C1(new_n787), .C2(new_n788), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  XOR2_X1   g609(.A(KEYINPUT115), .B(G140), .Z(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(G42));
  NOR4_X1   g611(.A1(new_n767), .A2(new_n516), .A3(new_n422), .A4(new_n425), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n677), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT49), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n588), .A2(new_n694), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n799), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n803), .B(new_n675), .C1(new_n800), .C2(new_n802), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n699), .A2(new_n425), .A3(new_n677), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT119), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n772), .A2(new_n416), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n808), .A2(new_n723), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g624(.A(new_n810), .B(KEYINPUT50), .Z(new_n811));
  NOR2_X1   g625(.A1(new_n801), .A2(new_n423), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n739), .B(new_n809), .C1(new_n789), .C2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n699), .A2(new_n739), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n670), .A2(new_n516), .A3(new_n415), .A4(new_n674), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n615), .A2(new_n362), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n817), .A2(KEYINPUT120), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(KEYINPUT120), .ZN(new_n819));
  AOI211_X1 g633(.A(new_n635), .B(new_n718), .C1(new_n720), .C2(new_n722), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n814), .A2(new_n808), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n818), .A2(new_n819), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n811), .A2(new_n813), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n814), .A2(new_n815), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n413), .B1(new_n828), .B2(new_n616), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n821), .A2(new_n738), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT48), .ZN(new_n831));
  AOI211_X1 g645(.A(new_n829), .B(new_n831), .C1(new_n711), .C2(new_n809), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n826), .A2(new_n827), .A3(new_n832), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n412), .A2(new_n338), .A3(new_n651), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n627), .A3(new_n636), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n740), .A2(new_n644), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n742), .B2(new_n820), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n744), .A2(new_n748), .A3(new_n752), .A4(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n726), .A2(new_n700), .A3(new_n714), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n596), .A2(new_n516), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n766), .A2(new_n412), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n841), .A2(KEYINPUT116), .B1(new_n615), .B2(new_n362), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(KEYINPUT116), .B2(new_n841), .ZN(new_n843));
  INV_X1    g657(.A(new_n599), .ZN(new_n844));
  INV_X1    g658(.A(new_n595), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n840), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n591), .A2(new_n639), .A3(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n839), .A2(new_n709), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n691), .B1(new_n729), .B2(new_n730), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n667), .B2(new_n653), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n679), .B1(new_n480), .B2(new_n481), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n589), .A2(new_n851), .A3(new_n635), .A4(new_n650), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n675), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT52), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n849), .ZN(new_n855));
  AND4_X1   g669(.A1(KEYINPUT52), .A2(new_n668), .A3(new_n855), .A4(new_n853), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n838), .B(new_n848), .C1(new_n854), .C2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n857), .B(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n860), .A3(KEYINPUT54), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n857), .A2(new_n858), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n847), .A2(KEYINPUT53), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n854), .B2(new_n856), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n839), .A2(KEYINPUT118), .A3(new_n709), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT118), .B1(new_n839), .B2(new_n709), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n838), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n862), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n861), .B1(KEYINPUT54), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n860), .B1(new_n859), .B2(KEYINPUT54), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n833), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(G952), .A2(G953), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n804), .B1(new_n873), .B2(new_n874), .ZN(G75));
  NOR2_X1   g689(.A1(new_n189), .A2(G952), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n744), .A2(new_n748), .A3(new_n837), .A4(new_n752), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n706), .A2(new_n708), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n726), .A2(new_n700), .A3(new_n714), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n878), .B1(new_n882), .B2(new_n866), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n668), .A2(new_n855), .A3(new_n853), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT52), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n850), .A2(KEYINPUT52), .A3(new_n853), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n863), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n858), .A2(new_n857), .B1(new_n883), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n187), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT56), .B1(new_n890), .B2(G210), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n474), .A2(new_n476), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n477), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n877), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n890), .A2(KEYINPUT121), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n889), .B2(new_n187), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n426), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n894), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n895), .B1(new_n901), .B2(new_n903), .ZN(G51));
  XNOR2_X1  g718(.A(new_n870), .B(KEYINPUT54), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n758), .B(KEYINPUT57), .Z(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n292), .B2(new_n584), .ZN(new_n908));
  INV_X1    g722(.A(new_n757), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n899), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n876), .B1(new_n908), .B2(new_n910), .ZN(G54));
  NAND4_X1  g725(.A1(new_n896), .A2(KEYINPUT58), .A3(G475), .A4(new_n898), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n912), .A2(new_n353), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n353), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n876), .ZN(G60));
  XNOR2_X1  g729(.A(new_n600), .B(KEYINPUT59), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n905), .A2(new_n613), .A3(new_n608), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n877), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n917), .B1(new_n871), .B2(new_n872), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n919), .B1(new_n920), .B2(new_n614), .ZN(G63));
  XNOR2_X1  g735(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n922));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  OAI21_X1  g738(.A(KEYINPUT123), .B1(new_n889), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n506), .A2(new_n507), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n927));
  INV_X1    g741(.A(new_n924), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n869), .A2(new_n865), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n839), .A2(new_n847), .A3(new_n709), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n886), .B2(new_n887), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT53), .B1(new_n931), .B2(new_n838), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n927), .B(new_n928), .C1(new_n929), .C2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n925), .A2(new_n926), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n934), .A2(KEYINPUT124), .A3(new_n877), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n925), .A2(new_n933), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n634), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT124), .B1(new_n934), .B2(new_n877), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n922), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n937), .A2(KEYINPUT61), .A3(new_n877), .A4(new_n934), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(G66));
  INV_X1    g756(.A(G224), .ZN(new_n943));
  OAI21_X1  g757(.A(G953), .B1(new_n418), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n848), .B2(G953), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n892), .B1(G898), .B2(new_n189), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G69));
  NAND2_X1  g761(.A1(new_n527), .A2(new_n532), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(new_n342), .Z(new_n949));
  XNOR2_X1  g763(.A(new_n850), .B(KEYINPUT125), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n687), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n685), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n954), .A2(new_n579), .A3(new_n739), .A4(new_n843), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n783), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n795), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n949), .B1(new_n958), .B2(new_n189), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n949), .B1(new_n648), .B2(new_n189), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n765), .A2(new_n703), .A3(new_n851), .A4(new_n737), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n783), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n795), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n950), .A2(new_n749), .A3(new_n752), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n960), .B1(new_n965), .B2(new_n189), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n967));
  OR3_X1    g781(.A1(new_n959), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n959), .B2(new_n966), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(G72));
  NAND3_X1  g784(.A1(new_n963), .A2(new_n848), .A3(new_n964), .ZN(new_n971));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT63), .Z(new_n973));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n568), .B(KEYINPUT126), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n975), .A2(new_n539), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n876), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n569), .A2(new_n540), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n859), .A2(new_n973), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n975), .A2(new_n539), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n953), .A2(new_n957), .A3(new_n848), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n981), .B1(new_n982), .B2(new_n973), .ZN(new_n983));
  OAI21_X1  g797(.A(KEYINPUT127), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n983), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n985), .A2(new_n986), .A3(new_n979), .A4(new_n977), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n984), .A2(new_n987), .ZN(G57));
endmodule


