//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n449, new_n450, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n449));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  INV_X1    g026(.A(new_n450), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n452), .A2(G567), .ZN(G234));
  NAND2_X1  g028(.A1(new_n452), .A2(G2106), .ZN(G217));
  NAND4_X1  g029(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n455));
  XNOR2_X1  g030(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NAND4_X1  g032(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n457), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n457), .A2(G2106), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n473), .A2(new_n475), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(KEYINPUT68), .A2(G113), .A3(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g056(.A(G2105), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AND3_X1   g059(.A1(KEYINPUT68), .A2(G113), .A3(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(KEYINPUT68), .B1(G113), .B2(G2104), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n473), .A2(new_n475), .A3(G125), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n489), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n472), .B1(new_n484), .B2(new_n490), .ZN(G160));
  NAND2_X1  g066(.A1(new_n473), .A2(new_n475), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(new_n469), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G124), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n492), .A2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G136), .ZN(new_n496));
  OR2_X1    g071(.A1(G100), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n494), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G162));
  NAND4_X1  g075(.A1(new_n473), .A2(new_n475), .A3(G138), .A4(new_n469), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n468), .A2(new_n503), .A3(G138), .A4(new_n469), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n473), .A2(new_n475), .A3(G126), .A4(G2105), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  OR2_X1    g082(.A1(G102), .A2(G2105), .ZN(new_n508));
  INV_X1    g083(.A(G114), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G2105), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(new_n510), .A3(G2104), .ZN(new_n511));
  AND3_X1   g086(.A1(new_n506), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n507), .B1(new_n506), .B2(new_n511), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n505), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G164));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G50), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n525), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n523), .A2(new_n529), .ZN(G166));
  AND2_X1   g105(.A1(new_n520), .A2(new_n524), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  INV_X1    g107(.A(new_n527), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n532), .A2(new_n534), .A3(new_n535), .A4(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n517), .A2(new_n519), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G651), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n525), .A2(new_n546), .B1(new_n527), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n531), .A2(G81), .B1(new_n533), .B2(G43), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n541), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT71), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n553), .A2(KEYINPUT71), .A3(G651), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n550), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT72), .Z(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g141(.A(new_n566), .B(KEYINPUT73), .Z(G188));
  NAND3_X1  g142(.A1(new_n524), .A2(G53), .A3(G543), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT9), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n541), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n531), .A2(G91), .B1(new_n572), .B2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(new_n548), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n575), .A2(new_n576), .A3(new_n544), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT74), .B1(new_n545), .B2(new_n548), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G301));
  INV_X1    g154(.A(G166), .ZN(G303));
  OAI21_X1  g155(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n581));
  INV_X1    g156(.A(G49), .ZN(new_n582));
  INV_X1    g157(.A(G87), .ZN(new_n583));
  OAI221_X1 g158(.A(new_n581), .B1(new_n527), .B2(new_n582), .C1(new_n583), .C2(new_n525), .ZN(G288));
  AOI22_X1  g159(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n522), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  INV_X1    g162(.A(G48), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n525), .A2(new_n587), .B1(new_n527), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n522), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n525), .A2(new_n594), .B1(new_n527), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n531), .A2(new_n599), .A3(G92), .ZN(new_n600));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  OAI21_X1  g176(.A(KEYINPUT10), .B1(new_n525), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n541), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(G54), .A2(new_n533), .B1(new_n606), .B2(G651), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(KEYINPUT75), .B1(new_n609), .B2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  MUX2_X1   g186(.A(KEYINPUT75), .B(new_n610), .S(new_n611), .Z(G284));
  XNOR2_X1  g187(.A(G284), .B(KEYINPUT76), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G299), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n609), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n609), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n468), .A2(new_n466), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2100), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT77), .B(KEYINPUT13), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n493), .A2(G123), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT78), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n495), .A2(G135), .ZN(new_n632));
  OR2_X1    g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n633), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n493), .A2(KEYINPUT78), .A3(G123), .ZN(new_n635));
  NAND4_X1  g210(.A1(new_n631), .A2(new_n632), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n628), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT15), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n643), .A2(G2435), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(G2435), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT81), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT80), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n651), .B(new_n652), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n646), .A2(new_n648), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n649), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n649), .B2(new_n654), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n640), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n659), .A2(new_n655), .A3(new_n639), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n660), .A3(G14), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XOR2_X1   g238(.A(KEYINPUT82), .B(KEYINPUT17), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XOR2_X1   g241(.A(G2067), .B(G2678), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n665), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n666), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n663), .A2(new_n667), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n669), .B(new_n670), .C1(new_n666), .C2(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(KEYINPUT18), .B1(new_n670), .B2(new_n663), .ZN(new_n673));
  OR3_X1    g248(.A1(new_n670), .A2(KEYINPUT18), .A3(new_n663), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2096), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT83), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT20), .Z(new_n686));
  NOR2_X1   g261(.A1(new_n681), .A2(new_n682), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n688), .A2(new_n680), .A3(new_n683), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n686), .B(new_n689), .C1(new_n680), .C2(new_n688), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT84), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT85), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  INV_X1    g270(.A(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n694), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n692), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(G229));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n702), .A2(KEYINPUT23), .A3(G20), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT23), .ZN(new_n704));
  INV_X1    g279(.A(G20), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(G16), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n703), .B(new_n706), .C1(new_n615), .C2(new_n702), .ZN(new_n707));
  INV_X1    g282(.A(G1956), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G35), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G162), .B2(new_n710), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G2090), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT95), .Z(new_n716));
  NOR2_X1   g291(.A1(G29), .A2(G33), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(new_n469), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G139), .B2(new_n495), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n466), .A2(G103), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT25), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n717), .B1(new_n725), .B2(G29), .ZN(new_n726));
  NOR2_X1   g301(.A1(G5), .A2(G16), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G171), .B2(G16), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n726), .A2(G2072), .B1(G1961), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n713), .A2(G2090), .ZN(new_n730));
  NAND2_X1  g305(.A1(G168), .A2(G16), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G16), .B2(G21), .ZN(new_n732));
  INV_X1    g307(.A(G1966), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT94), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n468), .A2(G141), .A3(new_n469), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT26), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n468), .A2(G129), .A3(G2105), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n466), .A2(G105), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n737), .A2(new_n740), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G29), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G29), .B2(G32), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT27), .B(G1996), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n730), .B(new_n736), .C1(KEYINPUT93), .C2(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n716), .A2(new_n729), .A3(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n746), .A2(new_n747), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n726), .A2(G2072), .ZN(new_n753));
  INV_X1    g328(.A(G11), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n752), .B(new_n753), .C1(KEYINPUT31), .C2(new_n754), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n755), .B1(KEYINPUT31), .B2(new_n754), .C1(new_n733), .C2(new_n732), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n702), .A2(G19), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n559), .B2(new_n702), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(G1341), .Z(new_n759));
  NAND3_X1  g334(.A1(new_n468), .A2(G128), .A3(G2105), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n468), .A2(G140), .A3(new_n469), .ZN(new_n761));
  OR2_X1    g336(.A1(G104), .A2(G2105), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n762), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT89), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n710), .A2(G26), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT28), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G2067), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n759), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G2078), .ZN(new_n773));
  NOR2_X1   g348(.A1(G164), .A2(new_n710), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G27), .B2(new_n710), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n734), .A2(new_n735), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT90), .B(KEYINPUT24), .Z(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(G34), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(G34), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n778), .A2(new_n710), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT91), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G160), .B2(G29), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n780), .A2(new_n781), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI221_X1 g360(.A(new_n776), .B1(new_n773), .B2(new_n775), .C1(G2084), .C2(new_n785), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n750), .A2(new_n756), .A3(new_n772), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n702), .A2(G6), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n590), .B2(new_n702), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT32), .B(G1981), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n789), .B(new_n790), .Z(new_n791));
  NOR2_X1   g366(.A1(G16), .A2(G22), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G166), .B2(G16), .ZN(new_n793));
  INV_X1    g368(.A(G1971), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G16), .A2(G23), .ZN(new_n796));
  XNOR2_X1  g371(.A(G288), .B(KEYINPUT87), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT33), .B(G1976), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n791), .B(new_n795), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT34), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n493), .A2(G119), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n495), .A2(G131), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n469), .A2(G107), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n805), .B(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT86), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n710), .A2(G25), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n809), .A2(G29), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n810), .B2(new_n811), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT35), .B(G1991), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n813), .B(new_n814), .Z(new_n815));
  NOR2_X1   g390(.A1(G16), .A2(G24), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n597), .B2(G16), .ZN(new_n817));
  INV_X1    g392(.A(G1986), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n804), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n820), .A2(new_n823), .A3(new_n821), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT30), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n825), .A2(G28), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(G28), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n826), .A2(new_n827), .A3(new_n710), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n636), .B2(new_n710), .ZN(new_n829));
  INV_X1    g404(.A(new_n728), .ZN(new_n830));
  INV_X1    g405(.A(G1961), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n787), .A2(new_n822), .A3(new_n824), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n785), .A2(G2084), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT92), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n748), .A2(KEYINPUT93), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n702), .A2(G4), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n609), .B2(new_n702), .ZN(new_n838));
  INV_X1    g413(.A(G1348), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NOR4_X1   g416(.A1(new_n833), .A2(new_n835), .A3(new_n836), .A4(new_n841), .ZN(G311));
  INV_X1    g417(.A(new_n833), .ZN(new_n843));
  INV_X1    g418(.A(new_n835), .ZN(new_n844));
  INV_X1    g419(.A(new_n836), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n840), .ZN(G150));
  INV_X1    g421(.A(G67), .ZN(new_n847));
  INV_X1    g422(.A(G80), .ZN(new_n848));
  OAI22_X1  g423(.A1(new_n541), .A2(new_n847), .B1(new_n848), .B2(new_n516), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT96), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI221_X1 g426(.A(KEYINPUT96), .B1(new_n848), .B2(new_n516), .C1(new_n541), .C2(new_n847), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n851), .A2(G651), .A3(new_n852), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n531), .A2(G93), .B1(new_n533), .B2(G55), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n855), .B1(new_n853), .B2(new_n854), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G860), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  AOI21_X1  g436(.A(new_n558), .B1(new_n854), .B2(new_n853), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n558), .B1(new_n857), .B2(new_n858), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n609), .A2(G559), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n861), .B1(new_n869), .B2(G860), .ZN(G145));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n744), .A2(new_n764), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n506), .A2(new_n511), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(new_n502), .B2(new_n504), .ZN(new_n874));
  INV_X1    g449(.A(new_n764), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n743), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n874), .B1(new_n872), .B2(new_n876), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT101), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n881));
  INV_X1    g456(.A(new_n873), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n505), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n876), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n875), .A2(new_n743), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n881), .B1(new_n886), .B2(new_n877), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n724), .B1(new_n880), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT102), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT101), .B1(new_n878), .B2(new_n879), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n886), .A2(new_n881), .A3(new_n877), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n893), .A3(new_n724), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n493), .A2(G130), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n495), .A2(G142), .ZN(new_n897));
  OAI21_X1  g472(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n469), .A2(G118), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n896), .B(new_n897), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n809), .B(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n625), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n904), .ZN(new_n906));
  INV_X1    g481(.A(new_n625), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT100), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT100), .B1(new_n878), .B2(new_n879), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n725), .A3(new_n910), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n895), .A2(new_n905), .A3(new_n908), .A4(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n893), .B1(new_n892), .B2(new_n724), .ZN(new_n913));
  AOI211_X1 g488(.A(KEYINPUT102), .B(new_n725), .C1(new_n890), .C2(new_n891), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n908), .A2(new_n905), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g492(.A(KEYINPUT98), .B(KEYINPUT99), .Z(new_n918));
  XNOR2_X1  g493(.A(new_n636), .B(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(G160), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(G162), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n912), .A2(new_n917), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n912), .A2(new_n917), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT104), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n921), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n871), .B(new_n923), .C1(new_n925), .C2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g504(.A1(G303), .A2(G290), .ZN(new_n930));
  NAND2_X1  g505(.A1(G166), .A2(new_n597), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n930), .A2(G305), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G305), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n797), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n930), .A2(new_n931), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n590), .ZN(new_n936));
  XOR2_X1   g511(.A(G288), .B(KEYINPUT87), .Z(new_n937));
  NAND3_X1  g512(.A1(new_n930), .A2(G305), .A3(new_n931), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n941));
  XOR2_X1   g516(.A(new_n941), .B(KEYINPUT105), .Z(new_n942));
  NOR2_X1   g517(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT106), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n865), .B(new_n620), .ZN(new_n945));
  INV_X1    g520(.A(new_n603), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n946), .A2(new_n573), .A3(new_n569), .A4(new_n607), .ZN(new_n947));
  OAI21_X1  g522(.A(G299), .B1(new_n608), .B2(new_n603), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT41), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n947), .A2(KEYINPUT41), .A3(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n947), .A2(new_n948), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n952), .B2(new_n945), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n942), .A2(new_n944), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n942), .B2(new_n944), .ZN(new_n955));
  INV_X1    g530(.A(G868), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT107), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(new_n859), .B2(new_n956), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n957), .B2(new_n960), .ZN(G295));
  OAI21_X1  g536(.A(new_n958), .B1(new_n957), .B2(new_n960), .ZN(G331));
  INV_X1    g537(.A(KEYINPUT43), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n950), .A2(new_n949), .ZN(new_n964));
  AND2_X1   g539(.A1(G286), .A2(G171), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n965), .B1(G168), .B2(G301), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n865), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(G301), .A2(G168), .ZN(new_n968));
  INV_X1    g543(.A(new_n965), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n970), .A2(new_n864), .A3(new_n863), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n964), .A2(new_n967), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT108), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n967), .A2(new_n971), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n952), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n964), .A2(new_n967), .A3(new_n971), .A4(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n973), .A2(new_n940), .A3(new_n975), .A4(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n978), .A2(new_n871), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n972), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n940), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT109), .B1(new_n934), .B2(new_n939), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n963), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT110), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n940), .B(new_n981), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n973), .A2(new_n975), .A3(new_n977), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n979), .A2(new_n963), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT44), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n963), .B1(new_n979), .B2(new_n989), .ZN(new_n992));
  AND4_X1   g567(.A1(new_n963), .A2(new_n984), .A3(new_n871), .A4(new_n978), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI22_X1  g569(.A1(new_n986), .A2(new_n991), .B1(KEYINPUT44), .B2(new_n994), .ZN(G397));
  INV_X1    g570(.A(KEYINPUT122), .ZN(new_n996));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n883), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n998), .A2(G160), .A3(G40), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT45), .B1(new_n514), .B2(new_n997), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT113), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n874), .A2(new_n1002), .A3(G1384), .ZN(new_n1003));
  INV_X1    g578(.A(new_n472), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT69), .B1(new_n489), .B2(G2105), .ZN(new_n1005));
  AOI211_X1 g580(.A(new_n483), .B(new_n469), .C1(new_n487), .C2(new_n488), .ZN(new_n1006));
  OAI211_X1 g581(.A(G40), .B(new_n1004), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n514), .A2(new_n997), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n1002), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1001), .A2(new_n1012), .A3(new_n773), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1007), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n883), .A2(new_n997), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n1002), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1016), .B(new_n1018), .C1(new_n1002), .C2(new_n1010), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1014), .A2(G2078), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1384), .B1(new_n505), .B2(new_n882), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR4_X1   g601(.A1(new_n874), .A2(KEYINPUT114), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1007), .B1(KEYINPUT50), .B2(new_n1010), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1961), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1022), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1015), .A2(new_n1031), .A3(G301), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n482), .A2(G40), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT120), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n1004), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1018), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1034), .B1(new_n1033), .B2(new_n1004), .ZN(new_n1037));
  NOR4_X1   g612(.A1(new_n1036), .A2(new_n1037), .A3(new_n1003), .A4(new_n1021), .ZN(new_n1038));
  AOI211_X1 g613(.A(new_n1030), .B(new_n1038), .C1(new_n1014), .C2(new_n1013), .ZN(new_n1039));
  INV_X1    g614(.A(G171), .ZN(new_n1040));
  OAI211_X1 g615(.A(KEYINPUT54), .B(new_n1032), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1007), .A2(new_n1017), .ZN(new_n1042));
  INV_X1    g617(.A(G8), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1044), .B1(new_n937), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT52), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G305), .A2(G1981), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n590), .A2(new_n696), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1048), .A2(KEYINPUT49), .A3(new_n1049), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n1044), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT52), .B1(G288), .B2(new_n1045), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1044), .B(new_n1055), .C1(new_n937), .C2(new_n1045), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1047), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1001), .A2(new_n1012), .ZN(new_n1058));
  INV_X1    g633(.A(G2090), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1028), .A2(new_n1059), .A3(new_n1029), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1058), .A2(new_n794), .B1(KEYINPUT115), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1028), .A2(new_n1029), .A3(new_n1062), .A4(new_n1059), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1043), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(G303), .A2(G8), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1065), .B(KEYINPUT55), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1057), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1019), .A2(new_n733), .ZN(new_n1069));
  INV_X1    g644(.A(G2084), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1028), .A2(new_n1070), .A3(new_n1029), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(new_n1071), .A3(G168), .ZN(new_n1072));
  AOI21_X1  g647(.A(G168), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1072), .B(G8), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1072), .A2(G8), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1971), .B1(new_n1001), .B2(new_n1012), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1007), .B1(KEYINPUT50), .B2(new_n1017), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n514), .A2(new_n1025), .A3(new_n997), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(G2090), .ZN(new_n1082));
  OAI21_X1  g657(.A(G8), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1066), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1041), .A2(new_n1068), .A3(new_n1077), .A4(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1038), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1030), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1015), .A2(G301), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1086), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1015), .A2(new_n1031), .ZN(new_n1092));
  INV_X1    g667(.A(G301), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT121), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1091), .B1(new_n1094), .B2(new_n1089), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n996), .B1(new_n1085), .B2(new_n1095), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1041), .A2(new_n1077), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1089), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1039), .A2(KEYINPUT121), .A3(G301), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n1086), .A3(new_n1099), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n999), .A2(KEYINPUT113), .A3(new_n1000), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1009), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n794), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1060), .A2(KEYINPUT115), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1103), .A2(new_n1063), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(G8), .A3(new_n1067), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1057), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1106), .A2(new_n1107), .A3(new_n1084), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1097), .A2(new_n1100), .A3(KEYINPUT122), .A4(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1956), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(G299), .B(KEYINPUT57), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1008), .A2(new_n1011), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n839), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT117), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1042), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT117), .B1(new_n1007), .B2(new_n1017), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(new_n770), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1116), .A2(new_n1123), .A3(new_n609), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1111), .A2(KEYINPUT118), .A3(new_n1115), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1115), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(new_n1127), .B2(new_n1110), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(new_n1128), .A3(new_n1112), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1112), .B1(new_n1127), .B2(new_n1110), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1116), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT58), .B(G1341), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n999), .A2(G1996), .A3(new_n1000), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n559), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1137), .A2(KEYINPUT119), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1131), .A2(new_n1132), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1129), .A2(KEYINPUT61), .A3(new_n1116), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1137), .A2(KEYINPUT119), .ZN(new_n1141));
  OR3_X1    g716(.A1(new_n1136), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1118), .A2(new_n1143), .A3(new_n609), .A4(new_n1122), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1139), .A2(new_n1140), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1123), .A2(new_n609), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1123), .A2(new_n609), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1143), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1124), .B(new_n1129), .C1(new_n1145), .C2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1096), .A2(new_n1109), .A3(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT63), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI211_X1 g728(.A(new_n1043), .B(G286), .C1(new_n1069), .C2(new_n1071), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT63), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1106), .A2(new_n1107), .A3(new_n1084), .A4(new_n1154), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1153), .A2(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1107), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1054), .A2(new_n1045), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1049), .B1(new_n1159), .B2(G288), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1044), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT116), .B1(new_n1157), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1164), .B1(new_n1077), .B2(KEYINPUT62), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1165), .B(new_n1108), .C1(KEYINPUT62), .C2(new_n1077), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1105), .A2(G8), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1155), .B1(new_n1167), .B2(new_n1066), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1068), .A2(new_n1168), .A3(new_n1154), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1156), .A2(new_n1155), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT116), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1171), .A2(new_n1172), .A3(new_n1158), .A4(new_n1161), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1150), .A2(new_n1163), .A3(new_n1166), .A4(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1018), .A2(new_n1007), .ZN(new_n1175));
  INV_X1    g750(.A(G1996), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1177), .A2(new_n743), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n1178), .A2(KEYINPUT111), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1175), .B(KEYINPUT112), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n764), .B(new_n770), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1181), .B1(new_n744), .B2(new_n1176), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1178), .A2(KEYINPUT111), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1179), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n809), .B(new_n814), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1180), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n597), .B(new_n818), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1188), .B1(new_n1175), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1174), .A2(new_n1190), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1177), .B(KEYINPUT46), .Z(new_n1192));
  NAND2_X1  g767(.A1(new_n1181), .A2(new_n744), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1192), .B1(new_n1180), .B2(new_n1193), .ZN(new_n1194));
  XOR2_X1   g769(.A(KEYINPUT123), .B(KEYINPUT47), .Z(new_n1195));
  XNOR2_X1  g770(.A(new_n1194), .B(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1185), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n809), .A2(new_n814), .ZN(new_n1198));
  OAI22_X1  g773(.A1(new_n1197), .A2(new_n1198), .B1(G2067), .B2(new_n764), .ZN(new_n1199));
  AND2_X1   g774(.A1(new_n1199), .A2(new_n1180), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1175), .A2(new_n818), .A3(new_n597), .ZN(new_n1201));
  XOR2_X1   g776(.A(KEYINPUT125), .B(KEYINPUT48), .Z(new_n1202));
  XNOR2_X1  g777(.A(new_n1201), .B(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1188), .B(KEYINPUT124), .ZN(new_n1204));
  AOI211_X1 g779(.A(new_n1196), .B(new_n1200), .C1(new_n1203), .C2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1191), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n1208));
  OAI211_X1 g782(.A(G319), .B(new_n700), .C1(new_n992), .C2(new_n993), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n661), .A2(new_n677), .ZN(new_n1210));
  INV_X1    g784(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g785(.A1(new_n928), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g786(.A(new_n1208), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1213));
  AND2_X1   g787(.A1(new_n926), .A2(new_n921), .ZN(new_n1214));
  NAND3_X1  g788(.A1(new_n912), .A2(new_n917), .A3(new_n924), .ZN(new_n1215));
  AOI21_X1  g789(.A(G37), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g790(.A(new_n1210), .B1(new_n1216), .B2(new_n923), .ZN(new_n1217));
  AND2_X1   g791(.A1(new_n987), .A2(new_n988), .ZN(new_n1218));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n871), .ZN(new_n1219));
  OAI21_X1  g793(.A(KEYINPUT43), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g794(.A1(new_n979), .A2(new_n963), .A3(new_n984), .ZN(new_n1221));
  AOI21_X1  g795(.A(new_n463), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND4_X1  g796(.A1(new_n1217), .A2(new_n1222), .A3(KEYINPUT126), .A4(new_n700), .ZN(new_n1223));
  AND2_X1   g797(.A1(new_n1213), .A2(new_n1223), .ZN(G308));
  NAND2_X1  g798(.A1(new_n1213), .A2(new_n1223), .ZN(G225));
endmodule


