//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n458), .A2(KEYINPUT67), .B1(new_n448), .B2(new_n454), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(KEYINPUT67), .B2(new_n458), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  OAI21_X1  g036(.A(KEYINPUT68), .B1(new_n461), .B2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n461), .A2(G2104), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n462), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(new_n467), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n466), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n464), .A2(G2105), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NOR3_X1   g051(.A1(new_n470), .A2(new_n474), .A3(new_n476), .ZN(G160));
  INV_X1    g052(.A(new_n468), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n466), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n462), .A2(new_n465), .A3(G2105), .A4(new_n467), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n484));
  OR2_X1    g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n484), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n482), .B1(new_n487), .B2(G124), .ZN(new_n488));
  XOR2_X1   g063(.A(new_n488), .B(KEYINPUT70), .Z(G162));
  NAND2_X1  g064(.A1(new_n471), .A2(new_n467), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR4_X1   g066(.A1(new_n490), .A2(KEYINPUT4), .A3(new_n491), .A4(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n491), .A2(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n462), .A2(new_n465), .A3(new_n467), .A4(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n493), .B1(new_n495), .B2(KEYINPUT72), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n461), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n499), .A2(new_n500), .A3(new_n462), .A4(new_n494), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n492), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G2105), .ZN(new_n505));
  NOR3_X1   g080(.A1(new_n466), .A2(KEYINPUT71), .A3(G114), .ZN(new_n506));
  OAI221_X1 g081(.A(G2104), .B1(G102), .B2(G2105), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G126), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(new_n483), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n502), .A2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n515), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n520), .A2(new_n523), .ZN(G166));
  NAND2_X1  g099(.A1(new_n518), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT73), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n514), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n518), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n531));
  INV_X1    g106(.A(new_n517), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n534));
  AND3_X1   g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n530), .A2(new_n533), .A3(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  AND2_X1   g113(.A1(new_n529), .A2(G52), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n540), .A2(new_n522), .B1(new_n519), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  NAND2_X1  g118(.A1(new_n529), .A2(G43), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n532), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n519), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n547), .A2(G651), .B1(new_n548), .B2(G81), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G860), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n548), .A2(G91), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT76), .B(G65), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n532), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(G78), .B2(G543), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n558), .B1(new_n561), .B2(new_n522), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n514), .A2(G53), .ZN(new_n563));
  XOR2_X1   g138(.A(new_n563), .B(KEYINPUT9), .Z(new_n564));
  NOR2_X1   g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G299));
  OAI21_X1  g141(.A(KEYINPUT77), .B1(new_n539), .B2(new_n542), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NOR3_X1   g143(.A1(new_n539), .A2(KEYINPUT77), .A3(new_n542), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(G301));
  OAI221_X1 g145(.A(new_n515), .B1(new_n519), .B2(new_n516), .C1(new_n521), .C2(new_n522), .ZN(G303));
  OAI21_X1  g146(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n517), .A2(new_n518), .A3(G87), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n518), .A2(G49), .A3(G543), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  AND2_X1   g150(.A1(KEYINPUT5), .A2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(KEYINPUT5), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(G61), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(KEYINPUT78), .B1(G73), .B2(G543), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n517), .A2(new_n580), .A3(G61), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n522), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n519), .A2(new_n583), .B1(new_n525), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  AND2_X1   g162(.A1(new_n529), .A2(G47), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n589), .A2(new_n522), .B1(new_n519), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  INV_X1    g168(.A(G301), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n517), .A2(G66), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT80), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n522), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(new_n529), .B2(G54), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(KEYINPUT81), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n602));
  INV_X1    g177(.A(G54), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n526), .B2(new_n528), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n602), .B1(new_n604), .B2(new_n599), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OR3_X1    g182(.A1(new_n519), .A2(KEYINPUT79), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT79), .B1(new_n519), .B2(new_n607), .ZN(new_n609));
  AND3_X1   g184(.A1(new_n608), .A2(KEYINPUT10), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(KEYINPUT10), .B1(new_n608), .B2(new_n609), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n595), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT82), .ZN(G284));
  INV_X1    g191(.A(new_n615), .ZN(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n565), .B2(G868), .ZN(G297));
  OAI21_X1  g194(.A(new_n618), .B1(new_n565), .B2(G868), .ZN(G280));
  AND2_X1   g195(.A1(new_n606), .A2(new_n612), .ZN(new_n621));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G860), .ZN(G148));
  NOR2_X1   g198(.A1(new_n550), .A2(G868), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n613), .A2(G559), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT83), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n624), .B1(new_n626), .B2(G868), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n478), .A2(G135), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT85), .ZN(new_n631));
  INV_X1    g206(.A(G111), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n630), .A2(new_n631), .B1(new_n632), .B2(G2105), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n631), .B2(new_n630), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n485), .A2(new_n486), .ZN(new_n635));
  INV_X1    g210(.A(G123), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n629), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n637), .A2(G2096), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(G2096), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n640));
  NOR3_X1   g215(.A1(new_n461), .A2(new_n464), .A3(G2105), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n640), .B(new_n641), .Z(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT13), .B(G2100), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n638), .A2(new_n639), .A3(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT87), .B(G2438), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n646), .B(new_n647), .Z(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2430), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2451), .B(G2454), .Z(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(G14), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n656), .A2(new_n659), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(G401));
  XOR2_X1   g238(.A(KEYINPUT88), .B(KEYINPUT18), .Z(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT89), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  INV_X1    g247(.A(new_n664), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n672), .B1(new_n667), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2096), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT19), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n681), .A2(new_n682), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  MUX2_X1   g263(.A(new_n688), .B(new_n687), .S(new_n680), .Z(new_n689));
  NOR2_X1   g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1981), .ZN(new_n691));
  INV_X1    g266(.A(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT90), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n693), .A2(new_n695), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  OR3_X1    g274(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n696), .B2(new_n697), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(G229));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G21), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G168), .B2(new_n703), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT102), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G1966), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT103), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G35), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G162), .B2(new_n709), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT29), .B(G2090), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n709), .A2(G32), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT26), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n718), .A2(new_n719), .B1(G105), .B2(new_n475), .ZN(new_n720));
  INV_X1    g295(.A(G141), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n468), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n487), .A2(KEYINPUT100), .A3(G129), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT100), .ZN(new_n724));
  INV_X1    g299(.A(G129), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n635), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n722), .B1(new_n723), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n715), .B1(new_n727), .B2(new_n709), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT27), .B(G1996), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT101), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n728), .B(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G27), .A2(G29), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G164), .B2(G29), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(G2078), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n621), .A2(G16), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G4), .B2(G16), .ZN(new_n736));
  INV_X1    g311(.A(G1348), .ZN(new_n737));
  OAI22_X1  g312(.A1(new_n736), .A2(new_n737), .B1(G2078), .B2(new_n733), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n734), .B(new_n738), .C1(new_n737), .C2(new_n736), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n703), .A2(G20), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT23), .Z(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G299), .B2(G16), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1956), .ZN(new_n743));
  INV_X1    g318(.A(G19), .ZN(new_n744));
  OR3_X1    g319(.A1(new_n744), .A2(KEYINPUT97), .A3(G16), .ZN(new_n745));
  OAI21_X1  g320(.A(KEYINPUT97), .B1(new_n744), .B2(G16), .ZN(new_n746));
  INV_X1    g321(.A(new_n550), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n745), .B(new_n746), .C1(new_n747), .C2(new_n703), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G1341), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n709), .A2(G26), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT28), .Z(new_n751));
  OAI21_X1  g326(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n752));
  INV_X1    g327(.A(G116), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G2105), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n478), .B2(G140), .ZN(new_n755));
  INV_X1    g330(.A(G128), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n635), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n751), .B1(new_n757), .B2(G29), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2067), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT31), .B(G11), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT104), .B(G28), .Z(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n761), .B2(KEYINPUT30), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(KEYINPUT105), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT105), .ZN(new_n765));
  OAI22_X1  g340(.A1(new_n762), .A2(new_n765), .B1(KEYINPUT30), .B2(new_n761), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n760), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G34), .ZN(new_n768));
  AOI21_X1  g343(.A(G29), .B1(new_n768), .B2(KEYINPUT24), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(KEYINPUT24), .B2(new_n768), .ZN(new_n770));
  INV_X1    g345(.A(G160), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(new_n709), .ZN(new_n772));
  INV_X1    g347(.A(G2084), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n767), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n743), .A2(new_n749), .A3(new_n759), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n703), .A2(G5), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G171), .B2(new_n703), .ZN(new_n777));
  INV_X1    g352(.A(G1961), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  OAI221_X1 g354(.A(new_n779), .B1(new_n709), .B2(new_n637), .C1(new_n773), .C2(new_n772), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n706), .A2(G1966), .ZN(new_n781));
  NAND2_X1  g356(.A1(G115), .A2(G2104), .ZN(new_n782));
  INV_X1    g357(.A(G127), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n490), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n466), .B1(new_n784), .B2(KEYINPUT99), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(KEYINPUT99), .B2(new_n784), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT98), .B(KEYINPUT25), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G139), .B2(new_n478), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G33), .B(new_n791), .S(G29), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2072), .ZN(new_n793));
  NOR4_X1   g368(.A1(new_n775), .A2(new_n780), .A3(new_n781), .A4(new_n793), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n714), .A2(new_n731), .A3(new_n739), .A4(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT96), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT36), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n709), .A2(G25), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n487), .A2(KEYINPUT91), .A3(G119), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT91), .ZN(new_n802));
  INV_X1    g377(.A(G119), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n635), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n806));
  INV_X1    g381(.A(G107), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(G2105), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n478), .B2(G131), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT92), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n800), .B1(new_n812), .B2(new_n709), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT35), .B(G1991), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT93), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n813), .B(new_n815), .Z(new_n816));
  NAND2_X1  g391(.A1(new_n703), .A2(G22), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G166), .B2(new_n703), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT95), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G1971), .ZN(new_n820));
  NOR2_X1   g395(.A1(G6), .A2(G16), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n586), .B2(G16), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT32), .B(G1981), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n703), .A2(G23), .ZN(new_n825));
  INV_X1    g400(.A(G288), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n703), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT33), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G1976), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n820), .A2(new_n824), .A3(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n703), .A2(G24), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n592), .B2(new_n703), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n692), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n832), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n799), .B1(new_n816), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n816), .A2(new_n837), .A3(new_n799), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n796), .B1(new_n839), .B2(new_n840), .ZN(G150));
  INV_X1    g416(.A(G150), .ZN(G311));
  NOR2_X1   g417(.A1(new_n613), .A2(new_n622), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n529), .A2(G55), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(new_n522), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n846), .B1(KEYINPUT107), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(KEYINPUT107), .ZN(new_n850));
  INV_X1    g425(.A(G93), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n850), .B1(new_n851), .B2(new_n519), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(new_n747), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n550), .B1(new_n849), .B2(new_n852), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n845), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n859));
  AOI21_X1  g434(.A(G860), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n859), .B2(new_n858), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n853), .A2(new_n551), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT37), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(G145));
  XNOR2_X1  g439(.A(new_n637), .B(new_n771), .ZN(new_n865));
  XNOR2_X1  g440(.A(G162), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n868));
  INV_X1    g443(.A(G118), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n868), .A2(KEYINPUT109), .B1(new_n869), .B2(G2105), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(KEYINPUT109), .B2(new_n868), .ZN(new_n871));
  INV_X1    g446(.A(G142), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n872), .B2(new_n468), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(new_n487), .B2(G130), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n805), .A2(new_n875), .A3(new_n809), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n875), .B1(new_n805), .B2(new_n809), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n642), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n810), .A2(new_n874), .ZN(new_n880));
  INV_X1    g455(.A(new_n642), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(new_n881), .A3(new_n876), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n791), .A2(KEYINPUT108), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n757), .B(G164), .Z(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(new_n885), .B2(new_n727), .ZN(new_n886));
  INV_X1    g461(.A(new_n757), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n887), .A2(G164), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n757), .A2(new_n502), .A3(new_n509), .ZN(new_n889));
  OR3_X1    g464(.A1(new_n888), .A2(new_n727), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n791), .A2(KEYINPUT108), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n886), .A2(new_n892), .A3(new_n890), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n883), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n886), .A2(new_n892), .A3(new_n890), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n892), .B1(new_n886), .B2(new_n890), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n879), .A2(new_n882), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n867), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT110), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n899), .B1(new_n897), .B2(new_n898), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n894), .A2(new_n883), .A3(new_n895), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(KEYINPUT110), .A3(new_n867), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n904), .A2(new_n905), .A3(new_n866), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT40), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n914));
  AOI211_X1 g489(.A(new_n914), .B(new_n911), .C1(new_n903), .C2(new_n907), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n913), .A2(new_n915), .ZN(G395));
  XNOR2_X1  g491(.A(new_n626), .B(new_n857), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n613), .A2(KEYINPUT111), .A3(new_n565), .ZN(new_n918));
  NAND3_X1  g493(.A1(G299), .A2(new_n606), .A3(new_n612), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT111), .B1(new_n613), .B2(new_n565), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n626), .B(new_n856), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT41), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(new_n920), .B2(new_n922), .ZN(new_n928));
  XOR2_X1   g503(.A(KEYINPUT112), .B(KEYINPUT41), .Z(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n923), .A2(new_n919), .A3(new_n918), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n592), .B(G305), .ZN(new_n934));
  XNOR2_X1  g509(.A(G303), .B(new_n826), .ZN(new_n935));
  XOR2_X1   g510(.A(new_n934), .B(new_n935), .Z(new_n936));
  XOR2_X1   g511(.A(new_n936), .B(KEYINPUT42), .Z(new_n937));
  AND3_X1   g512(.A1(new_n925), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n937), .B1(new_n925), .B2(new_n933), .ZN(new_n939));
  OAI21_X1  g514(.A(G868), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(G868), .B2(new_n853), .ZN(G295));
  OAI21_X1  g516(.A(new_n940), .B1(G868), .B2(new_n853), .ZN(G331));
  OR3_X1    g517(.A1(new_n539), .A2(KEYINPUT77), .A3(new_n542), .ZN(new_n943));
  AOI21_X1  g518(.A(G286), .B1(new_n943), .B2(new_n567), .ZN(new_n944));
  NOR2_X1   g519(.A1(G168), .A2(G171), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n855), .B(new_n854), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(G168), .B1(new_n568), .B2(new_n569), .ZN(new_n947));
  INV_X1    g522(.A(new_n945), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n856), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n932), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n936), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n921), .A2(new_n923), .B1(new_n946), .B2(new_n949), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n946), .A2(new_n949), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n928), .B2(new_n931), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n936), .B1(new_n957), .B2(new_n953), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n955), .A2(new_n958), .A3(new_n910), .ZN(new_n959));
  XOR2_X1   g534(.A(KEYINPUT113), .B(KEYINPUT43), .Z(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n930), .B1(new_n920), .B2(new_n922), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n923), .A2(new_n927), .A3(new_n919), .A4(new_n918), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n950), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n936), .B1(new_n966), .B2(new_n953), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n967), .A2(new_n955), .A3(new_n910), .A4(new_n960), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n962), .A2(new_n963), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n955), .A3(new_n910), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n955), .A2(new_n958), .A3(new_n910), .A4(new_n960), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n963), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n969), .A2(new_n973), .ZN(G397));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n502), .B2(new_n509), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G40), .ZN(new_n979));
  NOR4_X1   g554(.A1(new_n470), .A2(new_n474), .A3(new_n979), .A4(new_n476), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G2067), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n757), .B(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT115), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n983), .B1(new_n986), .B2(new_n727), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT46), .ZN(new_n988));
  INV_X1    g563(.A(G1996), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n982), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n987), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT47), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n990), .A2(new_n988), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT125), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n992), .B1(new_n991), .B2(new_n994), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n986), .A2(new_n989), .ZN(new_n997));
  INV_X1    g572(.A(new_n990), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n987), .A2(new_n997), .B1(new_n727), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n810), .B(new_n815), .Z(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n982), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n982), .A2(new_n692), .A3(new_n592), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT127), .ZN(new_n1004));
  XOR2_X1   g579(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1005));
  XNOR2_X1  g580(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  OAI22_X1  g581(.A1(new_n995), .A2(new_n996), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n999), .A2(new_n812), .A3(new_n815), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n887), .A2(new_n984), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n983), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1013), .B(new_n975), .C1(new_n502), .C2(new_n509), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1014), .A2(new_n980), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n976), .A2(KEYINPUT116), .A3(KEYINPUT50), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT116), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n773), .B(new_n1015), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT45), .B(new_n975), .C1(new_n502), .C2(new_n509), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n978), .A2(new_n980), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1966), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1018), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1012), .B1(new_n1023), .B2(G286), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1018), .A2(G168), .A3(new_n1022), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(G8), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1012), .B1(new_n1025), .B2(G8), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT62), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1028), .ZN(new_n1030));
  AOI21_X1  g605(.A(G168), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1031));
  OAI211_X1 g606(.A(G8), .B(new_n1025), .C1(new_n1031), .C2(new_n1012), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT62), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1030), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n1035));
  INV_X1    g610(.A(G8), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(G166), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1041), .A2(new_n980), .A3(new_n1014), .ZN(new_n1042));
  INV_X1    g617(.A(G2090), .ZN(new_n1043));
  INV_X1    g618(.A(G1971), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1042), .A2(new_n1043), .B1(new_n1020), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1040), .B1(new_n1045), .B2(new_n1036), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1043), .B(new_n1015), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1020), .A2(new_n1044), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1038), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT117), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1037), .A2(new_n1053), .A3(new_n1038), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1049), .A2(G8), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT49), .ZN(new_n1058));
  INV_X1    g633(.A(G1981), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n579), .A2(new_n581), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G651), .ZN(new_n1061));
  INV_X1    g636(.A(new_n585), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n582), .A2(G1981), .A3(new_n585), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1058), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n980), .B(new_n975), .C1(new_n502), .C2(new_n509), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1061), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1067));
  OAI21_X1  g642(.A(G1981), .B1(new_n582), .B2(new_n585), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(KEYINPUT49), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1065), .A2(G8), .A3(new_n1066), .A4(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n572), .A2(new_n573), .A3(new_n574), .A4(G1976), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1071), .B(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(G8), .C1(new_n976), .C2(new_n981), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT52), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1070), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1976), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT52), .B1(G288), .B2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1066), .A2(G8), .A3(new_n1073), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT119), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1079), .A2(KEYINPUT119), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1076), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1046), .A2(new_n1057), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G2078), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n978), .A2(new_n1084), .A3(new_n980), .A4(new_n1019), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1019), .A2(new_n980), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1088), .A2(KEYINPUT53), .A3(new_n1084), .A4(new_n978), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1014), .A2(new_n980), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1041), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n976), .A2(KEYINPUT116), .A3(KEYINPUT50), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1090), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1087), .B(new_n1089), .C1(new_n1094), .C2(G1961), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n594), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1083), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1029), .A2(new_n1034), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n1100));
  NAND2_X1  g675(.A1(G168), .A2(G8), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1100), .B1(new_n1023), .B2(new_n1102), .ZN(new_n1103));
  AOI211_X1 g678(.A(KEYINPUT121), .B(new_n1101), .C1(new_n1018), .C2(new_n1022), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1099), .B1(new_n1105), .B2(new_n1083), .ZN(new_n1106));
  AOI211_X1 g681(.A(new_n1036), .B(new_n1055), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1080), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1079), .A2(KEYINPUT119), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1075), .B(new_n1070), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1049), .A2(G8), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1099), .B1(new_n1112), .B2(new_n1040), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1111), .B(new_n1113), .C1(new_n1104), .C2(new_n1103), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1106), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1066), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1070), .A2(new_n1077), .A3(new_n826), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1064), .B(KEYINPUT120), .ZN(new_n1118));
  AOI211_X1 g693(.A(new_n1036), .B(new_n1116), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1082), .B2(new_n1107), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1098), .A2(new_n1115), .A3(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n978), .A2(KEYINPUT123), .A3(new_n980), .A4(new_n1019), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT53), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1085), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n778), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n978), .A2(new_n980), .A3(new_n1019), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1127), .A2(KEYINPUT53), .A3(new_n1122), .A4(new_n1084), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .A4(G301), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1096), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(G171), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1126), .A2(G301), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(KEYINPUT54), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1083), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1132), .A2(new_n1133), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1139), .A2(KEYINPUT124), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1116), .A2(new_n984), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n1094), .B2(G1348), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n613), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1125), .A2(new_n737), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1146), .A2(KEYINPUT60), .A3(new_n621), .A4(new_n1141), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1144), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1015), .A2(new_n1041), .ZN(new_n1150));
  INV_X1    g725(.A(G1956), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(KEYINPUT56), .B(G2072), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1127), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n565), .B(KEYINPUT57), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1152), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1155), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1149), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1158), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1160), .A2(KEYINPUT61), .A3(new_n1156), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT58), .B(G1341), .ZN(new_n1162));
  OAI22_X1  g737(.A1(new_n1020), .A2(G1996), .B1(new_n1116), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n747), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT59), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1148), .A2(new_n1159), .A3(new_n1161), .A4(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT122), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1142), .A2(new_n1167), .A3(new_n621), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1160), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1167), .B1(new_n1142), .B2(new_n621), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1156), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1139), .A2(KEYINPUT124), .B1(new_n1166), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1121), .B1(new_n1140), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT114), .B1(G290), .B2(G1986), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n592), .A2(new_n692), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n999), .B(new_n1001), .C1(new_n983), .C2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1011), .B1(new_n1173), .B2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g753(.A(G319), .B1(new_n661), .B2(new_n662), .ZN(new_n1180));
  NOR2_X1   g754(.A1(new_n1180), .A2(G227), .ZN(new_n1181));
  AND3_X1   g755(.A1(new_n700), .A2(new_n701), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g756(.A(new_n907), .ZN(new_n1183));
  AOI21_X1  g757(.A(KEYINPUT110), .B1(new_n906), .B2(new_n867), .ZN(new_n1184));
  OAI21_X1  g758(.A(new_n912), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g759(.A1(new_n962), .A2(new_n968), .ZN(new_n1186));
  NAND3_X1  g760(.A1(new_n1182), .A2(new_n1185), .A3(new_n1186), .ZN(G225));
  INV_X1    g761(.A(G225), .ZN(G308));
endmodule


