//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n546, new_n548, new_n549, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n588,
    new_n589, new_n592, new_n594, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1132;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n452));
  AND2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  XNOR2_X1  g028(.A(G325), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT67), .Z(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G137), .ZN(new_n460));
  NAND2_X1  g035(.A1(G101), .A2(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n467), .B1(new_n464), .B2(new_n466), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n462), .B1(new_n472), .B2(G2105), .ZN(G160));
  NAND2_X1  g048(.A1(new_n464), .A2(new_n466), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n474), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(new_n475), .B2(G112), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n477), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OAI211_X1 g058(.A(G138), .B(new_n475), .C1(new_n468), .C2(new_n469), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g061(.A1(KEYINPUT4), .A2(G138), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n464), .A2(new_n466), .A3(new_n487), .A4(new_n475), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT69), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n459), .A2(new_n496), .A3(G126), .A4(G2105), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n486), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(G62), .A3(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n506), .A2(new_n513), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n509), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  INV_X1    g094(.A(new_n515), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n506), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G51), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n521), .A2(new_n524), .A3(new_n525), .A4(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  AOI22_X1  g104(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n503), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT71), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT72), .B(G52), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n523), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n520), .A2(G90), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  INV_X1    g113(.A(G43), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n538), .A2(new_n515), .B1(new_n522), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT73), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n503), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  AND3_X1   g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G36), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(G188));
  XNOR2_X1  g125(.A(new_n513), .B(KEYINPUT74), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n503), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n520), .A2(G91), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n523), .A2(G53), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(G299));
  NAND2_X1  g132(.A1(new_n520), .A2(G87), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n523), .A2(G49), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(G288));
  NAND2_X1  g136(.A1(G73), .A2(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n510), .A2(new_n512), .ZN(new_n563));
  INV_X1    g138(.A(G61), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n506), .A2(G48), .A3(G543), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n506), .A2(new_n513), .A3(G86), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G305));
  NAND2_X1  g144(.A1(new_n520), .A2(G85), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n523), .A2(G47), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n570), .B(new_n571), .C1(new_n503), .C2(new_n572), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(KEYINPUT75), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(KEYINPUT75), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G290));
  NAND2_X1  g151(.A1(G301), .A2(G868), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n551), .A2(G66), .ZN(new_n578));
  NAND2_X1  g153(.A1(G79), .A2(G543), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n503), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(G54), .B2(new_n523), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n520), .A2(G92), .ZN(new_n582));
  XOR2_X1   g157(.A(new_n582), .B(KEYINPUT10), .Z(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n577), .B1(new_n585), .B2(G868), .ZN(G284));
  OAI21_X1  g161(.A(new_n577), .B1(new_n585), .B2(G868), .ZN(G321));
  NAND2_X1  g162(.A1(G286), .A2(G868), .ZN(new_n588));
  XNOR2_X1  g163(.A(G299), .B(KEYINPUT76), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(G868), .ZN(G297));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(G868), .ZN(G280));
  INV_X1    g166(.A(G559), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n585), .B1(new_n592), .B2(G860), .ZN(G148));
  OAI21_X1  g168(.A(G868), .B1(new_n584), .B2(G559), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(G868), .B2(new_n544), .ZN(G323));
  XNOR2_X1  g170(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g171(.A1(new_n474), .A2(KEYINPUT68), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n599), .A2(G2104), .A3(new_n475), .ZN(new_n600));
  XOR2_X1   g175(.A(new_n600), .B(KEYINPUT12), .Z(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT13), .ZN(new_n602));
  NOR2_X1   g177(.A1(KEYINPUT77), .A2(G2100), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n476), .A2(G123), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n478), .A2(G135), .ZN(new_n606));
  OR2_X1    g181(.A1(G99), .A2(G2105), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n607), .B(G2104), .C1(G111), .C2(new_n475), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G2096), .B1(KEYINPUT77), .B2(G2100), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n604), .B(new_n610), .C1(G2096), .C2(new_n609), .ZN(G156));
  XNOR2_X1  g186(.A(KEYINPUT15), .B(G2430), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2435), .ZN(new_n613));
  XOR2_X1   g188(.A(G2427), .B(G2438), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(KEYINPUT14), .ZN(new_n616));
  XNOR2_X1  g191(.A(G2443), .B(G2446), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2451), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2454), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n618), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(G1341), .B(G1348), .Z(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT80), .Z(new_n626));
  NOR2_X1   g201(.A1(new_n622), .A2(new_n624), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT79), .ZN(new_n628));
  AND3_X1   g203(.A1(new_n626), .A2(G14), .A3(new_n628), .ZN(G401));
  XOR2_X1   g204(.A(G2067), .B(G2678), .Z(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2084), .B(G2090), .Z(new_n632));
  AND2_X1   g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2072), .B(G2078), .Z(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT81), .B(KEYINPUT18), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT82), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(KEYINPUT17), .B1(new_n631), .B2(new_n632), .ZN(new_n640));
  AND2_X1   g215(.A1(new_n640), .A2(new_n634), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(new_n634), .ZN(new_n642));
  NOR3_X1   g217(.A1(new_n641), .A2(new_n642), .A3(new_n633), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2096), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2100), .ZN(G227));
  XNOR2_X1  g221(.A(G1956), .B(G2474), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT83), .ZN(new_n648));
  XOR2_X1   g223(.A(G1961), .B(G1966), .Z(new_n649));
  AND2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G1971), .B(G1976), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT19), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT20), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n648), .A2(new_n649), .ZN(new_n655));
  AOI22_X1  g230(.A1(new_n653), .A2(new_n654), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  OR3_X1    g231(.A1(new_n650), .A2(new_n655), .A3(new_n652), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n656), .B(new_n657), .C1(new_n654), .C2(new_n653), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT21), .B(G1986), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G1991), .B(G1996), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT84), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n660), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT22), .B(G1981), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n663), .B(new_n664), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G229));
  OR2_X1    g241(.A1(G16), .A2(G22), .ZN(new_n667));
  INV_X1    g242(.A(G16), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n667), .B1(G303), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G1971), .ZN(new_n670));
  MUX2_X1   g245(.A(G6), .B(G305), .S(G16), .Z(new_n671));
  XOR2_X1   g246(.A(KEYINPUT32), .B(G1981), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(G16), .A2(G23), .ZN(new_n675));
  INV_X1    g250(.A(G288), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n675), .B1(new_n676), .B2(G16), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT33), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  OAI22_X1  g254(.A1(new_n674), .A2(new_n679), .B1(KEYINPUT88), .B2(KEYINPUT34), .ZN(new_n680));
  NAND2_X1  g255(.A1(KEYINPUT88), .A2(KEYINPUT34), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n680), .B(new_n681), .Z(new_n682));
  NOR2_X1   g257(.A1(G16), .A2(G24), .ZN(new_n683));
  INV_X1    g258(.A(G290), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(G16), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT87), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(G2104), .B1(new_n475), .B2(G107), .ZN(new_n688));
  INV_X1    g263(.A(G95), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(new_n475), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT85), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n476), .A2(G119), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n478), .A2(G131), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G25), .B(new_n694), .S(G29), .Z(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT35), .B(G1991), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT86), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n682), .A2(new_n687), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n699), .B(new_n700), .Z(new_n701));
  AND2_X1   g276(.A1(new_n668), .A2(G21), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G286), .B2(G16), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(G1966), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT31), .B(G11), .Z(new_n705));
  INV_X1    g280(.A(G28), .ZN(new_n706));
  OR3_X1    g281(.A1(new_n706), .A2(KEYINPUT95), .A3(KEYINPUT30), .ZN(new_n707));
  OAI21_X1  g282(.A(KEYINPUT95), .B1(new_n706), .B2(KEYINPUT30), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI211_X1 g284(.A(G29), .B(new_n709), .C1(KEYINPUT30), .C2(new_n706), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n704), .A2(new_n705), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  INV_X1    g287(.A(G1961), .ZN(new_n713));
  NAND2_X1  g288(.A1(G171), .A2(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G5), .B2(G16), .ZN(new_n715));
  OAI221_X1 g290(.A(new_n711), .B1(new_n712), .B2(new_n609), .C1(new_n713), .C2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT96), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n712), .A2(G26), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n476), .A2(G128), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT91), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n478), .A2(G140), .ZN(new_n724));
  NOR2_X1   g299(.A1(G104), .A2(G2105), .ZN(new_n725));
  OAI21_X1  g300(.A(G2104), .B1(new_n475), .B2(G116), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n720), .B1(new_n728), .B2(new_n712), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G2067), .ZN(new_n730));
  INV_X1    g305(.A(G34), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(KEYINPUT24), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(KEYINPUT24), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n712), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G160), .B2(new_n712), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G2084), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n712), .A2(G35), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n712), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT97), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT29), .ZN(new_n740));
  AOI211_X1 g315(.A(new_n730), .B(new_n736), .C1(new_n740), .C2(G2090), .ZN(new_n741));
  NOR2_X1   g316(.A1(G16), .A2(G19), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n544), .B2(G16), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT90), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1341), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n668), .A2(KEYINPUT23), .A3(G20), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT23), .ZN(new_n747));
  INV_X1    g322(.A(G20), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(G16), .ZN(new_n749));
  INV_X1    g324(.A(G299), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n746), .B(new_n749), .C1(new_n750), .C2(new_n668), .ZN(new_n751));
  INV_X1    g326(.A(G1956), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n717), .A2(new_n741), .A3(new_n745), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n668), .A2(G4), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n585), .B2(new_n668), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1348), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n715), .A2(new_n713), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n740), .B2(G2090), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n754), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(G164), .A2(G29), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G27), .B2(G29), .ZN(new_n762));
  INV_X1    g337(.A(G2078), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OR2_X1    g339(.A1(G29), .A2(G33), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n478), .A2(G139), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT25), .Z(new_n768));
  AOI22_X1  g343(.A1(new_n599), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT93), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n766), .B(new_n768), .C1(new_n770), .C2(new_n475), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n765), .B1(new_n771), .B2(new_n712), .ZN(new_n772));
  INV_X1    g347(.A(G2072), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n772), .A2(new_n773), .B1(new_n763), .B2(new_n762), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n701), .A2(new_n760), .A3(new_n764), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n772), .A2(new_n773), .ZN(new_n776));
  AOI22_X1  g351(.A1(G129), .A2(new_n476), .B1(new_n478), .B2(G141), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n475), .A2(G105), .A3(G2104), .ZN(new_n778));
  NAND3_X1  g353(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT26), .Z(new_n780));
  NAND3_X1  g355(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT94), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(new_n712), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n712), .B2(G32), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT27), .B(G1996), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n785), .B(new_n786), .Z(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n775), .A2(new_n776), .A3(new_n788), .ZN(G311));
  AND3_X1   g364(.A1(new_n701), .A2(new_n774), .A3(new_n760), .ZN(new_n790));
  INV_X1    g365(.A(new_n776), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n790), .A2(new_n791), .A3(new_n787), .A4(new_n764), .ZN(G150));
  NAND2_X1  g367(.A1(new_n520), .A2(G93), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n523), .A2(G55), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n793), .B(new_n794), .C1(new_n503), .C2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT99), .B(G860), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT37), .Z(new_n799));
  NOR2_X1   g374(.A1(new_n584), .A2(new_n592), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n544), .B(new_n796), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n802), .B(new_n803), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(KEYINPUT39), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT100), .ZN(new_n806));
  INV_X1    g381(.A(new_n797), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n804), .B2(KEYINPUT39), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n799), .B1(new_n806), .B2(new_n808), .ZN(G145));
  OR2_X1    g384(.A1(new_n783), .A2(new_n694), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n783), .A2(new_n694), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n478), .A2(G142), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT101), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n476), .A2(G130), .ZN(new_n816));
  OR2_X1    g391(.A1(G106), .A2(G2105), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n817), .B(G2104), .C1(G118), .C2(new_n475), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n478), .A2(KEYINPUT101), .A3(G142), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n815), .A2(new_n816), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n812), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n820), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n810), .A2(new_n822), .A3(new_n811), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT102), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n499), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n827), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n821), .A2(new_n823), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n771), .B(new_n728), .ZN(new_n832));
  INV_X1    g407(.A(new_n601), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n828), .A2(new_n834), .A3(new_n835), .A4(new_n830), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT105), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n609), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n837), .A2(new_n838), .A3(new_n839), .A4(new_n609), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(G160), .B(G162), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G37), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n842), .A2(new_n845), .A3(new_n843), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g426(.A1(new_n796), .A2(G868), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n684), .A2(new_n676), .ZN(new_n853));
  NAND2_X1  g428(.A1(G290), .A2(G288), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT106), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n853), .A2(KEYINPUT106), .A3(new_n854), .ZN(new_n858));
  XNOR2_X1  g433(.A(G303), .B(G305), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n859), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n855), .A2(new_n856), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(KEYINPUT42), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(KEYINPUT42), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n585), .A2(new_n750), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n584), .A2(G299), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT41), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n868), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT41), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n584), .A2(G559), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n803), .B(new_n875), .ZN(new_n876));
  MUX2_X1   g451(.A(new_n874), .B(new_n869), .S(new_n876), .Z(new_n877));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n865), .B(new_n866), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n879), .B(new_n880), .Z(new_n881));
  AOI21_X1  g456(.A(new_n852), .B1(new_n881), .B2(G868), .ZN(G295));
  AOI21_X1  g457(.A(new_n852), .B1(new_n881), .B2(G868), .ZN(G331));
  NAND3_X1  g458(.A1(new_n871), .A2(KEYINPUT109), .A3(new_n873), .ZN(new_n884));
  XNOR2_X1  g459(.A(G301), .B(G168), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n803), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n803), .A2(new_n885), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n884), .B(new_n888), .C1(KEYINPUT109), .C2(new_n873), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n872), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n863), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n874), .A2(new_n888), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n894), .A3(new_n864), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n848), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT43), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n871), .A2(new_n873), .B1(new_n886), .B2(new_n887), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n863), .B1(new_n898), .B2(new_n890), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(new_n899), .A3(new_n848), .ZN(new_n900));
  OR3_X1    g475(.A1(new_n900), .A2(KEYINPUT110), .A3(KEYINPUT43), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT110), .B1(new_n900), .B2(KEYINPUT43), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n897), .A2(new_n901), .A3(KEYINPUT44), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(KEYINPUT43), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT108), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n893), .A2(new_n906), .A3(new_n848), .A4(new_n895), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n900), .A2(new_n908), .A3(KEYINPUT43), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n903), .B1(new_n911), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g487(.A(KEYINPUT127), .ZN(new_n913));
  OR2_X1    g488(.A1(G290), .A2(G1986), .ZN(new_n914));
  NAND2_X1  g489(.A1(G290), .A2(G1986), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(G1384), .B1(new_n486), .B2(new_n498), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT111), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n917), .B(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n920));
  INV_X1    g495(.A(G40), .ZN(new_n921));
  AOI211_X1 g496(.A(new_n921), .B(new_n462), .C1(new_n472), .C2(G2105), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n916), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n728), .B(G2067), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT113), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n783), .ZN(new_n927));
  INV_X1    g502(.A(G1996), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n923), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n923), .A2(G1996), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n932), .A2(new_n783), .ZN(new_n933));
  OR2_X1    g508(.A1(new_n933), .A2(KEYINPUT112), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n694), .A2(new_n696), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n694), .A2(new_n696), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n930), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(KEYINPUT112), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n931), .A2(new_n934), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(G303), .A2(G8), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n940), .B(KEYINPUT55), .Z(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n917), .B(new_n920), .ZN(new_n943));
  AOI21_X1  g518(.A(G1971), .B1(new_n943), .B2(new_n922), .ZN(new_n944));
  AOI211_X1 g519(.A(KEYINPUT50), .B(G1384), .C1(new_n486), .C2(new_n498), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT50), .ZN(new_n946));
  OAI211_X1 g521(.A(G40), .B(G160), .C1(new_n917), .C2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT118), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT118), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n922), .B(new_n949), .C1(new_n946), .C2(new_n917), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n945), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G2090), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n944), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G8), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n942), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n462), .ZN(new_n956));
  INV_X1    g531(.A(new_n471), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n957), .B1(new_n599), .B2(G125), .ZN(new_n958));
  OAI211_X1 g533(.A(G40), .B(new_n956), .C1(new_n958), .C2(new_n475), .ZN(new_n959));
  INV_X1    g534(.A(G1384), .ZN(new_n960));
  AOI21_X1  g535(.A(G2105), .B1(new_n597), .B2(new_n598), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT4), .B1(new_n961), .B2(G138), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n495), .A2(new_n497), .ZN(new_n963));
  INV_X1    g538(.A(new_n493), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n960), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n959), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n967));
  INV_X1    g542(.A(new_n945), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n952), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n920), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n917), .A2(KEYINPUT45), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n970), .A2(new_n922), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n969), .B1(new_n972), .B2(G1971), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT114), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(KEYINPUT114), .B(new_n969), .C1(new_n972), .C2(G1971), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n975), .A2(G8), .A3(new_n941), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(G305), .A2(G1981), .ZN(new_n978));
  INV_X1    g553(.A(G1981), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n566), .A2(new_n979), .A3(new_n567), .A4(new_n568), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT49), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT49), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n978), .A2(new_n983), .A3(new_n980), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n986));
  AOI211_X1 g561(.A(new_n986), .B(new_n954), .C1(new_n922), .C2(new_n917), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n917), .A2(G40), .A3(G160), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT115), .B1(new_n988), .B2(G8), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n985), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1976), .ZN(new_n991));
  NOR2_X1   g566(.A1(G288), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(G8), .B1(new_n966), .B2(new_n959), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n986), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n988), .A2(KEYINPUT115), .A3(G8), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n990), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT116), .B(G1976), .ZN(new_n999));
  NAND2_X1  g574(.A1(G288), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n997), .ZN(new_n1001));
  AOI211_X1 g576(.A(new_n992), .B(new_n1001), .C1(new_n994), .C2(new_n995), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n955), .A2(new_n977), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1961), .B1(new_n967), .B2(new_n968), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n959), .A2(G2078), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n943), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1011));
  XNOR2_X1  g586(.A(G301), .B(KEYINPUT54), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1012), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n919), .A2(new_n920), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1015), .A2(KEYINPUT53), .A3(new_n971), .A4(new_n1008), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n1010), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G2084), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n967), .A2(new_n1018), .A3(new_n968), .ZN(new_n1019));
  OAI211_X1 g594(.A(G168), .B(new_n1019), .C1(new_n972), .C2(G1966), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(G8), .ZN(new_n1021));
  AND2_X1   g596(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1022));
  NOR2_X1   g597(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1020), .A2(G8), .A3(new_n1023), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1019), .B1(new_n972), .B2(G1966), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(G8), .A3(G286), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1013), .B(new_n1017), .C1(new_n1025), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1348), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n947), .B2(new_n945), .ZN(new_n1032));
  INV_X1    g607(.A(new_n988), .ZN(new_n1033));
  INV_X1    g608(.A(G2067), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1032), .A2(KEYINPUT60), .A3(new_n1035), .ZN(new_n1036));
  OR2_X1    g611(.A1(new_n1036), .A2(KEYINPUT121), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1036), .A2(KEYINPUT121), .A3(new_n584), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n584), .B1(new_n1036), .B2(KEYINPUT121), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT60), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT61), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT56), .B(G2072), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n970), .A2(new_n922), .A3(new_n1046), .A4(new_n971), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1047), .A2(KEYINPUT119), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(KEYINPUT119), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1048), .A2(new_n1049), .B1(new_n951), .B2(G1956), .ZN(new_n1050));
  XNOR2_X1  g625(.A(G299), .B(KEYINPUT57), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1045), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n951), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n752), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n943), .A2(new_n1055), .A3(new_n922), .A4(new_n1046), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1047), .A2(KEYINPUT119), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n1059));
  XNOR2_X1  g634(.A(G299), .B(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1054), .A2(new_n1058), .A3(KEYINPUT61), .A4(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1052), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n970), .A2(new_n928), .A3(new_n922), .A4(new_n971), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT58), .B(G1341), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1033), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n544), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT59), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(new_n1068), .A3(new_n544), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1067), .A2(new_n1069), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1044), .A2(new_n1062), .A3(new_n1070), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1053), .A2(new_n752), .B1(new_n1057), .B2(new_n1056), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n584), .B1(new_n1072), .B2(new_n1060), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1051), .B(KEYINPUT120), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1073), .A2(new_n1041), .B1(new_n1074), .B2(new_n1050), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1030), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT62), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(new_n1028), .A4(new_n1026), .ZN(new_n1080));
  AND4_X1   g655(.A1(G171), .A2(new_n1077), .A3(new_n1011), .A4(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1005), .B1(new_n1076), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT117), .B1(new_n998), .B2(new_n1002), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n987), .A2(new_n989), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT52), .B1(new_n1084), .B2(new_n992), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n996), .A2(new_n997), .A3(new_n1000), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .A4(new_n990), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1083), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1089), .A2(new_n977), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n990), .A2(new_n991), .A3(new_n676), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1084), .B1(new_n1091), .B2(new_n980), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1083), .A2(new_n1088), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1027), .A2(G8), .A3(G168), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT63), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n975), .A2(G8), .A3(new_n976), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n1097), .B2(new_n942), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1093), .A2(new_n977), .A3(new_n1095), .A4(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1096), .B1(new_n1004), .B2(new_n1094), .ZN(new_n1100));
  AOI211_X1 g675(.A(new_n1090), .B(new_n1092), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n924), .B(new_n939), .C1(new_n1082), .C2(new_n1101), .ZN(new_n1102));
  XOR2_X1   g677(.A(new_n936), .B(KEYINPUT123), .Z(new_n1103));
  NAND4_X1  g678(.A1(new_n931), .A2(new_n934), .A3(new_n938), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n728), .A2(new_n1034), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT124), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(new_n1108), .A3(new_n1105), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1107), .A2(new_n930), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT125), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n927), .A2(new_n930), .B1(new_n1111), .B2(KEYINPUT46), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(KEYINPUT46), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n932), .B(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT47), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n939), .A2(KEYINPUT126), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n914), .A2(new_n923), .ZN(new_n1118));
  XOR2_X1   g693(.A(new_n1118), .B(KEYINPUT48), .Z(new_n1119));
  NAND2_X1  g694(.A1(new_n939), .A2(KEYINPUT126), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1110), .A2(new_n1116), .A3(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n913), .B1(new_n1102), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1082), .A2(new_n1101), .ZN(new_n1124));
  INV_X1    g699(.A(new_n924), .ZN(new_n1125));
  INV_X1    g700(.A(new_n939), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1122), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1127), .A2(new_n1128), .A3(KEYINPUT127), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1123), .A2(new_n1129), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g705(.A1(G401), .A2(new_n457), .A3(G227), .ZN(new_n1132));
  NAND4_X1  g706(.A1(new_n910), .A2(new_n850), .A3(new_n665), .A4(new_n1132), .ZN(G225));
  INV_X1    g707(.A(G225), .ZN(G308));
endmodule


