//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1240, new_n1241, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(G1), .ZN(new_n213));
  NOR3_X1   g0013(.A1(new_n213), .A2(new_n209), .A3(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n211), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G97), .A2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n221), .B(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n220), .B(new_n225), .C1(G58), .C2(G232), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(G1), .B2(G20), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT1), .Z(new_n228));
  AOI211_X1 g0028(.A(new_n216), .B(new_n228), .C1(new_n212), .C2(new_n215), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n219), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G58), .ZN(new_n239));
  INV_X1    g0039(.A(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G97), .B(G107), .ZN(new_n242));
  INV_X1    g0042(.A(G87), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n218), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n241), .B(new_n245), .Z(G351));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(G222), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(G223), .ZN(new_n251));
  OAI221_X1 g0051(.A(new_n249), .B1(new_n240), .B2(new_n247), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n208), .B1(G33), .B2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT65), .B(G41), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n213), .B(G274), .C1(new_n255), .C2(G45), .ZN(new_n256));
  INV_X1    g0056(.A(new_n253), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n213), .B1(G41), .B2(G45), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G226), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n254), .A2(new_n256), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n203), .A2(G20), .ZN(new_n264));
  INV_X1    g0064(.A(G150), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT8), .B(G58), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n264), .B1(new_n265), .B2(new_n267), .C1(new_n268), .C2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n208), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n213), .A2(G13), .A3(G20), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n272), .A2(new_n274), .B1(new_n202), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n274), .B1(new_n213), .B2(G20), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G50), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n263), .A2(G190), .B1(new_n281), .B2(KEYINPUT9), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT70), .ZN(new_n283));
  INV_X1    g0083(.A(G200), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n283), .B1(new_n263), .B2(new_n284), .ZN(new_n285));
  OR2_X1    g0085(.A1(new_n281), .A2(KEYINPUT9), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n262), .A2(KEYINPUT70), .A3(G200), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n282), .A2(new_n285), .A3(new_n286), .A4(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n288), .B(KEYINPUT10), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n280), .B1(new_n263), .B2(G169), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT66), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(G179), .B2(new_n262), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT13), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n247), .A2(G226), .A3(new_n248), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n247), .A2(G232), .A3(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(G97), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n296), .B(new_n297), .C1(new_n269), .C2(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n299), .A2(new_n253), .B1(new_n260), .B2(G238), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n295), .B1(new_n300), .B2(new_n256), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(new_n295), .A3(new_n256), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT14), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n302), .A2(G179), .A3(new_n303), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT14), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(new_n308), .A3(G169), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT12), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n275), .B2(G68), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n276), .A2(KEYINPUT12), .A3(new_n223), .ZN(new_n313));
  INV_X1    g0113(.A(new_n278), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n312), .B(new_n313), .C1(new_n314), .C2(new_n223), .ZN(new_n315));
  XOR2_X1   g0115(.A(new_n315), .B(KEYINPUT71), .Z(new_n316));
  AOI22_X1  g0116(.A1(new_n270), .A2(G77), .B1(new_n266), .B2(G50), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n209), .B2(G68), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n274), .ZN(new_n319));
  XOR2_X1   g0119(.A(new_n319), .B(KEYINPUT11), .Z(new_n320));
  NOR2_X1   g0120(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n321), .B(KEYINPUT72), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n310), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n304), .A2(G200), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n302), .A2(G190), .A3(new_n303), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(new_n321), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n294), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n268), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(new_n276), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n314), .B2(new_n328), .ZN(new_n330));
  INV_X1    g0130(.A(new_n274), .ZN(new_n331));
  INV_X1    g0131(.A(G58), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(new_n223), .ZN(new_n333));
  OAI21_X1  g0133(.A(G20), .B1(new_n333), .B2(new_n201), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n266), .A2(G159), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT3), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G33), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n339), .A3(KEYINPUT73), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT73), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(new_n269), .A3(KEYINPUT3), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n209), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n223), .B1(new_n343), .B2(KEYINPUT7), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT7), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n340), .A2(new_n345), .A3(new_n209), .A4(new_n342), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n336), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n331), .B1(new_n347), .B2(KEYINPUT16), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(KEYINPUT74), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n345), .A2(KEYINPUT74), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n349), .B(new_n350), .C1(new_n247), .C2(G20), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n337), .A2(new_n339), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n352), .A2(KEYINPUT74), .A3(new_n345), .A4(new_n209), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n353), .A3(G68), .ZN(new_n354));
  INV_X1    g0154(.A(new_n336), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT16), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n330), .B1(new_n348), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT75), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n248), .A2(G226), .ZN(new_n361));
  NOR2_X1   g0161(.A1(G223), .A2(G1698), .ZN(new_n362));
  AOI211_X1 g0162(.A(new_n361), .B(new_n362), .C1(new_n340), .C2(new_n342), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n269), .A2(new_n243), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n360), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n340), .A2(new_n342), .ZN(new_n366));
  INV_X1    g0166(.A(new_n361), .ZN(new_n367));
  INV_X1    g0167(.A(new_n362), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n364), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(KEYINPUT75), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n365), .A2(new_n253), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G190), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n260), .A2(G232), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n374), .A2(new_n256), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(G200), .B1(new_n372), .B2(new_n375), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n359), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT17), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT17), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n359), .B(new_n380), .C1(new_n376), .C2(new_n377), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n343), .A2(KEYINPUT7), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(G68), .A3(new_n346), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(KEYINPUT16), .A3(new_n355), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(new_n358), .A3(new_n274), .ZN(new_n386));
  INV_X1    g0186(.A(new_n330), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n372), .A2(G179), .A3(new_n375), .ZN(new_n389));
  INV_X1    g0189(.A(G169), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n372), .B2(new_n375), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n388), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n388), .B(KEYINPUT18), .C1(new_n389), .C2(new_n391), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n382), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n278), .A2(G77), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n398), .B(KEYINPUT68), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n276), .A2(new_n240), .ZN(new_n400));
  XOR2_X1   g0200(.A(KEYINPUT15), .B(G87), .Z(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n271), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n268), .A2(new_n267), .B1(new_n209), .B2(new_n240), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n274), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n399), .A2(new_n400), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G244), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n256), .B1(new_n259), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT67), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G179), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n247), .A2(G232), .A3(new_n248), .ZN(new_n413));
  INV_X1    g0213(.A(G107), .ZN(new_n414));
  OAI221_X1 g0214(.A(new_n413), .B1(new_n414), .B2(new_n247), .C1(new_n250), .C2(new_n224), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n253), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n411), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT69), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n418), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n407), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n411), .A2(new_n416), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n390), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(G200), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n425), .B(new_n407), .C1(new_n373), .C2(new_n422), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n327), .A2(new_n397), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n247), .A2(G250), .A3(G1698), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G283), .ZN(new_n432));
  AND2_X1   g0232(.A1(KEYINPUT4), .A2(G244), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n337), .A2(new_n339), .A3(new_n433), .A4(new_n248), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n366), .A2(G244), .A3(new_n248), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT4), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT79), .B1(new_n438), .B2(new_n257), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT79), .ZN(new_n440));
  AOI21_X1  g0240(.A(G1698), .B1(new_n340), .B2(new_n342), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT4), .B1(new_n441), .B2(G244), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n440), .B(new_n253), .C1(new_n442), .C2(new_n435), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G41), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT65), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT65), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G41), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT5), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G45), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G1), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n450), .A2(KEYINPUT80), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT80), .B1(new_n450), .B2(new_n452), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n445), .A2(KEYINPUT5), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n455), .A2(G274), .A3(new_n257), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n450), .A2(new_n452), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT80), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n450), .A2(KEYINPUT80), .A3(new_n452), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(new_n456), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(G257), .A3(new_n257), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n444), .A2(KEYINPUT81), .A3(new_n412), .A4(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT81), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n439), .A2(new_n463), .A3(new_n457), .A4(new_n443), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n466), .B1(new_n467), .B2(G179), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n331), .B(new_n275), .C1(G1), .C2(new_n269), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n276), .A2(new_n298), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n469), .A2(new_n298), .B1(KEYINPUT78), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT76), .A2(KEYINPUT6), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(KEYINPUT76), .A2(KEYINPUT6), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n473), .A2(G97), .A3(new_n414), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT77), .ZN(new_n476));
  INV_X1    g0276(.A(new_n474), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(new_n472), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT77), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n478), .A2(new_n479), .A3(G97), .A4(new_n414), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n242), .B1(new_n472), .B2(new_n477), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n476), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G20), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n351), .A2(new_n353), .A3(G107), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n266), .A2(G77), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n471), .B1(new_n486), .B2(new_n274), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n470), .A2(KEYINPUT78), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n253), .B1(new_n442), .B2(new_n435), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n463), .A2(new_n457), .A3(new_n490), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n487), .A2(new_n489), .B1(new_n491), .B2(new_n390), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n465), .A2(new_n468), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n366), .A2(new_n209), .A3(G68), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT19), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT82), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT82), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT19), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n271), .B2(new_n298), .ZN(new_n500));
  AND2_X1   g0300(.A1(G33), .A2(G97), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n496), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n209), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n243), .A2(new_n298), .A3(new_n414), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n494), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n274), .ZN(new_n507));
  INV_X1    g0307(.A(new_n469), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n401), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n401), .A2(new_n275), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n248), .A2(G244), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G238), .A2(G1698), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n366), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n269), .A2(new_n218), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n257), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n257), .B(G250), .C1(G1), .C2(new_n451), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n452), .A2(G274), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n390), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n523), .ZN(new_n525));
  AOI211_X1 g0325(.A(new_n513), .B(new_n515), .C1(new_n340), .C2(new_n342), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n253), .B1(new_n526), .B2(new_n518), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n527), .A3(new_n412), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n512), .A2(new_n524), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n525), .A2(new_n527), .A3(G190), .ZN(new_n530));
  OAI21_X1  g0330(.A(G200), .B1(new_n520), .B2(new_n523), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n510), .B1(new_n506), .B2(new_n274), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n469), .A2(new_n243), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n530), .A2(new_n531), .A3(new_n532), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT83), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n529), .A2(new_n535), .A3(KEYINPUT83), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n467), .A2(G200), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n463), .A2(new_n457), .A3(new_n490), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G190), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n540), .A2(new_n489), .A3(new_n487), .A4(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n493), .A2(new_n538), .A3(new_n539), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n462), .A2(G270), .A3(new_n257), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n248), .A2(G264), .ZN(new_n546));
  NOR2_X1   g0346(.A1(G257), .A2(G1698), .ZN(new_n547));
  AOI211_X1 g0347(.A(new_n546), .B(new_n547), .C1(new_n340), .C2(new_n342), .ZN(new_n548));
  INV_X1    g0348(.A(G303), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n247), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n253), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n457), .A2(new_n545), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n508), .A2(G116), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n432), .B(new_n209), .C1(G33), .C2(new_n298), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n554), .B(new_n274), .C1(new_n209), .C2(G116), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT20), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n555), .A2(new_n556), .ZN(new_n558));
  OAI221_X1 g0358(.A(new_n553), .B1(G116), .B2(new_n275), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n552), .A2(new_n559), .A3(G169), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT21), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n559), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n457), .A2(new_n545), .A3(G190), .A4(new_n551), .ZN(new_n564));
  INV_X1    g0364(.A(new_n552), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n563), .B(new_n564), .C1(new_n565), .C2(new_n284), .ZN(new_n566));
  AND4_X1   g0366(.A1(G179), .A2(new_n457), .A3(new_n545), .A4(new_n551), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n559), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n552), .A2(new_n559), .A3(KEYINPUT21), .A4(G169), .ZN(new_n569));
  AND4_X1   g0369(.A1(new_n562), .A2(new_n566), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n462), .A2(G264), .A3(new_n257), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n248), .A2(G257), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G250), .A2(G1698), .ZN(new_n573));
  AOI211_X1 g0373(.A(new_n572), .B(new_n573), .C1(new_n340), .C2(new_n342), .ZN(new_n574));
  INV_X1    g0374(.A(G294), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n269), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n253), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n457), .A2(new_n571), .A3(new_n577), .ZN(new_n578));
  OR2_X1    g0378(.A1(new_n578), .A2(new_n412), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT86), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(KEYINPUT86), .B(new_n253), .C1(new_n574), .C2(new_n576), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n583), .A2(new_n457), .A3(new_n571), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n579), .B1(new_n584), .B2(new_n390), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n270), .A2(G116), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n209), .A2(G107), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n587), .B(KEYINPUT23), .ZN(new_n588));
  NAND2_X1  g0388(.A1(KEYINPUT22), .A2(G87), .ZN(new_n589));
  AOI211_X1 g0389(.A(G20), .B(new_n589), .C1(new_n340), .C2(new_n342), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT84), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n337), .A2(new_n339), .A3(new_n209), .A4(G87), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT22), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n590), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n589), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n366), .A2(new_n209), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n592), .A2(new_n593), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT84), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n586), .B(new_n588), .C1(new_n595), .C2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT24), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n591), .B1(new_n590), .B2(new_n594), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n597), .A2(KEYINPUT84), .A3(new_n598), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n605), .A2(KEYINPUT24), .A3(new_n586), .A4(new_n588), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n602), .A2(new_n274), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT25), .B1(new_n275), .B2(G107), .ZN(new_n608));
  OR3_X1    g0408(.A1(new_n275), .A2(KEYINPUT25), .A3(G107), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n608), .B(new_n609), .C1(new_n469), .C2(new_n414), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT85), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n585), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n583), .A2(new_n373), .A3(new_n457), .A4(new_n571), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n578), .A2(new_n284), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n616), .A2(new_n611), .A3(new_n607), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n570), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n430), .A2(new_n544), .A3(new_n618), .ZN(G372));
  AOI21_X1  g0419(.A(new_n515), .B1(new_n340), .B2(new_n342), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n518), .B1(new_n620), .B2(new_n514), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT87), .B1(new_n621), .B2(new_n257), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT87), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n623), .B(new_n253), .C1(new_n526), .C2(new_n518), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n523), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n528), .B(new_n512), .C1(new_n625), .C2(G169), .ZN(new_n626));
  AOI211_X1 g0426(.A(new_n510), .B(new_n533), .C1(new_n506), .C2(new_n274), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n530), .B(new_n627), .C1(new_n625), .C2(new_n284), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n493), .A2(new_n617), .A3(new_n629), .A4(new_n543), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n562), .A2(new_n568), .A3(new_n569), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT88), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT88), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n562), .A2(new_n633), .A3(new_n568), .A4(new_n569), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n632), .A2(new_n613), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n538), .A2(new_n539), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT26), .B1(new_n637), .B2(new_n493), .ZN(new_n638));
  INV_X1    g0438(.A(new_n626), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n626), .A2(new_n628), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n493), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n636), .A2(new_n638), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n429), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n292), .ZN(new_n646));
  INV_X1    g0446(.A(new_n424), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n647), .A2(new_n326), .B1(new_n322), .B2(new_n310), .ZN(new_n648));
  INV_X1    g0448(.A(new_n382), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n396), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n646), .B1(new_n650), .B2(new_n289), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n645), .A2(new_n651), .ZN(G369));
  NAND2_X1  g0452(.A1(new_n632), .A2(new_n634), .ZN(new_n653));
  INV_X1    g0453(.A(G13), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(G20), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n213), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n653), .A2(new_n559), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n661), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n570), .B1(new_n563), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G330), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n612), .A2(new_n661), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n613), .A2(new_n669), .A3(new_n617), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT89), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT89), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n613), .A2(new_n669), .A3(new_n672), .A4(new_n617), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n613), .A2(new_n663), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n668), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n585), .A2(new_n612), .A3(new_n663), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n562), .A2(new_n568), .A3(new_n569), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n661), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n671), .A2(new_n673), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n678), .A2(new_n679), .A3(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n214), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n255), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n504), .A2(G116), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G1), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n206), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n644), .A2(KEYINPUT93), .A3(new_n663), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT93), .B1(new_n644), .B2(new_n663), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n691), .A2(new_n692), .A3(KEYINPUT29), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT29), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n642), .B1(new_n637), .B2(new_n493), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n465), .A2(new_n468), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(KEYINPUT26), .A3(new_n492), .A4(new_n629), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT94), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n493), .A2(new_n543), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n617), .A2(new_n629), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n613), .A2(new_n680), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n641), .A2(KEYINPUT94), .A3(KEYINPUT26), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n699), .A2(new_n626), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n694), .B1(new_n705), .B2(new_n663), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n693), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n571), .A2(new_n527), .A3(new_n525), .A4(new_n577), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT90), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n520), .A2(new_n523), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(KEYINPUT90), .A3(new_n577), .A4(new_n571), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n710), .A2(new_n567), .A3(new_n541), .A4(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(KEYINPUT91), .B1(new_n467), .B2(new_n578), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n716), .A2(new_n565), .A3(new_n625), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n467), .A2(KEYINPUT91), .A3(new_n578), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n718), .A2(new_n412), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n715), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT92), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n713), .A2(new_n721), .A3(new_n714), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n713), .B2(new_n714), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n661), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n618), .A2(new_n544), .A3(new_n661), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n713), .A2(new_n714), .ZN(new_n730));
  AOI211_X1 g0530(.A(new_n728), .B(new_n663), .C1(new_n720), .C2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n667), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n707), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n690), .B1(new_n736), .B2(G1), .ZN(G364));
  AOI21_X1  g0537(.A(new_n213), .B1(new_n655), .B2(G45), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n685), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n668), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(G330), .B2(new_n665), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n208), .B1(G20), .B2(new_n390), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n366), .A2(new_n684), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n207), .A2(new_n451), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n748), .B(new_n749), .C1(new_n241), .C2(new_n451), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n247), .A2(new_n214), .ZN(new_n751));
  XOR2_X1   g0551(.A(G355), .B(KEYINPUT95), .Z(new_n752));
  OAI221_X1 g0552(.A(new_n750), .B1(G116), .B2(new_n214), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n209), .A2(new_n412), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n373), .A2(new_n284), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n247), .B1(new_n757), .B2(G326), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n209), .A2(G179), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n758), .B1(new_n549), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n284), .A2(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n754), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT33), .B(G317), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n761), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G190), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n754), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G311), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n759), .A2(new_n762), .ZN(new_n770));
  INV_X1    g0570(.A(G283), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n768), .A2(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n759), .A2(new_n767), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n774), .A2(G329), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n754), .A2(G190), .A3(new_n284), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n772), .B(new_n775), .C1(G322), .C2(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n373), .A2(G179), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n209), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n766), .B(new_n778), .C1(new_n575), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n770), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G107), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n783), .B(new_n247), .C1(new_n243), .C2(new_n760), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT97), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT96), .B(G159), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n774), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT32), .Z(new_n788));
  NOR2_X1   g0588(.A1(new_n780), .A2(new_n298), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n776), .A2(new_n332), .B1(new_n763), .B2(new_n223), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n789), .B(new_n790), .C1(G50), .C2(new_n757), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n785), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n768), .A2(new_n240), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n781), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n747), .A2(new_n753), .B1(new_n794), .B2(new_n746), .ZN(new_n795));
  INV_X1    g0595(.A(new_n745), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n740), .B(new_n795), .C1(new_n665), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n742), .A2(new_n797), .ZN(G396));
  XNOR2_X1  g0598(.A(new_n417), .B(new_n418), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n799), .A2(new_n423), .A3(new_n406), .A4(new_n661), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT100), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n421), .A2(KEYINPUT100), .A3(new_n423), .A4(new_n661), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n406), .A2(new_n661), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT99), .Z(new_n806));
  NAND3_X1  g0606(.A1(new_n424), .A2(new_n426), .A3(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n691), .B2(new_n692), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n804), .A2(new_n807), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n644), .A2(new_n663), .A3(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n740), .B1(new_n812), .B2(new_n733), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT101), .Z(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n733), .B2(new_n812), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n366), .B1(new_n332), .B2(new_n780), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n782), .A2(G68), .ZN(new_n817));
  INV_X1    g0617(.A(G132), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n818), .B2(new_n773), .ZN(new_n819));
  INV_X1    g0619(.A(new_n768), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G137), .A2(new_n757), .B1(new_n820), .B2(new_n786), .ZN(new_n821));
  INV_X1    g0621(.A(G143), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n822), .B2(new_n776), .C1(new_n265), .C2(new_n763), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT34), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n816), .B(new_n819), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n825), .B1(new_n824), .B2(new_n823), .C1(new_n202), .C2(new_n760), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n760), .A2(new_n414), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n776), .A2(new_n575), .B1(new_n773), .B2(new_n769), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n827), .B(new_n828), .C1(G116), .C2(new_n820), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n247), .B(new_n789), .C1(G303), .C2(new_n757), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n763), .A2(KEYINPUT98), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n763), .A2(KEYINPUT98), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(G283), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n782), .A2(G87), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n829), .A2(new_n830), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n826), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n746), .A2(new_n743), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n838), .A2(new_n746), .B1(new_n240), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n740), .B(new_n840), .C1(new_n810), .C2(new_n744), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n815), .A2(new_n841), .ZN(G384));
  INV_X1    g0642(.A(new_n391), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n372), .A2(G179), .A3(new_n375), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(new_n659), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n388), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT37), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n846), .A2(new_n847), .A3(new_n378), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n348), .B1(KEYINPUT16), .B2(new_n347), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n387), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n845), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n847), .B1(new_n852), .B2(new_n378), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n659), .ZN(new_n856));
  AND4_X1   g0656(.A1(KEYINPUT103), .A2(new_n397), .A3(new_n856), .A4(new_n851), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n659), .B1(new_n382), .B2(new_n396), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT103), .B1(new_n858), .B2(new_n851), .ZN(new_n859));
  OAI211_X1 g0659(.A(KEYINPUT38), .B(new_n855), .C1(new_n857), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n858), .A2(new_n388), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n847), .B1(new_n846), .B2(new_n378), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n849), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n861), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT40), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n322), .A2(new_n661), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n323), .A2(new_n868), .A3(new_n326), .ZN(new_n869));
  INV_X1    g0669(.A(new_n326), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n322), .B(new_n661), .C1(new_n310), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n663), .B1(new_n720), .B2(new_n724), .ZN(new_n873));
  INV_X1    g0673(.A(new_n544), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n613), .A2(new_n617), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n874), .A2(new_n875), .A3(new_n570), .A4(new_n663), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n873), .B1(new_n876), .B2(KEYINPUT31), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n726), .A2(new_n728), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n810), .B(new_n872), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n867), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT104), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n397), .A2(new_n856), .A3(new_n851), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT103), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n858), .A2(KEYINPUT103), .A3(new_n851), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n886), .B2(new_n855), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n861), .B(new_n854), .C1(new_n884), .C2(new_n885), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n881), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n855), .B1(new_n857), .B2(new_n859), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n861), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(KEYINPUT104), .A3(new_n860), .ZN(new_n892));
  INV_X1    g0692(.A(new_n879), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n880), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n873), .A2(KEYINPUT31), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n729), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n429), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n896), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(G330), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT39), .B1(new_n887), .B2(new_n888), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n323), .A2(new_n661), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n647), .A2(KEYINPUT102), .A3(new_n663), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n647), .A2(new_n663), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT102), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n811), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n889), .A2(new_n892), .A3(new_n872), .A4(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n394), .A2(new_n395), .A3(new_n659), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n907), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n429), .B1(new_n693), .B2(new_n706), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n651), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n915), .B(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n902), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n902), .A2(new_n918), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n919), .B1(new_n921), .B2(KEYINPUT105), .ZN(new_n922));
  OAI221_X1 g0722(.A(new_n922), .B1(KEYINPUT105), .B2(new_n921), .C1(new_n213), .C2(new_n655), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n218), .B1(new_n482), .B2(KEYINPUT35), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n924), .B(new_n210), .C1(KEYINPUT35), .C2(new_n482), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT36), .ZN(new_n926));
  OAI21_X1  g0726(.A(G77), .B1(new_n332), .B2(new_n223), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n927), .A2(new_n206), .B1(G50), .B2(new_n223), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(G1), .A3(new_n654), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n923), .A2(new_n926), .A3(new_n929), .ZN(G367));
  NOR2_X1   g0730(.A1(new_n627), .A2(new_n663), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT106), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n639), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n640), .B2(new_n932), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n487), .A2(new_n489), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n661), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n493), .A2(new_n543), .A3(new_n937), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n465), .A2(new_n468), .A3(new_n492), .A4(new_n661), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT107), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n938), .A2(KEYINPUT107), .A3(new_n939), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n682), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT42), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n942), .A2(new_n943), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(new_n585), .A3(new_n612), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n661), .B1(new_n949), .B2(new_n493), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n935), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n678), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n952), .A3(new_n948), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n935), .B1(new_n678), .B2(new_n944), .C1(new_n947), .C2(new_n950), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n954), .B1(new_n953), .B2(new_n955), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n685), .B(KEYINPUT41), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT109), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n682), .A2(new_n679), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n962), .A2(new_n944), .A3(KEYINPUT44), .ZN(new_n963));
  AOI21_X1  g0763(.A(KEYINPUT44), .B1(new_n962), .B2(new_n944), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n962), .B2(new_n944), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n948), .A2(new_n679), .A3(new_n682), .A4(new_n966), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n961), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n968), .A2(new_n969), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n962), .A2(new_n944), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT44), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n962), .A2(new_n944), .A3(KEYINPUT44), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n972), .A2(new_n977), .A3(KEYINPUT109), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n971), .A2(new_n978), .A3(new_n952), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n972), .A2(new_n977), .ZN(new_n980));
  OAI21_X1  g0780(.A(KEYINPUT110), .B1(new_n980), .B2(new_n952), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n677), .A2(new_n681), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n682), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n668), .A2(KEYINPUT111), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n983), .A2(new_n682), .B1(new_n668), .B2(KEYINPUT111), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n986), .B1(new_n987), .B2(new_n985), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n735), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n971), .A2(new_n978), .A3(KEYINPUT110), .A4(new_n952), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n982), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n960), .B1(new_n991), .B2(new_n736), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n958), .B1(new_n992), .B2(new_n739), .ZN(new_n993));
  INV_X1    g0793(.A(new_n740), .ZN(new_n994));
  INV_X1    g0794(.A(new_n760), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(G116), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT46), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n996), .A2(new_n997), .B1(new_n414), .B2(new_n780), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G311), .B2(new_n757), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n366), .B1(new_n996), .B2(new_n997), .ZN(new_n1000));
  INV_X1    g0800(.A(G317), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n776), .A2(new_n549), .B1(new_n773), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n770), .A2(new_n298), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AND3_X1   g0804(.A1(new_n999), .A2(new_n1000), .A3(new_n1004), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n771), .B2(new_n768), .C1(new_n575), .C2(new_n833), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n770), .A2(new_n240), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n834), .A2(new_n786), .ZN(new_n1008));
  INV_X1    g0808(.A(G137), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n760), .A2(new_n332), .B1(new_n773), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G50), .B2(new_n820), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n352), .B1(new_n777), .B2(G150), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n780), .A2(new_n223), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G143), .B2(new_n757), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1008), .A2(new_n1011), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1006), .B1(new_n1007), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT47), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n994), .B1(new_n1017), .B2(new_n746), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n748), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n747), .B1(new_n214), .B2(new_n402), .C1(new_n236), .C2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT112), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1018), .B(new_n1021), .C1(new_n796), .C2(new_n934), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n993), .A2(new_n1022), .ZN(G387));
  INV_X1    g0823(.A(KEYINPUT113), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n735), .A2(new_n988), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n989), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n735), .A2(KEYINPUT113), .A3(new_n988), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1027), .A2(new_n685), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n988), .A2(new_n738), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n774), .A2(G326), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G322), .A2(new_n757), .B1(new_n820), .B2(G303), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n1001), .B2(new_n776), .C1(new_n833), .C2(new_n769), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT48), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n771), .B2(new_n780), .C1(new_n575), .C2(new_n760), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT49), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n366), .B(new_n1031), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n1036), .B2(new_n1035), .C1(new_n218), .C2(new_n770), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n366), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n777), .A2(G50), .B1(new_n995), .B2(G77), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n223), .B2(new_n768), .C1(new_n265), .C2(new_n773), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n780), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n401), .ZN(new_n1043));
  INV_X1    g0843(.A(G159), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1043), .B1(new_n1044), .B2(new_n756), .C1(new_n268), .C2(new_n763), .ZN(new_n1045));
  OR4_X1    g0845(.A1(new_n1039), .A2(new_n1041), .A3(new_n1003), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1038), .A2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g0847(.A(G116), .B(new_n504), .C1(G68), .C2(G77), .ZN(new_n1048));
  OR3_X1    g0848(.A1(new_n268), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1049));
  OAI21_X1  g0849(.A(KEYINPUT50), .B1(new_n268), .B2(G50), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n451), .A4(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1019), .B1(new_n233), .B2(G45), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n751), .A2(new_n687), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(G107), .B2(new_n214), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1047), .A2(new_n746), .B1(new_n747), .B2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1056), .B(new_n740), .C1(new_n677), .C2(new_n796), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1029), .A2(new_n1030), .A3(new_n1057), .ZN(G393));
  XNOR2_X1  g0858(.A(new_n980), .B(new_n678), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n991), .B(new_n685), .C1(new_n989), .C2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n944), .A2(new_n745), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G294), .A2(new_n820), .B1(new_n774), .B2(G322), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n218), .B2(new_n780), .C1(new_n771), .C2(new_n760), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G303), .B2(new_n834), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n776), .A2(new_n769), .B1(new_n756), .B2(new_n1001), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT52), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1064), .A2(new_n352), .A3(new_n783), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1042), .A2(G77), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1068), .B(new_n366), .C1(new_n268), .C2(new_n768), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G50), .B2(new_n834), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n776), .A2(new_n1044), .B1(new_n756), .B2(new_n265), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT51), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n760), .A2(new_n223), .B1(new_n773), .B2(new_n822), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT114), .Z(new_n1074));
  NAND4_X1  g0874(.A1(new_n1070), .A2(new_n836), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1067), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n994), .B1(new_n1076), .B2(new_n746), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1061), .A2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n245), .A2(new_n748), .B1(G97), .B2(new_n684), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1078), .B1(new_n747), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n1059), .B2(new_n739), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1060), .A2(new_n1081), .ZN(G390));
  NAND3_X1  g0882(.A1(new_n898), .A2(G330), .A3(new_n810), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n872), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n705), .A2(new_n663), .A3(new_n810), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n909), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n667), .B(new_n808), .C1(new_n729), .C2(new_n732), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n1088), .B2(new_n872), .ZN(new_n1089));
  OAI211_X1 g0889(.A(G330), .B(new_n810), .C1(new_n877), .C2(new_n731), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n1084), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n898), .A2(G330), .A3(new_n810), .A4(new_n872), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1085), .A2(new_n1089), .B1(new_n1093), .B2(new_n912), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n429), .A2(G330), .A3(new_n898), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n916), .A2(new_n651), .A3(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n906), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n866), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1084), .B1(new_n1086), .B2(new_n909), .ZN(new_n1100));
  OAI21_X1  g0900(.A(KEYINPUT115), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1087), .A2(new_n872), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT115), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n906), .B1(new_n860), .B2(new_n865), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1090), .A2(new_n1084), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n912), .A2(new_n872), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n1098), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(new_n904), .A3(new_n903), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n1106), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1092), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1113));
  OR3_X1    g0913(.A1(new_n1097), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1097), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n685), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n903), .A2(new_n743), .A3(new_n904), .ZN(new_n1117));
  INV_X1    g0917(.A(G128), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n247), .B1(new_n756), .B2(new_n1118), .C1(new_n780), .C2(new_n1044), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT54), .B(G143), .Z(new_n1120));
  AOI21_X1  g0920(.A(new_n1119), .B1(new_n820), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n995), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT53), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n760), .B2(new_n265), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G50), .A2(new_n782), .B1(new_n774), .B2(G125), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1121), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1127), .B1(new_n818), .B2(new_n776), .C1(new_n1009), .C2(new_n833), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n352), .B1(new_n760), .B2(new_n243), .C1(new_n771), .C2(new_n756), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n817), .B1(new_n298), .B2(new_n768), .C1(new_n218), .C2(new_n776), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G294), .B2(new_n774), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1131), .B(new_n1068), .C1(new_n414), .C2(new_n833), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1128), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1133), .A2(new_n746), .B1(new_n268), .B2(new_n839), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1117), .A2(new_n740), .A3(new_n1134), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n1136), .B2(new_n739), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1137), .A2(KEYINPUT116), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT116), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1139), .B(new_n1135), .C1(new_n1136), .C2(new_n739), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1116), .B1(new_n1138), .B2(new_n1140), .ZN(G378));
  NAND3_X1  g0941(.A1(new_n907), .A2(new_n913), .A3(new_n914), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT55), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n294), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n293), .A2(KEYINPUT55), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n281), .A2(new_n659), .ZN(new_n1146));
  OR3_X1    g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1146), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1147), .A2(new_n1150), .A3(new_n1148), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n896), .A2(G330), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1154), .B1(new_n896), .B2(G330), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1142), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n894), .A2(new_n895), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n880), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(G330), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1154), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n896), .A2(G330), .A3(new_n1154), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n915), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n738), .B1(new_n1157), .B2(new_n1164), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n366), .A2(new_n255), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n782), .A2(G58), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n240), .B2(new_n760), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1166), .B(new_n1168), .C1(G283), .C2(new_n774), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT118), .Z(new_n1170));
  OAI22_X1  g0970(.A1(new_n756), .A2(new_n218), .B1(new_n763), .B2(new_n298), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1013), .B(new_n1171), .C1(G107), .C2(new_n777), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(new_n402), .C2(new_n768), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT58), .Z(new_n1174));
  OAI22_X1  g0974(.A1(new_n776), .A2(new_n1118), .B1(new_n768), .B2(new_n1009), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n995), .B2(new_n1120), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G125), .A2(new_n757), .B1(new_n764), .B2(G132), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(new_n265), .C2(new_n780), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1178), .A2(KEYINPUT59), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n774), .A2(G124), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(KEYINPUT59), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(G33), .A2(G41), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT117), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n782), .B2(new_n786), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .A4(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1166), .A2(new_n202), .A3(new_n1183), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n746), .B1(new_n1174), .B2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT119), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n994), .B1(new_n202), .B2(new_n839), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT120), .Z(new_n1191));
  OAI211_X1 g0991(.A(new_n1189), .B(new_n1191), .C1(new_n1154), .C2(new_n744), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT122), .ZN(new_n1193));
  OAI21_X1  g0993(.A(KEYINPUT123), .B1(new_n1165), .B2(new_n1193), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1155), .A2(new_n1156), .A3(new_n1142), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n915), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n739), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT123), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1193), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1194), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1096), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1115), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT57), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1203), .B(KEYINPUT57), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n685), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1201), .A2(new_n1208), .ZN(G375));
  NAND2_X1  g1009(.A1(new_n1084), .A2(new_n743), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n366), .B1(new_n202), .B2(new_n780), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1167), .B1(new_n265), .B2(new_n768), .C1(new_n1044), .C2(new_n760), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(G128), .C2(new_n774), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT124), .Z(new_n1214));
  AOI22_X1  g1014(.A1(new_n834), .A2(new_n1120), .B1(G132), .B2(new_n757), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(new_n1009), .C2(new_n776), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n760), .A2(new_n298), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n776), .A2(new_n771), .B1(new_n768), .B2(new_n414), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(G303), .C2(new_n774), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n247), .B(new_n1007), .C1(G294), .C2(new_n757), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n834), .A2(G116), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1219), .A2(new_n1043), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1216), .A2(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1223), .A2(new_n746), .B1(new_n223), .B2(new_n839), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1210), .A2(new_n740), .A3(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1094), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1225), .B1(new_n1226), .B2(new_n739), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n959), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1227), .B1(new_n1229), .B2(new_n1097), .ZN(G381));
  XNOR2_X1  g1030(.A(G375), .B(KEYINPUT125), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1116), .A2(new_n1137), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(G390), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(G396), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1029), .A2(new_n1236), .A3(new_n1030), .A4(new_n1057), .ZN(new_n1237));
  OR4_X1    g1037(.A1(G384), .A2(G387), .A3(G381), .A4(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1235), .A2(new_n1238), .ZN(G407));
  INV_X1    g1039(.A(G213), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n1233), .B2(new_n660), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1238), .B2(new_n1235), .ZN(G409));
  NAND2_X1  g1042(.A1(G393), .A2(G396), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1243), .A2(new_n1237), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n993), .A2(new_n1022), .A3(G390), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G390), .B1(new_n993), .B2(new_n1022), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1244), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G387), .A2(new_n1234), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n993), .A2(G390), .A3(new_n1022), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT126), .B1(new_n1243), .B2(new_n1237), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1245), .A2(KEYINPUT126), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1247), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1253), .A2(KEYINPUT61), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1240), .A2(G343), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1201), .A2(new_n1208), .A3(G378), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1199), .B(new_n1197), .C1(new_n1204), .C2(new_n960), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1232), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1255), .B1(new_n1256), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(G384), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT60), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n686), .B1(new_n1228), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1226), .A2(new_n1202), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1263), .B(new_n1264), .C1(new_n1262), .C2(new_n1228), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1227), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1261), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(G384), .A2(new_n1227), .A3(new_n1265), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1260), .A2(KEYINPUT63), .A3(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT63), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1255), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1255), .A2(G2897), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1268), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G384), .B1(new_n1265), .B2(new_n1227), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1277), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1267), .A2(new_n1268), .A3(new_n1276), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1272), .B1(new_n1275), .B2(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1275), .A2(new_n1269), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1254), .B(new_n1271), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1260), .A2(new_n1287), .A3(new_n1270), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1289), .B1(new_n1260), .B2(new_n1282), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1287), .B1(new_n1260), .B2(new_n1270), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1288), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1253), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1286), .B1(new_n1292), .B2(new_n1293), .ZN(G405));
  AND3_X1   g1094(.A1(new_n1201), .A2(new_n1208), .A3(G378), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1232), .B1(new_n1201), .B2(new_n1208), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1270), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G375), .A2(new_n1258), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(new_n1256), .A3(new_n1269), .ZN(new_n1299));
  AOI211_X1 g1099(.A(KEYINPUT127), .B(new_n1253), .C1(new_n1297), .C2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT127), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1301), .B1(new_n1302), .B2(new_n1293), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1293), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1300), .A2(new_n1303), .A3(new_n1304), .ZN(G402));
endmodule


