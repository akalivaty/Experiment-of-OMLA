//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n586, new_n587,
    new_n588, new_n589, new_n591, new_n592, new_n594, new_n595, new_n596,
    new_n597, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G22gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(G141gat), .B(G148gat), .ZN(new_n207));
  XOR2_X1   g006(.A(G155gat), .B(G162gat), .Z(new_n208));
  INV_X1    g007(.A(G155gat), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT2), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI211_X1 g010(.A(new_n207), .B(new_n208), .C1(KEYINPUT76), .C2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(KEYINPUT76), .B2(new_n211), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n211), .A2(KEYINPUT75), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n214), .A2(new_n207), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n211), .A2(KEYINPUT75), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n208), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G197gat), .B(G204gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n219), .A2(KEYINPUT72), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(KEYINPUT72), .ZN(new_n221));
  AND2_X1   g020(.A1(G211gat), .A2(G218gat), .ZN(new_n222));
  OAI22_X1  g021(.A1(new_n220), .A2(new_n221), .B1(KEYINPUT22), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(new_n223), .B(KEYINPUT73), .Z(new_n224));
  XOR2_X1   g023(.A(G211gat), .B(G218gat), .Z(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n223), .B(KEYINPUT73), .ZN(new_n227));
  INV_X1    g026(.A(new_n225), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT29), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n226), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n218), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT79), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n233), .A2(new_n234), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n226), .A2(new_n229), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT29), .B1(new_n218), .B2(new_n232), .ZN(new_n239));
  OAI22_X1  g038(.A1(new_n235), .A2(new_n236), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(G228gat), .A2(G233gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n218), .A2(new_n232), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(new_n230), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n239), .A2(KEYINPUT80), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n238), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n249), .A2(new_n242), .A3(new_n233), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n206), .B1(new_n243), .B2(new_n251), .ZN(new_n252));
  AOI211_X1 g051(.A(G22gat), .B(new_n250), .C1(new_n240), .C2(new_n242), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n205), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT81), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n243), .A2(new_n251), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G22gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n206), .A3(new_n251), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n259), .A3(new_n204), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT82), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT82), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n258), .A2(new_n262), .A3(new_n259), .A4(new_n204), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT83), .B1(new_n256), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n261), .A2(new_n263), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n254), .B(KEYINPUT81), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT83), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT27), .B(G183gat), .ZN(new_n272));
  INV_X1    g071(.A(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n274), .B(new_n275), .Z(new_n276));
  OR2_X1    g075(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n278));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(KEYINPUT26), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT26), .ZN(new_n282));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G183gat), .ZN(new_n285));
  OAI22_X1  g084(.A1(new_n281), .A2(new_n284), .B1(new_n285), .B2(new_n273), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n276), .A2(new_n277), .B1(new_n278), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(new_n278), .B2(new_n286), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n279), .A2(KEYINPUT23), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(KEYINPUT64), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT23), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n283), .B1(new_n280), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n285), .A2(new_n273), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(new_n295), .B2(KEYINPUT24), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT65), .B(KEYINPUT24), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n296), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n293), .A2(KEYINPUT25), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n296), .B1(KEYINPUT24), .B2(new_n295), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n299), .B1(new_n301), .B2(KEYINPUT25), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n288), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n230), .ZN(new_n304));
  NAND2_X1  g103(.A1(G226gat), .A2(G233gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n288), .A2(new_n302), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n306), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(new_n237), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT74), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n237), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n312), .B1(new_n308), .B2(new_n237), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G8gat), .B(G36gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(G64gat), .B(G92gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n318), .A2(KEYINPUT30), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n314), .A2(new_n317), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(KEYINPUT30), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(G113gat), .B(G120gat), .Z(new_n323));
  INV_X1    g122(.A(KEYINPUT68), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G127gat), .B(G134gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT1), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n327), .B(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n213), .A2(new_n217), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n331), .B1(new_n332), .B2(KEYINPUT3), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n244), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n332), .A2(new_n330), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n334), .B1(KEYINPUT4), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(KEYINPUT77), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(KEYINPUT4), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT5), .ZN(new_n339));
  NAND2_X1  g138(.A1(G225gat), .A2(G233gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n341), .A2(KEYINPUT78), .ZN(new_n342));
  INV_X1    g141(.A(new_n337), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n218), .B2(new_n331), .ZN(new_n344));
  INV_X1    g143(.A(new_n340), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n345), .B1(new_n335), .B2(KEYINPUT4), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n334), .B(new_n347), .C1(new_n337), .C2(KEYINPUT4), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(KEYINPUT5), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n341), .A2(KEYINPUT78), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n342), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G1gat), .B(G29gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT0), .ZN(new_n353));
  XNOR2_X1  g152(.A(G57gat), .B(G85gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n353), .B(new_n354), .Z(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT6), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n342), .A2(new_n355), .A3(new_n349), .A4(new_n350), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n351), .A2(KEYINPUT6), .A3(new_n356), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n322), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n271), .A2(new_n363), .ZN(new_n364));
  OR2_X1    g163(.A1(new_n314), .A2(KEYINPUT37), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n314), .A2(KEYINPUT37), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(new_n317), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT84), .B1(new_n367), .B2(KEYINPUT38), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT38), .ZN(new_n369));
  INV_X1    g168(.A(new_n311), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT37), .B1(new_n370), .B2(new_n309), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n365), .A2(new_n369), .A3(new_n317), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n318), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n368), .A2(new_n362), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n367), .A2(KEYINPUT84), .A3(KEYINPUT38), .ZN(new_n375));
  INV_X1    g174(.A(new_n322), .ZN(new_n376));
  OR2_X1    g175(.A1(new_n338), .A2(new_n340), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n377), .B(KEYINPUT39), .C1(new_n345), .C2(new_n344), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n378), .B(new_n355), .C1(KEYINPUT39), .C2(new_n377), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT40), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n380), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n381), .A2(new_n357), .A3(new_n382), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n374), .A2(new_n375), .B1(new_n376), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n270), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT69), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n307), .B2(new_n331), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n307), .A2(new_n331), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n389), .B1(KEYINPUT69), .B2(new_n388), .ZN(new_n390));
  NAND2_X1  g189(.A1(G227gat), .A2(G233gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT34), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n393), .B1(new_n391), .B2(KEYINPUT71), .ZN(new_n394));
  OR2_X1    g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n394), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT70), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  XOR2_X1   g199(.A(G15gat), .B(G43gat), .Z(new_n401));
  XNOR2_X1  g200(.A(G71gat), .B(G99gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n390), .A2(new_n391), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n403), .B1(new_n404), .B2(KEYINPUT33), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT32), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OR2_X1    g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n405), .A2(new_n407), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n400), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n399), .A2(new_n409), .A3(new_n408), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT36), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n395), .A2(new_n396), .ZN(new_n415));
  INV_X1    g214(.A(new_n409), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n405), .A2(new_n407), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n408), .A2(new_n409), .A3(new_n397), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n414), .B1(KEYINPUT36), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n364), .A2(new_n385), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT35), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n413), .B1(new_n265), .B2(new_n269), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n319), .A2(new_n321), .B1(new_n360), .B2(new_n361), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n420), .A3(new_n425), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(new_n265), .B2(new_n269), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n424), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(G43gat), .B(G50gat), .Z(new_n432));
  INV_X1    g231(.A(KEYINPUT89), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT15), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  OR3_X1    g235(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT90), .ZN(new_n440));
  INV_X1    g239(.A(G29gat), .ZN(new_n441));
  INV_X1    g240(.A(G36gat), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n436), .B(new_n440), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(KEYINPUT91), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT88), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n437), .B1(new_n445), .B2(new_n438), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n438), .A2(new_n445), .ZN(new_n447));
  OAI22_X1  g246(.A1(new_n446), .A2(new_n447), .B1(new_n441), .B2(new_n442), .ZN(new_n448));
  INV_X1    g247(.A(new_n432), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(KEYINPUT15), .A3(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G15gat), .B(G22gat), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n452), .A2(G1gat), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT16), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n452), .B1(new_n454), .B2(G1gat), .ZN(new_n455));
  INV_X1    g254(.A(G8gat), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n453), .A2(new_n455), .B1(KEYINPUT92), .B2(new_n456), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n456), .A2(KEYINPUT92), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n457), .B(new_n458), .Z(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n451), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n451), .A2(new_n460), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n461), .B1(new_n462), .B2(KEYINPUT93), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(KEYINPUT93), .B2(new_n461), .ZN(new_n464));
  NAND2_X1  g263(.A1(G229gat), .A2(G233gat), .ZN(new_n465));
  XOR2_X1   g264(.A(new_n465), .B(KEYINPUT13), .Z(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n444), .A2(new_n450), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT17), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n462), .B1(new_n469), .B2(new_n460), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n470), .A2(KEYINPUT18), .A3(new_n465), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  XOR2_X1   g271(.A(G169gat), .B(G197gat), .Z(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G113gat), .B(G141gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(KEYINPUT86), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n475), .B(new_n477), .Z(new_n478));
  XNOR2_X1  g277(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n479));
  XOR2_X1   g278(.A(new_n478), .B(new_n479), .Z(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT18), .B1(new_n470), .B2(new_n465), .ZN(new_n482));
  OR3_X1    g281(.A1(new_n472), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n472), .B2(new_n482), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(G232gat), .A2(G233gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(KEYINPUT41), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(KEYINPUT99), .ZN(new_n488));
  XOR2_X1   g287(.A(G134gat), .B(G162gat), .Z(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT101), .ZN(new_n491));
  NAND2_X1  g290(.A1(G99gat), .A2(G106gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT8), .ZN(new_n493));
  OR2_X1    g292(.A1(G85gat), .A2(G92gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT100), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(G85gat), .A3(G92gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT7), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT7), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n496), .A2(new_n499), .A3(G85gat), .A4(G92gat), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n495), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G99gat), .B(G106gat), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n491), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n498), .A2(new_n500), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n493), .A2(new_n494), .ZN(new_n505));
  AND4_X1   g304(.A1(new_n491), .A2(new_n504), .A3(new_n502), .A4(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT102), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n505), .ZN(new_n508));
  INV_X1    g307(.A(new_n502), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT101), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT102), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n501), .A2(new_n491), .A3(new_n502), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n508), .A2(new_n509), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n507), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n469), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n515), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n468), .A2(new_n517), .B1(KEYINPUT41), .B2(new_n486), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G190gat), .B(G218gat), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT103), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n490), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n519), .B(new_n520), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n524), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G57gat), .B(G64gat), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(G71gat), .A2(G78gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(G71gat), .A2(G78gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(KEYINPUT94), .A2(KEYINPUT9), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n531), .B(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n459), .B1(KEYINPUT21), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT96), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n538), .B(KEYINPUT97), .Z(new_n539));
  INV_X1    g338(.A(new_n536), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G231gat), .A2(G233gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G127gat), .B(G155gat), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n539), .B(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G183gat), .B(G211gat), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT98), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n549), .B(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n528), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT10), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT105), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n502), .B1(new_n508), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(new_n555), .B2(new_n508), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n557), .B(new_n536), .C1(new_n503), .C2(new_n506), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n515), .A2(KEYINPUT104), .A3(new_n540), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT104), .B1(new_n515), .B2(new_n540), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n554), .B(new_n558), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n536), .A2(KEYINPUT10), .ZN(new_n562));
  OR3_X1    g361(.A1(new_n515), .A2(KEYINPUT106), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT106), .B1(new_n515), .B2(new_n562), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n559), .A2(new_n560), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n569), .A2(new_n558), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n568), .B1(new_n570), .B2(new_n567), .ZN(new_n571));
  XNOR2_X1  g370(.A(G120gat), .B(G148gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(G176gat), .B(G204gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n574), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(KEYINPUT107), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT107), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n571), .A2(new_n579), .A3(new_n574), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n431), .A2(new_n485), .A3(new_n553), .A4(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(new_n362), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n584), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g384(.A1(new_n583), .A2(new_n322), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT42), .B1(new_n586), .B2(new_n456), .ZN(new_n587));
  XOR2_X1   g386(.A(KEYINPUT16), .B(G8gat), .Z(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  MUX2_X1   g388(.A(KEYINPUT42), .B(new_n587), .S(new_n589), .Z(G1325gat));
  OAI21_X1  g389(.A(G15gat), .B1(new_n583), .B2(new_n423), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n421), .A2(G15gat), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n591), .B1(new_n583), .B2(new_n592), .ZN(G1326gat));
  OR3_X1    g392(.A1(new_n583), .A2(KEYINPUT108), .A3(new_n270), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT108), .B1(new_n583), .B2(new_n270), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT43), .B(G22gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(G1327gat));
  INV_X1    g397(.A(new_n552), .ZN(new_n599));
  NOR3_X1   g398(.A1(new_n599), .A2(new_n527), .A3(new_n581), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n431), .A2(new_n485), .A3(new_n600), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n601), .A2(G29gat), .A3(new_n362), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT45), .Z(new_n603));
  NAND3_X1  g402(.A1(new_n431), .A2(KEYINPUT44), .A3(new_n528), .ZN(new_n604));
  INV_X1    g403(.A(new_n485), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n599), .A2(new_n605), .A3(new_n581), .ZN(new_n606));
  INV_X1    g405(.A(new_n413), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n270), .A2(new_n427), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n430), .B1(new_n608), .B2(KEYINPUT35), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT109), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n422), .B1(new_n270), .B2(new_n384), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n609), .A2(new_n610), .B1(new_n611), .B2(new_n364), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT109), .B1(new_n428), .B2(new_n430), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n527), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n604), .B(new_n606), .C1(new_n614), .C2(KEYINPUT44), .ZN(new_n615));
  OAI21_X1  g414(.A(G29gat), .B1(new_n615), .B2(new_n362), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n603), .A2(new_n616), .ZN(G1328gat));
  OAI21_X1  g416(.A(G36gat), .B1(new_n615), .B2(new_n322), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT46), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n376), .A2(new_n442), .ZN(new_n620));
  OR3_X1    g419(.A1(new_n601), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n619), .B1(new_n601), .B2(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT110), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n618), .A2(KEYINPUT110), .A3(new_n623), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(G1329gat));
  NAND2_X1  g427(.A1(new_n422), .A2(G43gat), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n601), .A2(new_n421), .ZN(new_n630));
  OAI22_X1  g429(.A1(new_n615), .A2(new_n629), .B1(G43gat), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g431(.A1(new_n271), .A2(G50gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n601), .A2(new_n270), .ZN(new_n634));
  OAI22_X1  g433(.A1(new_n615), .A2(new_n633), .B1(G50gat), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g435(.A(new_n430), .ZN(new_n637));
  AOI211_X1 g436(.A(new_n363), .B(new_n413), .C1(new_n265), .C2(new_n269), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n637), .B(new_n610), .C1(new_n638), .C2(new_n425), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n613), .A2(new_n424), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT111), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n553), .A2(new_n605), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n582), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n641), .B1(new_n640), .B2(new_n643), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n362), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g448(.A1(new_n640), .A2(new_n643), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT111), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n322), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT112), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n651), .A2(KEYINPUT112), .A3(new_n652), .A4(new_n653), .ZN(new_n657));
  OR2_X1    g456(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n658), .B1(new_n656), .B2(new_n657), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(G1333gat));
  INV_X1    g460(.A(G71gat), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n651), .A2(new_n662), .A3(new_n420), .A4(new_n652), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n644), .A2(new_n645), .A3(new_n423), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n663), .B1(new_n664), .B2(new_n662), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT50), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI211_X1 g466(.A(KEYINPUT50), .B(new_n663), .C1(new_n664), .C2(new_n662), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(G1334gat));
  NAND2_X1  g468(.A1(new_n646), .A2(new_n271), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g470(.A1(new_n599), .A2(new_n485), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n582), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n604), .B(new_n674), .C1(new_n614), .C2(KEYINPUT44), .ZN(new_n675));
  OAI21_X1  g474(.A(G85gat), .B1(new_n675), .B2(new_n362), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT51), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n673), .B1(KEYINPUT113), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n640), .A2(new_n528), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT113), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n680), .A3(KEYINPUT51), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(KEYINPUT51), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n614), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n681), .A2(new_n683), .A3(new_n581), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n362), .A2(G85gat), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n676), .B1(new_n684), .B2(new_n685), .ZN(G1336gat));
  OAI21_X1  g485(.A(G92gat), .B1(new_n675), .B2(new_n322), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n322), .A2(G92gat), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n681), .A2(new_n683), .A3(new_n581), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT52), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT52), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n687), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(G1337gat));
  INV_X1    g493(.A(G99gat), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n675), .A2(new_n695), .A3(new_n423), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n684), .A2(new_n421), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(new_n695), .ZN(G1338gat));
  OAI21_X1  g497(.A(G106gat), .B1(new_n675), .B2(new_n270), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n270), .A2(G106gat), .A3(new_n582), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n681), .A2(new_n683), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT53), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT53), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n699), .A2(new_n704), .A3(new_n701), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(G1339gat));
  NOR2_X1   g505(.A1(new_n642), .A2(new_n581), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n472), .A2(new_n482), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n464), .A2(new_n466), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n470), .A2(new_n465), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI22_X1  g510(.A1(new_n708), .A2(new_n480), .B1(new_n711), .B2(new_n478), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n525), .A2(new_n712), .A3(new_n526), .ZN(new_n713));
  INV_X1    g512(.A(new_n567), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n561), .A2(new_n565), .A3(new_n714), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n568), .A2(KEYINPUT114), .A3(KEYINPUT54), .A4(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n574), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n714), .B1(new_n561), .B2(new_n565), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT54), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n718), .A2(new_n719), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT114), .B1(new_n722), .B2(new_n715), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n575), .B1(new_n724), .B2(KEYINPUT55), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT55), .ZN(new_n726));
  OAI211_X1 g525(.A(KEYINPUT115), .B(new_n726), .C1(new_n721), .C2(new_n723), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n721), .B2(new_n723), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT115), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n725), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT116), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT116), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n725), .A2(new_n730), .A3(new_n733), .A4(new_n727), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n713), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n732), .A2(new_n485), .A3(new_n734), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n712), .A2(new_n581), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT117), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n528), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n737), .A2(KEYINPUT117), .A3(new_n738), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n736), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT118), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n599), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n739), .A2(new_n740), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(new_n527), .A3(new_n742), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n735), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT118), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n707), .B1(new_n745), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n426), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n376), .A2(new_n362), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(G113gat), .B1(new_n754), .B2(new_n485), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT119), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n750), .B2(new_n271), .ZN(new_n757));
  INV_X1    g556(.A(new_n707), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n747), .A2(new_n744), .A3(new_n735), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n552), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n743), .A2(new_n744), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(KEYINPUT119), .A3(new_n270), .ZN(new_n763));
  AOI211_X1 g562(.A(new_n421), .B(new_n753), .C1(new_n757), .C2(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n485), .A2(G113gat), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n755), .B1(new_n764), .B2(new_n765), .ZN(G1340gat));
  AOI21_X1  g565(.A(G120gat), .B1(new_n754), .B2(new_n581), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n581), .A2(G120gat), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n764), .B2(new_n768), .ZN(G1341gat));
  INV_X1    g568(.A(G127gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n770), .A3(new_n599), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n764), .A2(new_n599), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n772), .B2(new_n770), .ZN(G1342gat));
  NOR2_X1   g572(.A1(new_n750), .A2(new_n753), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n751), .A2(G134gat), .A3(new_n527), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n776), .B(KEYINPUT56), .Z(new_n777));
  NOR2_X1   g576(.A1(new_n753), .A2(new_n421), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n750), .A2(new_n756), .A3(new_n271), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT119), .B1(new_n762), .B2(new_n270), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n528), .B(new_n778), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT120), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n781), .A2(new_n782), .A3(G134gat), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n781), .B2(G134gat), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n777), .B1(new_n783), .B2(new_n784), .ZN(G1343gat));
  INV_X1    g584(.A(G141gat), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n422), .A2(new_n753), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n750), .B2(new_n270), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT121), .B1(new_n721), .B2(new_n723), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n485), .B(new_n576), .C1(KEYINPUT55), .C2(new_n791), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n791), .A2(KEYINPUT55), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n738), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n527), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n735), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n552), .ZN(new_n797));
  AOI211_X1 g596(.A(new_n789), .B(new_n270), .C1(new_n797), .C2(new_n758), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n788), .B1(new_n790), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n786), .B1(new_n800), .B2(new_n485), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n422), .A2(new_n270), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n750), .A2(new_n753), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n605), .A2(G141gat), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT58), .B1(new_n801), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT57), .B1(new_n762), .B2(new_n271), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n787), .B1(new_n809), .B2(new_n798), .ZN(new_n810));
  OAI21_X1  g609(.A(G141gat), .B1(new_n810), .B2(new_n605), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n812), .A3(new_n806), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n808), .A2(new_n813), .ZN(G1344gat));
  NOR3_X1   g613(.A1(new_n753), .A2(G148gat), .A3(new_n582), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n762), .A2(new_n802), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G148gat), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n800), .B2(new_n581), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT57), .B1(new_n750), .B2(new_n270), .ZN(new_n820));
  INV_X1    g619(.A(new_n731), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n713), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n599), .B1(new_n795), .B2(new_n822), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n789), .B(new_n271), .C1(new_n823), .C2(new_n707), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n820), .A2(new_n581), .A3(new_n787), .A4(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n817), .B1(new_n825), .B2(G148gat), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n816), .B1(new_n819), .B2(new_n826), .ZN(G1345gat));
  INV_X1    g626(.A(new_n804), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n828), .A2(KEYINPUT122), .A3(new_n552), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(G155gat), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT122), .B1(new_n828), .B2(new_n552), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n552), .A2(new_n209), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n830), .A2(new_n831), .B1(new_n800), .B2(new_n832), .ZN(G1346gat));
  OAI21_X1  g632(.A(G162gat), .B1(new_n810), .B2(new_n527), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n804), .A2(new_n210), .A3(new_n528), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1347gat));
  NOR3_X1   g635(.A1(new_n750), .A2(new_n647), .A3(new_n322), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n426), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT123), .ZN(new_n839));
  INV_X1    g638(.A(G169gat), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n485), .A2(new_n840), .ZN(new_n841));
  OR3_X1    g640(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n839), .B1(new_n838), .B2(new_n841), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n647), .A2(new_n322), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n420), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n845), .B1(new_n757), .B2(new_n763), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n485), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n842), .B(new_n843), .C1(new_n847), .C2(new_n840), .ZN(G1348gat));
  INV_X1    g647(.A(new_n838), .ZN(new_n849));
  AOI21_X1  g648(.A(G176gat), .B1(new_n849), .B2(new_n581), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n846), .A2(G176gat), .A3(new_n581), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT124), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n846), .A2(new_n853), .A3(G176gat), .A4(new_n581), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n850), .B1(new_n852), .B2(new_n854), .ZN(G1349gat));
  AOI21_X1  g654(.A(new_n285), .B1(new_n846), .B2(new_n599), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n837), .A2(new_n272), .A3(new_n426), .A4(new_n599), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT60), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n860));
  AOI211_X1 g659(.A(new_n552), .B(new_n845), .C1(new_n757), .C2(new_n763), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n860), .B(new_n857), .C1(new_n861), .C2(new_n285), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n862), .ZN(G1350gat));
  NAND3_X1  g662(.A1(new_n849), .A2(new_n273), .A3(new_n528), .ZN(new_n864));
  AOI211_X1 g663(.A(KEYINPUT61), .B(new_n273), .C1(new_n846), .C2(new_n528), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT61), .ZN(new_n866));
  INV_X1    g665(.A(new_n845), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n528), .B(new_n867), .C1(new_n779), .C2(new_n780), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n866), .B1(new_n868), .B2(G190gat), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n864), .B1(new_n865), .B2(new_n869), .ZN(G1351gat));
  INV_X1    g669(.A(KEYINPUT126), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n837), .A2(new_n802), .ZN(new_n872));
  XNOR2_X1  g671(.A(KEYINPUT125), .B(G197gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n485), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n871), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  OR3_X1    g674(.A1(new_n872), .A2(new_n871), .A3(new_n874), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n820), .A2(new_n824), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n422), .A2(new_n647), .A3(new_n322), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n877), .A2(new_n485), .A3(new_n878), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n875), .B(new_n876), .C1(new_n879), .C2(new_n873), .ZN(G1352gat));
  NAND3_X1  g679(.A1(new_n877), .A2(new_n581), .A3(new_n878), .ZN(new_n881));
  XNOR2_X1  g680(.A(KEYINPUT127), .B(G204gat), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR4_X1   g682(.A1(new_n803), .A2(new_n322), .A3(new_n582), .A4(new_n882), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n762), .A2(new_n362), .A3(new_n884), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n885), .B(KEYINPUT62), .Z(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(new_n886), .ZN(G1353gat));
  OR3_X1    g686(.A1(new_n872), .A2(G211gat), .A3(new_n552), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n820), .A2(new_n599), .A3(new_n824), .A4(new_n878), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n889), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT63), .B1(new_n889), .B2(G211gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(G1354gat));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n528), .A3(new_n878), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(G218gat), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n527), .A2(G218gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n872), .B2(new_n895), .ZN(G1355gat));
endmodule


