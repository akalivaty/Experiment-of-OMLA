//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT91), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT92), .ZN(new_n206));
  AOI21_X1  g005(.A(G8gat), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n205), .B1(new_n203), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n207), .B(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G43gat), .B(G50gat), .Z(new_n211));
  INV_X1    g010(.A(KEYINPUT15), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT89), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  OR3_X1    g015(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(KEYINPUT90), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(KEYINPUT90), .B2(new_n217), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n211), .A2(new_n212), .ZN(new_n220));
  NAND2_X1  g019(.A1(G29gat), .A2(G36gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(KEYINPUT88), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n214), .A2(new_n219), .A3(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n217), .A2(new_n215), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n220), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n210), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n210), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(KEYINPUT17), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n230), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G229gat), .A2(G233gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(KEYINPUT93), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT94), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT18), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(new_n239), .B2(new_n238), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n235), .A2(new_n237), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n210), .B(new_n229), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n237), .B(KEYINPUT13), .Z(new_n244));
  AOI22_X1  g043(.A1(new_n242), .A2(KEYINPUT18), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G141gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(G197gat), .ZN(new_n248));
  XOR2_X1   g047(.A(KEYINPUT11), .B(G169gat), .Z(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT12), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT95), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n251), .B1(new_n245), .B2(new_n252), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n246), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n246), .A2(new_n253), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  OR2_X1    g056(.A1(G57gat), .A2(G64gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(G57gat), .A2(G64gat), .ZN(new_n259));
  AND2_X1   g058(.A1(G71gat), .A2(G78gat), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n258), .B(new_n259), .C1(new_n260), .C2(KEYINPUT9), .ZN(new_n261));
  NOR2_X1   g060(.A1(G71gat), .A2(G78gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(KEYINPUT96), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n260), .A2(new_n262), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT21), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n210), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT98), .ZN(new_n268));
  NAND2_X1  g067(.A1(G231gat), .A2(G233gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT97), .ZN(new_n270));
  XOR2_X1   g069(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n268), .B(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n265), .A2(KEYINPUT21), .ZN(new_n274));
  XNOR2_X1  g073(.A(G127gat), .B(G155gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G183gat), .B(G211gat), .Z(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n273), .A2(new_n278), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G85gat), .A2(G92gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT7), .ZN(new_n284));
  NOR2_X1   g083(.A1(G85gat), .A2(G92gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(G99gat), .A2(G106gat), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n285), .B1(KEYINPUT8), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G99gat), .B(G106gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n234), .A2(new_n232), .A3(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(G232gat), .A2(G233gat), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n228), .A2(new_n290), .B1(KEYINPUT41), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G190gat), .B(G218gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n293), .A2(KEYINPUT41), .ZN(new_n298));
  XNOR2_X1  g097(.A(G134gat), .B(G162gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n297), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n282), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n265), .A2(new_n290), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n304), .A2(KEYINPUT100), .A3(KEYINPUT10), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT99), .B1(new_n284), .B2(new_n287), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n265), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n291), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n265), .A2(new_n290), .A3(new_n307), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT10), .B1(new_n311), .B2(KEYINPUT100), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G230gat), .ZN(new_n314));
  INV_X1    g113(.A(G233gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n309), .A2(new_n311), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(G230gat), .A3(G233gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G120gat), .B(G148gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(G176gat), .B(G204gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(KEYINPUT101), .B(KEYINPUT102), .Z(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n319), .A2(new_n324), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n303), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n330));
  XNOR2_X1  g129(.A(G15gat), .B(G43gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(G71gat), .B(G99gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  AND3_X1   g132(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT24), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT65), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT65), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n336), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT23), .ZN(new_n346));
  NAND2_X1  g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT23), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n348), .B1(G169gat), .B2(G176gat), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT25), .B1(new_n344), .B2(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n346), .A2(KEYINPUT25), .A3(new_n349), .A4(new_n347), .ZN(new_n352));
  INV_X1    g151(.A(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT66), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT66), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(G183gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n334), .A2(new_n341), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n352), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT67), .B1(new_n351), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n358), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(new_n350), .A3(KEYINPUT25), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT67), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n365));
  NAND3_X1  g164(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n366), .B1(G183gat), .B2(G190gat), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n342), .B1(new_n337), .B2(new_n338), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n365), .B1(new_n369), .B2(new_n343), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n363), .B(new_n364), .C1(new_n370), .C2(KEYINPUT25), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n345), .A2(KEYINPUT26), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT26), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n347), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n372), .B(new_n337), .C1(new_n374), .C2(new_n345), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n357), .A2(KEYINPUT27), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT27), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G183gat), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n354), .A2(new_n356), .A3(new_n376), .A4(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT28), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT66), .B(G190gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT27), .B(G183gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT28), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n375), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT68), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI211_X1 g186(.A(KEYINPUT68), .B(new_n375), .C1(new_n381), .C2(new_n384), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n361), .B(new_n371), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G134gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(G127gat), .ZN(new_n391));
  INV_X1    g190(.A(G127gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G134gat), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT69), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n390), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(G113gat), .B(G120gat), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n395), .B(new_n396), .C1(KEYINPUT1), .C2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G113gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G120gat), .ZN(new_n400));
  INV_X1    g199(.A(G120gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G113gat), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n402), .A3(KEYINPUT70), .ZN(new_n403));
  OR3_X1    g202(.A1(new_n401), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT1), .ZN(new_n405));
  XNOR2_X1  g204(.A(G127gat), .B(G134gat), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n398), .A2(new_n407), .A3(KEYINPUT71), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT71), .B1(new_n398), .B2(new_n407), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n389), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n375), .ZN(new_n414));
  INV_X1    g213(.A(new_n384), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT28), .B1(new_n382), .B2(new_n383), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT68), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n385), .A2(new_n386), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n420), .A2(new_n411), .A3(new_n371), .A4(new_n361), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n413), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G227gat), .A2(G233gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(KEYINPUT64), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n333), .B1(new_n425), .B2(KEYINPUT32), .ZN(new_n426));
  INV_X1    g225(.A(new_n424), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n427), .B1(new_n413), .B2(new_n421), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT72), .B1(new_n428), .B2(KEYINPUT33), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT72), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT33), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n425), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n426), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n413), .A2(new_n427), .A3(new_n421), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n434), .B(KEYINPUT34), .Z(new_n435));
  OAI211_X1 g234(.A(new_n425), .B(KEYINPUT32), .C1(new_n431), .C2(new_n333), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n435), .B1(new_n433), .B2(new_n436), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n330), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n435), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n430), .B1(new_n425), .B2(new_n431), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n428), .A2(KEYINPUT72), .A3(KEYINPUT33), .ZN(new_n442));
  INV_X1    g241(.A(new_n333), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT32), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n443), .B1(new_n428), .B2(new_n444), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n441), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n436), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n440), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n449));
  INV_X1    g248(.A(new_n330), .ZN(new_n450));
  NOR2_X1   g249(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n448), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G226gat), .A2(G233gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n457), .B(KEYINPUT74), .Z(new_n458));
  NAND2_X1  g257(.A1(new_n389), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n458), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n351), .A2(new_n360), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(new_n385), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n460), .B1(new_n462), .B2(KEYINPUT29), .ZN(new_n463));
  XNOR2_X1  g262(.A(G197gat), .B(G204gat), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT22), .ZN(new_n465));
  INV_X1    g264(.A(G211gat), .ZN(new_n466));
  INV_X1    g265(.A(G218gat), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G211gat), .B(G218gat), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(new_n464), .A3(new_n468), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n463), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n458), .A2(KEYINPUT29), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n389), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n474), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n458), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n475), .A2(new_n480), .A3(KEYINPUT75), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT75), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n477), .A2(new_n482), .A3(new_n478), .A4(new_n479), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G8gat), .B(G36gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(G64gat), .B(G92gat), .ZN(new_n486));
  XOR2_X1   g285(.A(new_n485), .B(new_n486), .Z(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n487), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n481), .A2(new_n483), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(KEYINPUT30), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT30), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n484), .A2(new_n492), .A3(new_n487), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G1gat), .B(G29gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT0), .ZN(new_n496));
  XNOR2_X1  g295(.A(G57gat), .B(G85gat), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n496), .B(new_n497), .Z(new_n498));
  INV_X1    g297(.A(G141gat), .ZN(new_n499));
  INV_X1    g298(.A(G148gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT2), .ZN(new_n502));
  NAND2_X1  g301(.A1(G141gat), .A2(G148gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G162gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G155gat), .ZN(new_n506));
  INV_X1    g305(.A(G155gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(G162gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT76), .B(G162gat), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n502), .B1(new_n511), .B2(G155gat), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n501), .A2(new_n506), .A3(new_n508), .A4(new_n503), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT77), .ZN(new_n515));
  INV_X1    g314(.A(new_n513), .ZN(new_n516));
  AND2_X1   g315(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n518));
  OAI21_X1  g317(.A(G155gat), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT2), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT77), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(new_n510), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n515), .A2(KEYINPUT3), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT3), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n525), .B(new_n510), .C1(new_n512), .C2(new_n513), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT78), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n515), .A2(new_n523), .A3(new_n527), .A4(KEYINPUT3), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n398), .A2(new_n407), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n410), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n516), .A2(new_n520), .B1(new_n509), .B2(new_n504), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n533), .A2(KEYINPUT4), .A3(new_n534), .A4(new_n408), .ZN(new_n535));
  NAND2_X1  g334(.A1(G225gat), .A2(G233gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n521), .A2(new_n398), .A3(new_n510), .A4(new_n407), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT4), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n532), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT5), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n515), .A2(new_n523), .A3(new_n531), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n538), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n543), .B1(new_n545), .B2(new_n537), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n538), .A2(new_n539), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n534), .A3(new_n408), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n548), .B1(new_n549), .B2(new_n539), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n532), .A2(new_n543), .A3(new_n536), .A4(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n498), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT6), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT6), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n547), .A2(new_n551), .A3(new_n498), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT79), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n554), .B(new_n555), .C1(new_n552), .C2(new_n556), .ZN(new_n557));
  AOI211_X1 g356(.A(KEYINPUT79), .B(new_n498), .C1(new_n547), .C2(new_n551), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n553), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n494), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G78gat), .B(G106gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(G228gat), .A2(G233gat), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT29), .B1(new_n472), .B2(new_n473), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n563), .A2(KEYINPUT3), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(new_n534), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT29), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n474), .B1(new_n526), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n562), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n526), .A2(new_n566), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n562), .B1(new_n569), .B2(new_n478), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n515), .B(new_n523), .C1(KEYINPUT3), .C2(new_n563), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT81), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT81), .B1(new_n570), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n568), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(G22gat), .ZN(new_n575));
  INV_X1    g374(.A(G22gat), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n576), .B(new_n568), .C1(new_n572), .C2(new_n573), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n578), .B1(new_n575), .B2(new_n577), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n561), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT82), .B(G50gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n570), .A2(new_n571), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT81), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT81), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n576), .B1(new_n588), .B2(new_n568), .ZN(new_n589));
  INV_X1    g388(.A(new_n577), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n583), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n561), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n581), .A2(new_n582), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n582), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n579), .A2(new_n580), .A3(new_n561), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n592), .B1(new_n591), .B2(new_n593), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n560), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT83), .B1(new_n456), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT37), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n487), .B1(new_n484), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n459), .A2(new_n463), .A3(new_n478), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n477), .A2(new_n474), .A3(new_n479), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT37), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT85), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT38), .B1(new_n606), .B2(new_n607), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n603), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n535), .A2(new_n540), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n524), .A2(new_n528), .B1(new_n407), .B2(new_n398), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n611), .B1(new_n612), .B2(new_n530), .ZN(new_n613));
  INV_X1    g412(.A(new_n546), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n551), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT84), .ZN(new_n616));
  INV_X1    g415(.A(new_n498), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT84), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n547), .A2(new_n618), .A3(new_n551), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n555), .A2(new_n554), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n610), .A2(new_n622), .A3(new_n553), .A4(new_n488), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT86), .ZN(new_n624));
  AOI22_X1  g423(.A1(new_n620), .A2(new_n621), .B1(KEYINPUT6), .B2(new_n552), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT86), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n625), .A2(new_n626), .A3(new_n488), .A4(new_n610), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n603), .B1(new_n602), .B2(new_n484), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT38), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT40), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n536), .B1(new_n532), .B2(new_n550), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n617), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT39), .B1(new_n545), .B2(new_n537), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n634), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n498), .B1(new_n615), .B2(KEYINPUT84), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n631), .A2(new_n636), .B1(new_n637), .B2(new_n619), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n636), .A2(new_n631), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n638), .A2(new_n639), .A3(new_n493), .A4(new_n491), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n581), .A2(new_n582), .A3(new_n594), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n582), .B1(new_n581), .B2(new_n594), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n630), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n560), .A2(new_n595), .A3(new_n599), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT83), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(new_n455), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n601), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n448), .A2(new_n449), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(new_n595), .B2(new_n599), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n559), .A3(new_n494), .ZN(new_n652));
  INV_X1    g451(.A(new_n494), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT87), .B(KEYINPUT35), .Z(new_n654));
  NOR3_X1   g453(.A1(new_n653), .A2(new_n625), .A3(new_n654), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n652), .A2(KEYINPUT35), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI211_X1 g456(.A(new_n257), .B(new_n329), .C1(new_n649), .C2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n559), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G1gat), .ZN(G1324gat));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n658), .A2(new_n653), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT16), .B(G8gat), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n665), .A2(KEYINPUT42), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(G8gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(KEYINPUT42), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(G1325gat));
  INV_X1    g468(.A(new_n650), .ZN(new_n670));
  AOI21_X1  g469(.A(G15gat), .B1(new_n658), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT104), .Z(new_n672));
  NOR3_X1   g471(.A1(new_n437), .A2(new_n438), .A3(new_n452), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n450), .B1(new_n448), .B2(new_n449), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT105), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n439), .A2(new_n454), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n679), .A2(G15gat), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n672), .B1(new_n658), .B2(new_n680), .ZN(G1326gat));
  NAND2_X1  g480(.A1(new_n599), .A2(new_n595), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n658), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n439), .A2(new_n454), .A3(new_n676), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n676), .B1(new_n439), .B2(new_n454), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n646), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI22_X1  g489(.A1(new_n623), .A2(KEYINPUT86), .B1(KEYINPUT38), .B2(new_n628), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n643), .B1(new_n691), .B2(new_n627), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT106), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n645), .A2(new_n678), .A3(new_n694), .A4(new_n646), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n656), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n687), .B1(new_n696), .B2(new_n301), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n657), .A2(new_n649), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(KEYINPUT44), .A3(new_n302), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n282), .A2(new_n328), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n700), .A2(new_n257), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G29gat), .B1(new_n703), .B2(new_n559), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n698), .A2(new_n256), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n705), .A2(new_n301), .A3(new_n701), .ZN(new_n706));
  INV_X1    g505(.A(G29gat), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n706), .A2(new_n707), .A3(new_n659), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT45), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n704), .A2(new_n709), .ZN(G1328gat));
  INV_X1    g509(.A(G36gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n706), .A2(new_n711), .A3(new_n653), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT46), .Z(new_n713));
  OAI21_X1  g512(.A(G36gat), .B1(new_n703), .B2(new_n494), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1329gat));
  INV_X1    g514(.A(G43gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n706), .A2(new_n716), .A3(new_n670), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n679), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT108), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G43gat), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n718), .A2(KEYINPUT108), .ZN(new_n721));
  OAI211_X1 g520(.A(KEYINPUT47), .B(new_n717), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n717), .B(KEYINPUT107), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(G43gat), .B2(new_n718), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(KEYINPUT47), .B2(new_n724), .ZN(G1330gat));
  NAND3_X1  g524(.A1(new_n702), .A2(G50gat), .A3(new_n683), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n706), .A2(new_n683), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(G50gat), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g528(.A1(new_n690), .A2(new_n692), .A3(KEYINPUT106), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n600), .B1(new_n675), .B2(new_n677), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n694), .B1(new_n731), .B2(new_n645), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n657), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  AND4_X1   g532(.A1(new_n257), .A2(new_n733), .A3(new_n303), .A4(new_n327), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n659), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n653), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT49), .B(G64gat), .Z(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(G1333gat));
  INV_X1    g539(.A(G71gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n734), .A2(new_n741), .A3(new_n670), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n734), .A2(new_n679), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(new_n741), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n744), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g544(.A1(new_n734), .A2(new_n683), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT109), .B(G78gat), .Z(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1335gat));
  NOR2_X1   g547(.A1(new_n256), .A2(new_n281), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n302), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n733), .A2(KEYINPUT51), .A3(new_n302), .A4(new_n749), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n752), .A2(KEYINPUT110), .A3(new_n753), .ZN(new_n754));
  OR3_X1    g553(.A1(new_n750), .A2(KEYINPUT110), .A3(new_n751), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n328), .A2(G85gat), .A3(new_n559), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT111), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n256), .A2(new_n281), .A3(new_n328), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n697), .A2(new_n699), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760), .B2(new_n559), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(G1336gat));
  NOR3_X1   g561(.A1(new_n328), .A2(G92gat), .A3(new_n494), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n754), .A2(new_n755), .A3(new_n763), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n697), .A2(new_n653), .A3(new_n699), .A4(new_n759), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G92gat), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n767), .A2(KEYINPUT52), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(KEYINPUT52), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n764), .A2(new_n766), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n752), .A2(KEYINPUT113), .A3(new_n753), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n750), .A2(new_n772), .A3(new_n751), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(new_n763), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n765), .A2(KEYINPUT112), .A3(G92gat), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT112), .B1(new_n765), .B2(G92gat), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n771), .A2(KEYINPUT114), .A3(new_n763), .A4(new_n773), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n776), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n781), .A2(new_n782), .A3(KEYINPUT52), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n781), .B2(KEYINPUT52), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n770), .B1(new_n783), .B2(new_n784), .ZN(G1337gat));
  NOR3_X1   g584(.A1(new_n650), .A2(new_n328), .A3(G99gat), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n754), .A2(new_n755), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G99gat), .B1(new_n760), .B2(new_n678), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(G1338gat));
  NOR3_X1   g588(.A1(new_n682), .A2(G106gat), .A3(new_n328), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n754), .A2(new_n755), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  OAI21_X1  g591(.A(G106gat), .B1(new_n760), .B2(new_n682), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n771), .A2(new_n773), .A3(new_n790), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n793), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n796), .A2(KEYINPUT117), .A3(KEYINPUT53), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT117), .B1(new_n796), .B2(KEYINPUT53), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(G1339gat));
  NOR2_X1   g598(.A1(new_n329), .A2(new_n256), .ZN(new_n800));
  OAI211_X1 g599(.A(G230gat), .B(G233gat), .C1(new_n310), .C2(new_n312), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n316), .A2(KEYINPUT54), .A3(new_n801), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n802), .B(new_n324), .C1(KEYINPUT54), .C2(new_n316), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n325), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n256), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n241), .A2(new_n245), .A3(new_n251), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n235), .A2(new_n237), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n243), .A2(new_n244), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n250), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n810), .A2(new_n327), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n301), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n810), .A2(KEYINPUT118), .A3(new_n813), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n808), .A3(new_n302), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT118), .B1(new_n810), .B2(new_n813), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT119), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OR3_X1    g619(.A1(new_n818), .A2(KEYINPUT119), .A3(new_n819), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n816), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n800), .B1(new_n822), .B2(new_n282), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n823), .A2(new_n650), .A3(new_n683), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n653), .A2(new_n559), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n257), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(new_n399), .ZN(G1340gat));
  NOR2_X1   g627(.A1(new_n826), .A2(new_n328), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(new_n401), .ZN(G1341gat));
  NOR2_X1   g629(.A1(new_n826), .A2(new_n282), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(new_n392), .ZN(G1342gat));
  NOR2_X1   g631(.A1(new_n301), .A2(new_n653), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT120), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n824), .A2(new_n390), .A3(new_n659), .A4(new_n834), .ZN(new_n835));
  XOR2_X1   g634(.A(new_n835), .B(KEYINPUT56), .Z(new_n836));
  OAI21_X1  g635(.A(G134gat), .B1(new_n826), .B2(new_n301), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1343gat));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n282), .ZN(new_n839));
  INV_X1    g638(.A(new_n800), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n683), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n678), .A2(new_n825), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n499), .A3(new_n256), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n821), .A2(new_n820), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n808), .A2(KEYINPUT121), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n808), .A2(KEYINPUT121), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n256), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n302), .B1(new_n851), .B2(new_n814), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n282), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n840), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n682), .A2(new_n846), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI211_X1 g655(.A(new_n257), .B(new_n843), .C1(new_n847), .C2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n845), .B1(new_n857), .B2(new_n499), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT58), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n860), .B(new_n845), .C1(new_n857), .C2(new_n499), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(G1344gat));
  NOR2_X1   g661(.A1(new_n500), .A2(KEYINPUT59), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n843), .B1(new_n847), .B2(new_n856), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n863), .B1(new_n865), .B2(new_n328), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n800), .B(KEYINPUT122), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n818), .A2(new_n819), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n282), .B1(new_n852), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n682), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n855), .ZN(new_n871));
  OAI22_X1  g670(.A1(new_n870), .A2(KEYINPUT57), .B1(new_n823), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n843), .A2(new_n328), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(G148gat), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n873), .B1(new_n872), .B2(new_n874), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT59), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n866), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n844), .A2(new_n500), .A3(new_n327), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1345gat));
  OAI21_X1  g680(.A(G155gat), .B1(new_n865), .B2(new_n282), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n844), .A2(new_n507), .A3(new_n281), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1346gat));
  NOR2_X1   g683(.A1(new_n823), .A2(new_n682), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n679), .A2(new_n511), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n885), .A2(new_n659), .A3(new_n834), .A4(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n864), .A2(KEYINPUT124), .A3(new_n302), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n511), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT124), .B1(new_n864), .B2(new_n302), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(G1347gat));
  NOR2_X1   g690(.A1(new_n659), .A2(new_n494), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n824), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(G169gat), .B1(new_n893), .B2(new_n256), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n892), .B(KEYINPUT125), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n824), .A2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(G169gat), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n896), .A2(new_n897), .A3(new_n257), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n894), .A2(new_n898), .ZN(G1348gat));
  INV_X1    g698(.A(G176gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n893), .A2(new_n900), .A3(new_n327), .ZN(new_n901));
  OAI21_X1  g700(.A(G176gat), .B1(new_n896), .B2(new_n328), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1349gat));
  NAND3_X1  g702(.A1(new_n893), .A2(new_n383), .A3(new_n281), .ZN(new_n904));
  OAI21_X1  g703(.A(G183gat), .B1(new_n896), .B2(new_n282), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g706(.A1(new_n893), .A2(new_n382), .A3(new_n302), .ZN(new_n908));
  OAI21_X1  g707(.A(G190gat), .B1(new_n896), .B2(new_n301), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n909), .A2(KEYINPUT61), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n909), .A2(KEYINPUT61), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1351gat));
  NAND2_X1  g711(.A1(new_n678), .A2(new_n892), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n842), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(G197gat), .B1(new_n914), .B2(new_n256), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n872), .A2(KEYINPUT126), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n895), .A2(new_n678), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n872), .A2(KEYINPUT126), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n256), .A2(G197gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n915), .B1(new_n920), .B2(new_n921), .ZN(G1352gat));
  OAI21_X1  g721(.A(G204gat), .B1(new_n919), .B2(new_n328), .ZN(new_n923));
  NOR4_X1   g722(.A1(new_n842), .A2(G204gat), .A3(new_n328), .A4(new_n913), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT62), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1353gat));
  NAND3_X1  g725(.A1(new_n914), .A2(new_n466), .A3(new_n281), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n872), .A2(new_n281), .A3(new_n917), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n928), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT63), .B1(new_n928), .B2(G211gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(G1354gat));
  AOI21_X1  g730(.A(G218gat), .B1(new_n914), .B2(new_n302), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n301), .A2(new_n467), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n920), .B2(new_n933), .ZN(G1355gat));
endmodule


