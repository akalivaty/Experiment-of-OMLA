//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(KEYINPUT81), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  INV_X1    g007(.A(G211gat), .ZN(new_n209));
  INV_X1    g008(.A(G218gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n208), .B1(KEYINPUT22), .B2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(G211gat), .B(G218gat), .Z(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n212), .B(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT74), .ZN(new_n217));
  XOR2_X1   g016(.A(G141gat), .B(G148gat), .Z(new_n218));
  INV_X1    g017(.A(G155gat), .ZN(new_n219));
  INV_X1    g018(.A(G162gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n218), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G141gat), .B(G148gat), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n222), .B(new_n221), .C1(new_n226), .C2(KEYINPUT2), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n217), .B1(new_n228), .B2(KEYINPUT3), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n225), .A2(new_n227), .A3(KEYINPUT74), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT29), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n216), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n234), .B1(G228gat), .B2(G233gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n215), .A2(KEYINPUT29), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n230), .B1(new_n236), .B2(KEYINPUT80), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n216), .A2(KEYINPUT80), .A3(new_n233), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n228), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n225), .A2(new_n227), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n216), .A2(new_n233), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(new_n230), .ZN(new_n243));
  OAI211_X1 g042(.A(G228gat), .B(G233gat), .C1(new_n243), .C2(new_n234), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n240), .A2(G22gat), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(G22gat), .B1(new_n240), .B2(new_n244), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n207), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n240), .A2(new_n244), .ZN(new_n248));
  INV_X1    g047(.A(G22gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n204), .B(KEYINPUT81), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n240), .A2(G22gat), .A3(new_n244), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G226gat), .A2(G233gat), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n257), .B(KEYINPUT72), .Z(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G183gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT66), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT66), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G183gat), .ZN(new_n263));
  INV_X1    g062(.A(G190gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT24), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n266), .A2(KEYINPUT65), .A3(new_n267), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n265), .A2(new_n270), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n274));
  INV_X1    g073(.A(G169gat), .ZN(new_n275));
  INV_X1    g074(.A(G176gat), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT64), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT64), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(G169gat), .A3(G176gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT23), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n277), .A2(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n273), .A2(new_n274), .A3(new_n284), .A4(KEYINPUT25), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n273), .A2(KEYINPUT25), .A3(new_n284), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT25), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n268), .B(new_n271), .C1(G183gat), .C2(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n286), .A2(KEYINPUT67), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT27), .B(G183gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n292));
  OR2_X1    g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n292), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n264), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT28), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT27), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G183gat), .ZN(new_n299));
  AOI211_X1 g098(.A(KEYINPUT28), .B(G190gat), .C1(new_n299), .C2(KEYINPUT68), .ZN(new_n300));
  OR2_X1    g099(.A1(new_n299), .A2(KEYINPUT68), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n261), .A2(new_n263), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n300), .B(new_n301), .C1(new_n298), .C2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n280), .B(KEYINPUT26), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n277), .A2(new_n279), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n304), .A2(new_n305), .B1(G183gat), .B2(G190gat), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n285), .A2(new_n290), .B1(new_n297), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n259), .B1(new_n308), .B2(KEYINPUT29), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n289), .A2(new_n287), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(new_n285), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(G190gat), .B1(new_n293), .B2(new_n294), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n303), .B(new_n306), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT73), .B1(new_n316), .B2(new_n258), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n318));
  AOI211_X1 g117(.A(new_n318), .B(new_n259), .C1(new_n312), .C2(new_n315), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n309), .B(new_n216), .C1(new_n317), .C2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n258), .B1(new_n316), .B2(new_n233), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n308), .A2(new_n259), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n215), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G8gat), .B(G36gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(G64gat), .B(G92gat), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n325), .B(new_n326), .Z(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n320), .A2(new_n323), .A3(new_n327), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(KEYINPUT30), .A3(new_n330), .ZN(new_n331));
  OR3_X1    g130(.A1(new_n324), .A2(KEYINPUT30), .A3(new_n328), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT39), .ZN(new_n335));
  XOR2_X1   g134(.A(G127gat), .B(G134gat), .Z(new_n336));
  XNOR2_X1  g135(.A(G113gat), .B(G120gat), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n336), .B1(KEYINPUT1), .B2(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(G113gat), .B(G120gat), .Z(new_n339));
  INV_X1    g138(.A(KEYINPUT1), .ZN(new_n340));
  XNOR2_X1  g139(.A(G127gat), .B(G134gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n228), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n225), .A2(new_n338), .A3(new_n342), .A4(new_n227), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT75), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n335), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n343), .A2(new_n241), .A3(KEYINPUT4), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n346), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n343), .B1(KEYINPUT3), .B2(new_n228), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n355), .B1(new_n232), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n351), .B1(new_n357), .B2(new_n350), .ZN(new_n358));
  XNOR2_X1  g157(.A(G1gat), .B(G29gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT0), .ZN(new_n360));
  XNOR2_X1  g159(.A(G57gat), .B(G85gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  NAND2_X1  g161(.A1(new_n232), .A2(new_n356), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n346), .B(KEYINPUT4), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n365), .A2(new_n335), .A3(new_n349), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n358), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT40), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n362), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT77), .B(KEYINPUT5), .ZN(new_n371));
  OR3_X1    g170(.A1(new_n347), .A2(new_n350), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n371), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT76), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n374), .B1(new_n357), .B2(new_n350), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n363), .A2(new_n364), .A3(new_n350), .A4(new_n374), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n370), .B(new_n372), .C1(new_n375), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n367), .A2(new_n368), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n369), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n256), .B1(new_n334), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT6), .ZN(new_n382));
  OR2_X1    g181(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n363), .A2(new_n364), .A3(new_n350), .ZN(new_n384));
  INV_X1    g183(.A(new_n374), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n376), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n370), .B1(new_n387), .B2(new_n372), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n378), .A2(new_n382), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n383), .B(new_n330), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n324), .A2(KEYINPUT37), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n328), .B1(new_n324), .B2(KEYINPUT37), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT38), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n317), .A2(new_n319), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n215), .B1(new_n395), .B2(new_n321), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n321), .A2(new_n322), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(new_n216), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n398), .B1(new_n397), .B2(new_n216), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT37), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n393), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT38), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n391), .A2(new_n394), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT36), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT32), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n312), .A2(new_n343), .A3(new_n315), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT70), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n312), .A2(KEYINPUT70), .A3(new_n343), .A4(new_n315), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n316), .A2(new_n344), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(G227gat), .A2(G233gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n408), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT33), .B1(new_n414), .B2(new_n416), .ZN(new_n418));
  XOR2_X1   g217(.A(G15gat), .B(G43gat), .Z(new_n419));
  XNOR2_X1  g218(.A(G71gat), .B(G99gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n417), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n411), .A2(new_n413), .A3(new_n415), .A4(new_n412), .ZN(new_n424));
  XOR2_X1   g223(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(KEYINPUT71), .A2(KEYINPUT34), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n426), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AOI221_X4 g228(.A(new_n408), .B1(KEYINPUT33), .B2(new_n421), .C1(new_n414), .C2(new_n416), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n423), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n418), .A2(new_n422), .ZN(new_n432));
  INV_X1    g231(.A(new_n417), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n430), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n428), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n407), .B1(new_n431), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n429), .B1(new_n423), .B2(new_n430), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n434), .A2(new_n435), .A3(new_n428), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT36), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n381), .A2(new_n406), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT78), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n442), .B1(new_n389), .B2(new_n388), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n387), .A2(new_n372), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n362), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n445), .A2(KEYINPUT78), .A3(new_n382), .A4(new_n378), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(new_n446), .A3(new_n383), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n447), .A2(KEYINPUT79), .A3(new_n333), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT79), .B1(new_n447), .B2(new_n333), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n256), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n441), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT35), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n448), .A2(new_n449), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n439), .A3(new_n255), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT83), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n439), .A2(new_n438), .A3(new_n255), .A4(KEYINPUT83), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n452), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n383), .B1(new_n388), .B2(new_n389), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n333), .A2(new_n452), .A3(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(new_n454), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n451), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G15gat), .B(G22gat), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT16), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n464), .B1(new_n465), .B2(G1gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT88), .ZN(new_n467));
  INV_X1    g266(.A(new_n464), .ZN(new_n468));
  INV_X1    g267(.A(G1gat), .ZN(new_n469));
  AOI21_X1  g268(.A(G8gat), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT88), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n464), .B(new_n471), .C1(new_n465), .C2(G1gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n467), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT89), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT89), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n467), .A2(new_n470), .A3(new_n475), .A4(new_n472), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n466), .B1(G1gat), .B2(new_n464), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G8gat), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT91), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n477), .A2(KEYINPUT91), .A3(new_n479), .ZN(new_n482));
  XNOR2_X1  g281(.A(G43gat), .B(G50gat), .ZN(new_n483));
  INV_X1    g282(.A(G29gat), .ZN(new_n484));
  INV_X1    g283(.A(G36gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT14), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT14), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(G29gat), .B2(G36gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n484), .A2(new_n485), .ZN(new_n490));
  OAI211_X1 g289(.A(KEYINPUT15), .B(new_n483), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n489), .B(KEYINPUT87), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n490), .B1(new_n483), .B2(KEYINPUT15), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(KEYINPUT15), .B2(new_n483), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n491), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n481), .A2(new_n482), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n477), .A2(new_n479), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT90), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n477), .A2(KEYINPUT90), .A3(new_n479), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n495), .B(KEYINPUT17), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G229gat), .A2(G233gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n496), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT18), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n495), .ZN(new_n507));
  INV_X1    g306(.A(new_n482), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(new_n480), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n496), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n503), .B(KEYINPUT13), .Z(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n496), .A2(new_n502), .A3(KEYINPUT18), .A4(new_n503), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n506), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G169gat), .B(G197gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(G113gat), .B(G141gat), .Z(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT85), .B(KEYINPUT86), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n521), .B(KEYINPUT12), .Z(new_n522));
  NAND2_X1  g321(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n522), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n524), .A2(new_n513), .A3(new_n512), .A4(new_n506), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n463), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(G57gat), .A2(G64gat), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n530));
  NAND2_X1  g329(.A1(G57gat), .A2(G64gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(G57gat), .A2(G64gat), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT93), .B1(new_n533), .B2(new_n528), .ZN(new_n534));
  OR2_X1    g333(.A1(G71gat), .A2(G78gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(G71gat), .A2(G78gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n532), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT92), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT94), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n533), .A2(new_n528), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n542), .A2(new_n530), .B1(new_n536), .B2(new_n535), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT9), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n536), .A2(KEYINPUT92), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT92), .B1(new_n536), .B2(new_n545), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n543), .A2(new_n544), .A3(new_n548), .A4(new_n534), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n541), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n537), .B1(new_n548), .B2(new_n542), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT95), .B(KEYINPUT21), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g354(.A1(G231gat), .A2(G233gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G127gat), .B(G155gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT20), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n557), .B(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G183gat), .B(G211gat), .Z(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n560), .A2(new_n562), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT97), .B1(new_n550), .B2(new_n552), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n566));
  AOI211_X1 g365(.A(new_n566), .B(new_n551), .C1(new_n541), .C2(new_n549), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n481), .A2(new_n482), .B1(new_n568), .B2(KEYINPUT21), .ZN(new_n569));
  XOR2_X1   g368(.A(KEYINPUT96), .B(KEYINPUT19), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  OR3_X1    g370(.A1(new_n563), .A2(new_n564), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n571), .B1(new_n563), .B2(new_n564), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT8), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n576), .B1(G99gat), .B2(G106gat), .ZN(new_n577));
  AND2_X1   g376(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(G85gat), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G99gat), .B(G106gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT7), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT7), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(G85gat), .A3(G92gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n582), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(new_n581), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(G99gat), .ZN(new_n593));
  INV_X1    g392(.A(G106gat), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT8), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(new_n588), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n583), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n589), .A2(new_n598), .A3(KEYINPUT99), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n583), .B1(new_n582), .B2(new_n588), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT99), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n501), .A2(new_n604), .B1(KEYINPUT41), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n495), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G190gat), .B(G218gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(KEYINPUT100), .Z(new_n610));
  AND2_X1   g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n608), .A2(new_n610), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n605), .A2(KEYINPUT41), .ZN(new_n613));
  XNOR2_X1  g412(.A(G134gat), .B(G162gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OR3_X1    g415(.A1(new_n611), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n616), .B1(new_n611), .B2(new_n612), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n575), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G120gat), .B(G148gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n553), .A2(new_n602), .A3(new_n599), .ZN(new_n626));
  AND4_X1   g425(.A1(new_n583), .A2(new_n592), .A3(new_n588), .A4(new_n595), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n600), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n550), .A2(new_n628), .A3(new_n552), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT103), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n603), .A2(KEYINPUT10), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n635), .A2(new_n565), .A3(new_n567), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n551), .B1(new_n541), .B2(new_n549), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n629), .B(new_n637), .C1(new_n638), .C2(new_n603), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n626), .A2(KEYINPUT101), .A3(new_n637), .A4(new_n629), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n636), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n643), .A2(new_n632), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n625), .B1(new_n634), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT104), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n647), .B(new_n625), .C1(new_n634), .C2(new_n644), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n641), .A2(new_n642), .ZN(new_n650));
  INV_X1    g449(.A(new_n636), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n643), .A2(KEYINPUT102), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(new_n655), .A3(new_n631), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n634), .A2(new_n625), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n649), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n621), .A2(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n527), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n447), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n334), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n665), .A2(G8gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT105), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G8gat), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT42), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n669), .A2(KEYINPUT42), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(G1325gat));
  INV_X1    g471(.A(new_n661), .ZN(new_n673));
  INV_X1    g472(.A(new_n440), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT36), .B1(new_n438), .B2(new_n439), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT106), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(new_n674), .B2(new_n675), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G15gat), .B1(new_n673), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n431), .A2(new_n436), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n683), .A2(G15gat), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n681), .B1(new_n673), .B2(new_n684), .ZN(G1326gat));
  NAND2_X1  g484(.A1(new_n661), .A2(new_n256), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  INV_X1    g487(.A(new_n659), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n574), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n523), .A2(new_n525), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n463), .A2(new_n619), .ZN(new_n694));
  AND2_X1   g493(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n695));
  NOR2_X1   g494(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n695), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n463), .A2(new_n619), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n693), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G29gat), .B1(new_n703), .B2(new_n447), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n690), .A2(new_n620), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n527), .A2(new_n484), .A3(new_n662), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT45), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n707), .ZN(G1328gat));
  NAND2_X1  g507(.A1(new_n527), .A2(new_n705), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(G36gat), .A3(new_n333), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT46), .ZN(new_n711));
  OAI21_X1  g510(.A(G36gat), .B1(new_n703), .B2(new_n333), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(G1329gat));
  NOR3_X1   g512(.A1(new_n709), .A2(G43gat), .A3(new_n683), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n702), .A2(new_n679), .A3(new_n677), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n715), .B2(G43gat), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(G43gat), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n719), .B1(new_n702), .B2(new_n676), .ZN(new_n720));
  OAI22_X1  g519(.A1(new_n716), .A2(KEYINPUT47), .B1(new_n718), .B2(new_n720), .ZN(G1330gat));
  NOR3_X1   g520(.A1(new_n709), .A2(G50gat), .A3(new_n255), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT48), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n463), .A2(new_n619), .A3(new_n700), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n697), .B1(new_n463), .B2(new_n619), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n256), .B(new_n692), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G50gat), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n727), .A2(new_n728), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n724), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n727), .A2(G50gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n723), .B1(new_n733), .B2(new_n722), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1331gat));
  NOR2_X1   g534(.A1(new_n621), .A2(new_n526), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n463), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n659), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n447), .B(KEYINPUT109), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g542(.A1(new_n689), .A2(new_n333), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n737), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT49), .B(G64gat), .Z(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT110), .ZN(G1333gat));
  OAI21_X1  g548(.A(G71gat), .B1(new_n738), .B2(new_n680), .ZN(new_n750));
  INV_X1    g549(.A(G71gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n682), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n738), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1334gat));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n256), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g556(.A1(new_n575), .A2(new_n526), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n659), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n725), .B2(new_n726), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT111), .B1(new_n761), .B2(new_n447), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G85gat), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n761), .A2(KEYINPUT111), .A3(new_n447), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n463), .A2(new_n619), .A3(new_n758), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n463), .A2(KEYINPUT51), .A3(new_n619), .A4(new_n758), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n659), .A2(new_n581), .A3(new_n662), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT112), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n763), .A2(new_n764), .B1(new_n770), .B2(new_n772), .ZN(G1336gat));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n774));
  INV_X1    g573(.A(G92gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n744), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n770), .B2(new_n776), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n334), .B(new_n760), .C1(new_n725), .C2(new_n726), .ZN(new_n778));
  INV_X1    g577(.A(new_n580), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT52), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n776), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n769), .A2(KEYINPUT114), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n777), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n759), .B1(new_n699), .B2(new_n701), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n580), .B1(new_n784), .B2(new_n334), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n769), .B2(new_n781), .ZN(new_n787));
  AOI211_X1 g586(.A(KEYINPUT113), .B(new_n776), .C1(new_n767), .C2(new_n768), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n783), .B1(new_n789), .B2(new_n790), .ZN(G1337gat));
  OAI21_X1  g590(.A(G99gat), .B1(new_n761), .B2(new_n680), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n659), .A2(new_n682), .A3(new_n593), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n770), .B2(new_n793), .ZN(G1338gat));
  OAI211_X1 g593(.A(new_n256), .B(new_n760), .C1(new_n725), .C2(new_n726), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G106gat), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n689), .A2(G106gat), .A3(new_n255), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT115), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n770), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT53), .B1(new_n769), .B2(new_n797), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n801), .A2(new_n802), .A3(new_n796), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n801), .B2(new_n796), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n800), .B1(new_n803), .B2(new_n804), .ZN(G1339gat));
  NOR3_X1   g604(.A1(new_n621), .A2(new_n526), .A3(new_n659), .ZN(new_n806));
  INV_X1    g605(.A(new_n658), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n624), .B1(new_n644), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n808), .B1(new_n643), .B2(new_n632), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n631), .B1(new_n643), .B2(KEYINPUT102), .ZN(new_n812));
  AOI211_X1 g611(.A(new_n653), .B(new_n636), .C1(new_n641), .C2(new_n642), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g615(.A(KEYINPUT117), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n810), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n807), .B1(new_n818), .B2(KEYINPUT55), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT117), .B1(new_n656), .B2(new_n811), .ZN(new_n820));
  INV_X1    g619(.A(new_n817), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n809), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n510), .A2(new_n511), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n503), .B1(new_n496), .B2(new_n502), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n521), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n525), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n819), .A2(new_n824), .A3(new_n619), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n828), .B1(new_n649), .B2(new_n658), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n691), .B1(new_n822), .B2(new_n823), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(new_n819), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n830), .B1(new_n833), .B2(new_n619), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n806), .B1(new_n834), .B2(new_n574), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n256), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n662), .A2(new_n333), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n683), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(G113gat), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n839), .A2(new_n840), .A3(new_n691), .ZN(new_n841));
  INV_X1    g640(.A(new_n458), .ZN(new_n842));
  NOR4_X1   g641(.A1(new_n835), .A2(new_n334), .A3(new_n842), .A4(new_n740), .ZN(new_n843));
  AOI21_X1  g642(.A(G113gat), .B1(new_n843), .B2(new_n526), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n841), .A2(new_n844), .ZN(G1340gat));
  NAND3_X1  g644(.A1(new_n836), .A2(new_n659), .A3(new_n838), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n846), .A2(KEYINPUT118), .A3(G120gat), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT118), .B1(new_n846), .B2(G120gat), .ZN(new_n848));
  INV_X1    g647(.A(new_n843), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n689), .A2(G120gat), .ZN(new_n850));
  OAI22_X1  g649(.A1(new_n847), .A2(new_n848), .B1(new_n849), .B2(new_n850), .ZN(G1341gat));
  OAI21_X1  g650(.A(G127gat), .B1(new_n839), .B2(new_n574), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n574), .A2(G127gat), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n849), .B2(new_n853), .ZN(G1342gat));
  INV_X1    g653(.A(G134gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n843), .A2(new_n855), .A3(new_n619), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857));
  OR3_X1    g656(.A1(new_n856), .A2(new_n857), .A3(KEYINPUT56), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n856), .B2(KEYINPUT56), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n836), .A2(new_n619), .A3(new_n838), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT56), .B1(new_n860), .B2(G134gat), .ZN(new_n861));
  INV_X1    g660(.A(new_n856), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n858), .B(new_n859), .C1(new_n861), .C2(new_n862), .ZN(G1343gat));
  NOR2_X1   g662(.A1(new_n676), .A2(new_n837), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n255), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n868), .B1(new_n833), .B2(new_n619), .ZN(new_n869));
  INV_X1    g668(.A(new_n831), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n658), .B1(new_n822), .B2(new_n823), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n526), .B1(new_n818), .B2(KEYINPUT55), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(KEYINPUT120), .A3(new_n620), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n869), .A2(new_n830), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n574), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n660), .A2(new_n691), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n867), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n828), .B(new_n620), .C1(new_n823), .C2(new_n822), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n873), .A2(new_n620), .B1(new_n879), .B2(new_n819), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n877), .B1(new_n880), .B2(new_n575), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(new_n881), .B2(new_n256), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n526), .B(new_n864), .C1(new_n878), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(G141gat), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n255), .B1(new_n677), .B2(new_n679), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n333), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n691), .A2(G141gat), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT121), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n881), .A2(new_n741), .A3(new_n886), .A4(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n884), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n835), .A2(new_n740), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n893), .A2(KEYINPUT122), .A3(new_n886), .A4(new_n888), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(new_n883), .B2(G141gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n892), .B1(new_n890), .B2(new_n898), .ZN(G1344gat));
  NOR2_X1   g698(.A1(new_n689), .A2(G148gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n893), .A2(new_n886), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT123), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G148gat), .ZN(new_n904));
  INV_X1    g703(.A(new_n864), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n876), .A2(new_n877), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n866), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n865), .B1(new_n835), .B2(new_n255), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n904), .B1(new_n909), .B2(new_n659), .ZN(new_n910));
  XOR2_X1   g709(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n911));
  NAND2_X1  g710(.A1(new_n881), .A2(new_n866), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n659), .A3(new_n864), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n911), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n902), .B1(new_n910), .B2(new_n915), .ZN(G1345gat));
  OAI21_X1  g715(.A(new_n864), .B1(new_n878), .B2(new_n882), .ZN(new_n917));
  OAI21_X1  g716(.A(G155gat), .B1(new_n917), .B2(new_n574), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n893), .A2(new_n886), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n575), .A2(new_n219), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(G1346gat));
  OAI21_X1  g720(.A(G162gat), .B1(new_n917), .B2(new_n620), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n619), .A2(new_n220), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n919), .B2(new_n923), .ZN(G1347gat));
  NOR3_X1   g723(.A1(new_n741), .A2(new_n333), .A3(new_n683), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n836), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n926), .A2(new_n275), .A3(new_n691), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n835), .A2(new_n662), .A3(new_n842), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n334), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n526), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n927), .B1(new_n931), .B2(new_n275), .ZN(G1348gat));
  OAI21_X1  g731(.A(G176gat), .B1(new_n926), .B2(new_n689), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n928), .A2(new_n276), .A3(new_n744), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1349gat));
  OAI21_X1  g734(.A(new_n302), .B1(new_n926), .B2(new_n574), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n575), .A2(new_n295), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n929), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT60), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n936), .B(new_n940), .C1(new_n929), .C2(new_n937), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1350gat));
  NAND3_X1  g741(.A1(new_n930), .A2(new_n264), .A3(new_n619), .ZN(new_n943));
  OAI21_X1  g742(.A(G190gat), .B1(new_n926), .B2(new_n620), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(G1351gat));
  XNOR2_X1  g746(.A(KEYINPUT126), .B(G197gat), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n691), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n881), .A2(new_n447), .A3(new_n334), .A4(new_n885), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n951), .A2(new_n952), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n680), .A2(new_n334), .A3(new_n740), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n835), .A2(new_n867), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n959), .B(new_n526), .C1(new_n882), .C2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n949), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n956), .A2(new_n957), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n958), .B1(new_n908), .B2(new_n912), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n948), .B1(new_n964), .B2(new_n526), .ZN(new_n965));
  INV_X1    g764(.A(new_n950), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n835), .A2(new_n662), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n967), .A2(KEYINPUT125), .A3(new_n334), .A4(new_n885), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n966), .B1(new_n968), .B2(new_n953), .ZN(new_n969));
  OAI21_X1  g768(.A(KEYINPUT127), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n963), .A2(new_n970), .ZN(G1352gat));
  INV_X1    g770(.A(G204gat), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n967), .A2(new_n972), .A3(new_n744), .A4(new_n885), .ZN(new_n973));
  XOR2_X1   g772(.A(new_n973), .B(KEYINPUT62), .Z(new_n974));
  INV_X1    g773(.A(new_n964), .ZN(new_n975));
  OAI21_X1  g774(.A(G204gat), .B1(new_n975), .B2(new_n689), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n976), .ZN(G1353gat));
  OAI211_X1 g776(.A(new_n209), .B(new_n575), .C1(new_n954), .C2(new_n955), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n964), .A2(new_n575), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n979), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT63), .B1(new_n979), .B2(G211gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(G1354gat));
  OAI21_X1  g781(.A(G218gat), .B1(new_n975), .B2(new_n620), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n210), .B(new_n619), .C1(new_n954), .C2(new_n955), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1355gat));
endmodule


