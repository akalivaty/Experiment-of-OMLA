//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT71), .B(G125), .Z(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  AND3_X1   g003(.A1(new_n189), .A2(KEYINPUT1), .A3(G146), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n190), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n192), .A3(new_n193), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n188), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G224), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G953), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n205));
  OAI211_X1 g019(.A(KEYINPUT0), .B(G128), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  OR2_X1    g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n194), .A2(KEYINPUT64), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n209), .A3(new_n188), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n200), .A2(new_n203), .A3(new_n210), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n206), .A2(new_n209), .A3(new_n188), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n202), .B1(new_n212), .B2(new_n199), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n202), .A2(KEYINPUT7), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G110), .B(G122), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n217), .B(KEYINPUT8), .ZN(new_n218));
  INV_X1    g032(.A(G119), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G116), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(KEYINPUT5), .ZN(new_n221));
  INV_X1    g035(.A(G113), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G116), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G116), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n227), .A3(G119), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n220), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT5), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n223), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT2), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G113), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n228), .A2(new_n220), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G104), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT3), .B1(new_n237), .B2(G107), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n239));
  INV_X1    g053(.A(G107), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(G104), .ZN(new_n241));
  INV_X1    g055(.A(G101), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(G107), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n238), .A2(new_n241), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n237), .A2(G107), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n240), .A2(G104), .ZN(new_n246));
  OAI21_X1  g060(.A(G101), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n231), .A2(new_n236), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n231), .B2(new_n236), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n218), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n200), .A2(new_n210), .A3(new_n214), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n216), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n238), .A2(new_n241), .A3(new_n243), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(G101), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n228), .A2(new_n220), .A3(new_n235), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n235), .B1(new_n228), .B2(new_n220), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(G101), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n261), .A2(KEYINPUT4), .A3(new_n244), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT81), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n231), .A2(new_n236), .A3(new_n248), .ZN(new_n264));
  INV_X1    g078(.A(new_n235), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n229), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n236), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT81), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n261), .A2(KEYINPUT4), .A3(new_n244), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n267), .A2(new_n268), .A3(new_n269), .A4(new_n257), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n263), .A2(new_n217), .A3(new_n264), .A4(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT82), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n271), .A2(new_n272), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n254), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n187), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n270), .A2(new_n264), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n278), .A2(KEYINPUT82), .A3(new_n217), .A4(new_n263), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n271), .A2(new_n272), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n253), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n281), .A2(KEYINPUT84), .A3(G902), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(G210), .B1(G237), .B2(G902), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(KEYINPUT85), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT83), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n263), .A2(new_n264), .A3(new_n270), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT6), .ZN(new_n289));
  INV_X1    g103(.A(new_n217), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n279), .A2(new_n280), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n289), .B1(new_n288), .B2(new_n290), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n211), .A2(new_n213), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n287), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n295), .A2(new_n287), .A3(new_n296), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n283), .B(new_n286), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n275), .A2(new_n187), .A3(new_n276), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT84), .B1(new_n281), .B2(G902), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n295), .A2(new_n296), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT83), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n295), .A2(new_n287), .A3(new_n296), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n302), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n285), .B(KEYINPUT86), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n299), .B(KEYINPUT87), .C1(new_n306), .C2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT87), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n298), .A2(new_n297), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n310), .B(new_n307), .C1(new_n311), .C2(new_n302), .ZN(new_n312));
  INV_X1    g126(.A(G953), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n313), .A2(G952), .ZN(new_n314));
  INV_X1    g128(.A(G234), .ZN(new_n315));
  INV_X1    g129(.A(G237), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XOR2_X1   g131(.A(new_n317), .B(KEYINPUT98), .Z(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT67), .B(G953), .ZN(new_n319));
  AOI211_X1 g133(.A(new_n276), .B(new_n319), .C1(G234), .C2(G237), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT21), .B(G898), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G214), .B1(G237), .B2(G902), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n309), .A2(new_n312), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n206), .A2(new_n209), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT11), .ZN(new_n330));
  INV_X1    g144(.A(G134), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n330), .B1(new_n331), .B2(G137), .ZN(new_n332));
  INV_X1    g146(.A(G137), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(KEYINPUT11), .A3(G134), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(G137), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G131), .ZN(new_n337));
  INV_X1    g151(.A(G131), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n332), .A2(new_n334), .A3(new_n338), .A4(new_n335), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n329), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n335), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n331), .A2(G137), .ZN(new_n343));
  OAI21_X1  g157(.A(G131), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n345));
  OAI22_X1  g159(.A1(new_n204), .A2(G128), .B1(new_n345), .B2(new_n193), .ZN(new_n346));
  INV_X1    g160(.A(new_n198), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n339), .B(new_n344), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n341), .A2(KEYINPUT30), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n348), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n337), .A2(new_n339), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n206), .A2(new_n209), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT65), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT65), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n329), .A2(new_n354), .A3(new_n340), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n350), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n349), .B(new_n267), .C1(new_n356), .C2(KEYINPUT30), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n258), .A2(new_n259), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n358), .B(new_n348), .C1(new_n351), .C2(new_n352), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n319), .A2(G210), .A3(new_n316), .ZN(new_n360));
  XOR2_X1   g174(.A(KEYINPUT26), .B(G101), .Z(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n357), .A2(new_n359), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT31), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT31), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n357), .A2(new_n367), .A3(new_n359), .A4(new_n364), .ZN(new_n368));
  INV_X1    g182(.A(new_n359), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT28), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT28), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n359), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n370), .B(new_n372), .C1(new_n358), .C2(new_n356), .ZN(new_n373));
  INV_X1    g187(.A(new_n364), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n366), .A2(new_n368), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(G472), .A2(G902), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT32), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT32), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n376), .A2(new_n380), .A3(new_n377), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT70), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n359), .A2(new_n382), .A3(new_n371), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n348), .B1(new_n351), .B2(new_n352), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n267), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n371), .B1(new_n385), .B2(new_n359), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n372), .A2(KEYINPUT70), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n383), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n374), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(G902), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT69), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n373), .B2(new_n374), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n356), .A2(new_n358), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n359), .B(KEYINPUT28), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n394), .A2(KEYINPUT69), .A3(new_n364), .A4(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n389), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n364), .B1(new_n357), .B2(new_n359), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n391), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n379), .A2(new_n381), .B1(G472), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G217), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(G234), .B2(new_n276), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n319), .A2(G221), .A3(G234), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT22), .B(G137), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(G125), .A2(G140), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT71), .B(G125), .ZN(new_n410));
  INV_X1    g224(.A(G140), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(KEYINPUT16), .A2(G140), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n412), .A2(KEYINPUT16), .B1(new_n188), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(new_n191), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT23), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n219), .B2(G128), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n417), .B(new_n418), .C1(G119), .C2(new_n195), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G110), .ZN(new_n420));
  XOR2_X1   g234(.A(G119), .B(G128), .Z(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT24), .B(G110), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n415), .A2(new_n423), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n419), .A2(G110), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n422), .ZN(new_n426));
  AND2_X1   g240(.A1(G125), .A2(G140), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n191), .B1(new_n427), .B2(new_n408), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT72), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(KEYINPUT72), .B(new_n191), .C1(new_n427), .C2(new_n408), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n425), .A2(new_n426), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n188), .A2(new_n413), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n408), .B1(new_n188), .B2(G140), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT16), .ZN(new_n435));
  OAI211_X1 g249(.A(G146), .B(new_n433), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n407), .B1(new_n424), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n191), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n436), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n442), .B(new_n420), .C1(new_n421), .C2(new_n422), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n437), .A3(new_n406), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n439), .A2(new_n444), .A3(new_n276), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT25), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n439), .A2(new_n444), .A3(KEYINPUT25), .A4(new_n276), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n403), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n439), .A2(new_n444), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n450), .A2(G902), .A3(new_n402), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n400), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT9), .B(G234), .ZN(new_n455));
  OAI21_X1  g269(.A(G221), .B1(new_n455), .B2(G902), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n455), .A2(new_n401), .A3(G953), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT97), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G128), .B(G143), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(G134), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n461), .A2(KEYINPUT94), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(KEYINPUT94), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n225), .A2(new_n227), .A3(G122), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n224), .A2(G122), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n240), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT95), .ZN(new_n468));
  INV_X1    g282(.A(new_n464), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT14), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n464), .A2(KEYINPUT95), .A3(KEYINPUT14), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n465), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT96), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n473), .A2(new_n474), .B1(new_n470), .B2(new_n469), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n471), .A2(KEYINPUT96), .A3(new_n465), .A4(new_n472), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n467), .B1(new_n477), .B2(G107), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n460), .A2(new_n331), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT93), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n189), .A2(KEYINPUT13), .A3(G128), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n481), .B(KEYINPUT92), .C1(G128), .C2(new_n189), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT13), .B1(new_n189), .B2(G128), .ZN(new_n483));
  OAI221_X1 g297(.A(G134), .B1(KEYINPUT92), .B2(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n466), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n240), .B1(new_n464), .B2(new_n465), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n459), .B1(new_n478), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n489), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n240), .B1(new_n475), .B2(new_n476), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n458), .B(new_n491), .C1(new_n492), .C2(new_n467), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(new_n276), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G478), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(KEYINPUT15), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n496), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n490), .A2(new_n276), .A3(new_n493), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT20), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n313), .A2(KEYINPUT67), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT67), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G953), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n502), .A2(new_n504), .A3(G214), .A4(new_n316), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n189), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n319), .A2(G143), .A3(G214), .A4(new_n316), .ZN(new_n507));
  NAND2_X1  g321(.A1(KEYINPUT18), .A2(G131), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n507), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(KEYINPUT18), .A3(G131), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n188), .A2(G140), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n512), .A2(KEYINPUT88), .A3(G146), .A4(new_n409), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n430), .A2(new_n431), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT88), .B1(new_n434), .B2(G146), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n509), .B(new_n511), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT19), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n518), .A2(KEYINPUT89), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(KEYINPUT89), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n519), .B(new_n520), .C1(new_n427), .C2(new_n408), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n191), .B(new_n521), .C1(new_n412), .C2(new_n518), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n506), .A2(new_n507), .A3(new_n338), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n338), .B1(new_n506), .B2(new_n507), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n436), .B(new_n522), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n517), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(G113), .B(G122), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(new_n237), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n525), .A2(KEYINPUT17), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n441), .A2(new_n436), .A3(new_n532), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n524), .A2(KEYINPUT17), .A3(new_n525), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n529), .B(new_n517), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(G475), .A2(G902), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n501), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n537), .ZN(new_n539));
  AOI211_X1 g353(.A(KEYINPUT20), .B(new_n539), .C1(new_n531), .C2(new_n535), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G475), .ZN(new_n542));
  INV_X1    g356(.A(new_n525), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n523), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n415), .A2(new_n545), .A3(new_n532), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n529), .B1(new_n546), .B2(new_n517), .ZN(new_n547));
  AOI21_X1  g361(.A(G902), .B1(new_n547), .B2(KEYINPUT90), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n517), .B1(new_n533), .B2(new_n534), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n530), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT90), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n551), .A3(new_n535), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n542), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT91), .B1(new_n541), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n536), .A2(new_n537), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT20), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n536), .A2(new_n501), .A3(new_n537), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n550), .A2(new_n551), .A3(new_n535), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n276), .B1(new_n550), .B2(new_n551), .ZN(new_n560));
  OAI21_X1  g374(.A(G475), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT91), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n558), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n500), .B1(new_n554), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G469), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n196), .A2(new_n198), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n248), .A2(new_n566), .A3(KEYINPUT10), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT76), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n198), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n204), .A2(KEYINPUT76), .A3(new_n197), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n196), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n248), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT10), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT77), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n567), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n257), .A2(new_n206), .A3(new_n209), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT75), .B1(new_n262), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT75), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n329), .A2(new_n269), .A3(new_n579), .A4(new_n257), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AOI211_X1 g395(.A(new_n575), .B(KEYINPUT10), .C1(new_n571), .C2(new_n248), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n576), .A2(new_n581), .A3(new_n351), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT78), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n248), .A2(new_n566), .A3(KEYINPUT10), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT10), .B1(new_n571), .B2(new_n248), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n586), .B1(new_n587), .B2(KEYINPUT77), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(new_n582), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT78), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n589), .A2(new_n590), .A3(new_n351), .A4(new_n581), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n572), .B1(new_n566), .B2(new_n248), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n340), .ZN(new_n594));
  XOR2_X1   g408(.A(new_n594), .B(KEYINPUT12), .Z(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(G110), .B(G140), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT73), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n319), .A2(G227), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n598), .B(new_n599), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(KEYINPUT74), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n351), .B1(new_n589), .B2(new_n581), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n600), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n585), .B2(new_n591), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n604), .B1(new_n606), .B2(KEYINPUT79), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT79), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n608), .B(new_n605), .C1(new_n585), .C2(new_n591), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n602), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n565), .B1(new_n610), .B2(new_n276), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT80), .B(G469), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n606), .A2(new_n595), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n600), .B1(new_n592), .B2(new_n604), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n276), .B(new_n612), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n456), .B(new_n564), .C1(new_n611), .C2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n328), .A2(new_n454), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  INV_X1    g434(.A(new_n456), .ZN(new_n621));
  INV_X1    g435(.A(new_n601), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n592), .B2(new_n595), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n592), .A2(new_n600), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n603), .B1(new_n624), .B2(new_n608), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n606), .A2(KEYINPUT79), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(G469), .B1(new_n627), .B2(G902), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n621), .B1(new_n628), .B2(new_n615), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n376), .A2(new_n276), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(G472), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n378), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(G472), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n376), .B2(new_n276), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n632), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n634), .A2(new_n452), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n629), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n456), .B1(new_n611), .B2(new_n616), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT100), .B1(new_n642), .B2(new_n638), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n285), .B1(new_n311), .B2(new_n302), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n325), .B1(new_n646), .B2(new_n299), .ZN(new_n647));
  INV_X1    g461(.A(new_n323), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT101), .B1(new_n494), .B2(new_n495), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n494), .A2(KEYINPUT101), .A3(new_n495), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n477), .A2(G107), .ZN(new_n653));
  INV_X1    g467(.A(new_n467), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n458), .B1(new_n655), .B2(new_n491), .ZN(new_n656));
  INV_X1    g470(.A(new_n493), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n652), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n490), .A2(KEYINPUT33), .A3(new_n493), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n495), .A2(G902), .ZN(new_n661));
  AOI22_X1  g475(.A1(new_n650), .A2(new_n651), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n554), .A2(new_n563), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n647), .A2(new_n648), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n645), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT34), .B(G104), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  INV_X1    g482(.A(new_n500), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n558), .A2(new_n561), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n647), .A2(new_n648), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n644), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n240), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT102), .B(KEYINPUT35), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  NOR2_X1   g490(.A1(new_n327), .A2(new_n617), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n443), .B2(new_n437), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n424), .A2(KEYINPUT103), .A3(new_n438), .ZN(new_n680));
  OAI22_X1  g494(.A1(new_n679), .A2(new_n680), .B1(KEYINPUT36), .B2(new_n407), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT103), .B1(new_n424), .B2(new_n438), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n443), .A2(new_n678), .A3(new_n437), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n407), .A2(KEYINPUT36), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n402), .A2(G902), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n681), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n449), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n634), .A2(new_n690), .A3(new_n637), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n677), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT37), .B(G110), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G12));
  XOR2_X1   g509(.A(KEYINPUT104), .B(G900), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n320), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n318), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n558), .A2(new_n561), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n669), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n400), .A2(new_n689), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n629), .A2(new_n647), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  XNOR2_X1  g517(.A(new_n698), .B(KEYINPUT39), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n629), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT106), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT40), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n705), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n309), .A2(new_n312), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT38), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n379), .A2(new_n381), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n358), .B1(new_n341), .B2(new_n348), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n374), .B1(new_n369), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n365), .A2(KEYINPUT105), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n276), .ZN(new_n718));
  AOI21_X1  g532(.A(KEYINPUT105), .B1(new_n365), .B2(new_n716), .ZN(new_n719));
  OAI21_X1  g533(.A(G472), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n554), .A2(new_n563), .A3(new_n500), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n324), .A3(new_n689), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n713), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n708), .A2(new_n711), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT107), .B(G143), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G45));
  INV_X1    g542(.A(new_n698), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n662), .A2(new_n663), .A3(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n629), .A2(new_n647), .A3(new_n701), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G146), .ZN(G48));
  AOI211_X1 g546(.A(new_n323), .B(new_n325), .C1(new_n646), .C2(new_n299), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n276), .B1(new_n613), .B2(new_n614), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(G469), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n456), .A3(new_n615), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n736), .A2(new_n400), .A3(new_n453), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n733), .A2(new_n737), .A3(new_n664), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT41), .B(G113), .Z(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT108), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n738), .B(new_n740), .ZN(G15));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n735), .A2(new_n456), .A3(new_n615), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n454), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n742), .B1(new_n672), .B2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n733), .A2(new_n737), .A3(KEYINPUT109), .A4(new_n671), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  INV_X1    g562(.A(new_n299), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n304), .A2(new_n305), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n286), .B1(new_n750), .B2(new_n283), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n324), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n399), .A2(G472), .ZN(new_n753));
  INV_X1    g567(.A(new_n381), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n380), .B1(new_n376), .B2(new_n377), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n690), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n735), .A2(new_n648), .A3(new_n456), .A4(new_n615), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n554), .A2(new_n563), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n759), .A2(new_n500), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G119), .ZN(G21));
  INV_X1    g577(.A(new_n383), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT28), .B1(new_n369), .B2(new_n715), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n382), .B1(new_n359), .B2(new_n371), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n374), .B1(new_n767), .B2(KEYINPUT110), .ZN(new_n768));
  OAI211_X1 g582(.A(KEYINPUT110), .B(new_n383), .C1(new_n386), .C2(new_n387), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n366), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT111), .B(new_n366), .C1(new_n768), .C2(new_n770), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n368), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n636), .B1(new_n775), .B2(new_n377), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n743), .A2(new_n776), .A3(new_n452), .A4(new_n648), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n324), .B(new_n723), .C1(new_n749), .C2(new_n751), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT112), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n364), .B1(new_n388), .B2(new_n780), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n781), .A2(new_n769), .B1(KEYINPUT31), .B2(new_n365), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n368), .B1(new_n782), .B2(KEYINPUT111), .ZN(new_n783));
  INV_X1    g597(.A(new_n774), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n377), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n452), .A3(new_n631), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n759), .ZN(new_n787));
  AOI211_X1 g601(.A(new_n325), .B(new_n722), .C1(new_n646), .C2(new_n299), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n779), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G122), .ZN(G24));
  AOI211_X1 g606(.A(new_n636), .B(new_n689), .C1(new_n775), .C2(new_n377), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n793), .A2(new_n647), .A3(new_n730), .A4(new_n743), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G125), .ZN(G27));
  AND3_X1   g609(.A1(new_n712), .A2(new_n629), .A3(new_n324), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(KEYINPUT42), .A3(new_n454), .A4(new_n730), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n325), .B1(new_n309), .B2(new_n312), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(new_n454), .A3(new_n629), .A4(new_n730), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT42), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G131), .ZN(G33));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n804), .B1(new_n669), .B2(new_n699), .ZN(new_n805));
  INV_X1    g619(.A(new_n699), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(KEYINPUT113), .A3(new_n500), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n798), .A2(new_n454), .A3(new_n629), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G134), .ZN(G36));
  INV_X1    g624(.A(new_n798), .ZN(new_n811));
  INV_X1    g625(.A(new_n659), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT33), .B1(new_n490), .B2(new_n493), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n661), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n651), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n814), .B1(new_n815), .B2(new_n649), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n663), .ZN(new_n817));
  XOR2_X1   g631(.A(new_n817), .B(KEYINPUT43), .Z(new_n818));
  AOI21_X1  g632(.A(new_n689), .B1(new_n634), .B2(new_n637), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT44), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n811), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n818), .A2(KEYINPUT44), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT45), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n565), .B1(new_n610), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n825), .B2(new_n610), .ZN(new_n827));
  NAND2_X1  g641(.A1(G469), .A2(G902), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT46), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n615), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n829), .A2(new_n830), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n456), .B(new_n704), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n834), .A2(KEYINPUT114), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(KEYINPUT114), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n824), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(new_n333), .ZN(G39));
  NAND3_X1  g652(.A1(new_n760), .A2(new_n816), .A3(new_n698), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n839), .A2(new_n756), .A3(new_n452), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n798), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n456), .B1(new_n832), .B2(new_n833), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT47), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(KEYINPUT47), .B(new_n456), .C1(new_n832), .C2(new_n833), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n841), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(new_n411), .ZN(G42));
  NOR4_X1   g661(.A1(new_n817), .A2(new_n453), .A3(new_n325), .A4(new_n621), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n735), .A2(new_n615), .ZN(new_n849));
  XOR2_X1   g663(.A(new_n849), .B(KEYINPUT49), .Z(new_n850));
  NAND4_X1  g664(.A1(new_n713), .A2(new_n721), .A3(new_n848), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n778), .A2(new_n786), .A3(KEYINPUT112), .A4(new_n759), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n789), .B1(new_n787), .B2(new_n788), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n693), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n619), .A2(new_n762), .A3(new_n738), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n699), .A2(new_n500), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n756), .A2(new_n690), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n785), .A2(new_n631), .A3(new_n690), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n859), .B1(new_n860), .B2(new_n839), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n629), .A3(new_n798), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n809), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n797), .B2(new_n801), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n760), .A2(new_n669), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(new_n309), .A3(new_n312), .A4(new_n326), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT116), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n866), .A2(KEYINPUT116), .ZN(new_n869));
  OR3_X1    g683(.A1(new_n868), .A2(new_n644), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT115), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(new_n662), .B2(new_n663), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n760), .A2(new_n816), .A3(KEYINPUT115), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n327), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n645), .A2(new_n876), .B1(new_n745), .B2(new_n746), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n857), .A2(new_n864), .A3(new_n870), .A4(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n702), .A2(new_n731), .A3(new_n794), .ZN(new_n879));
  INV_X1    g693(.A(new_n449), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n698), .B(KEYINPUT117), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n687), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n714), .B2(new_n720), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n624), .A2(new_n608), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n626), .A3(new_n604), .ZN(new_n885));
  AOI21_X1  g699(.A(G902), .B1(new_n885), .B2(new_n602), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n615), .B1(new_n886), .B2(new_n565), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n883), .A2(new_n887), .A3(new_n456), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT118), .B1(new_n888), .B2(new_n778), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n788), .A2(new_n890), .A3(new_n629), .A4(new_n883), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n879), .A2(KEYINPUT52), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT52), .B1(new_n879), .B2(new_n892), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n852), .B1(new_n878), .B2(new_n895), .ZN(new_n896));
  AOI22_X1  g710(.A1(new_n665), .A2(new_n737), .B1(new_n758), .B2(new_n761), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n791), .A2(new_n897), .A3(new_n619), .A4(new_n693), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n876), .A2(new_n641), .A3(new_n643), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n747), .A2(new_n899), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n868), .A2(new_n644), .A3(new_n869), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT52), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n889), .A2(new_n891), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n702), .A2(new_n731), .A3(new_n794), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n879), .A2(new_n892), .A3(KEYINPUT52), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n702), .A2(new_n794), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n852), .B1(new_n909), .B2(KEYINPUT52), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n902), .A2(new_n908), .A3(new_n864), .A4(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n896), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n896), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT53), .B1(new_n909), .B2(KEYINPUT52), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n878), .A2(new_n895), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n913), .B1(new_n917), .B2(new_n912), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT51), .ZN(new_n919));
  INV_X1    g733(.A(new_n318), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n818), .A2(new_n452), .A3(new_n920), .A4(new_n776), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n743), .B(new_n325), .C1(KEYINPUT119), .C2(KEYINPUT50), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n713), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT50), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OR3_X1    g741(.A1(new_n923), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n811), .A2(new_n736), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n929), .A2(new_n920), .A3(new_n818), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n793), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n927), .B1(new_n923), .B2(new_n924), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n929), .A2(new_n452), .A3(new_n920), .A4(new_n721), .ZN(new_n933));
  OR3_X1    g747(.A1(new_n933), .A2(new_n760), .A3(new_n816), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n928), .A2(new_n931), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n844), .B(new_n845), .C1(new_n456), .C2(new_n849), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n921), .A2(new_n811), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n919), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n930), .A2(new_n454), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT48), .Z(new_n941));
  NAND2_X1  g755(.A1(new_n647), .A2(new_n743), .ZN(new_n942));
  INV_X1    g756(.A(new_n664), .ZN(new_n943));
  OAI221_X1 g757(.A(new_n314), .B1(new_n942), .B2(new_n921), .C1(new_n933), .C2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n939), .A2(new_n945), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n935), .A2(new_n919), .A3(new_n938), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n918), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(G952), .A2(G953), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n851), .B1(new_n948), .B2(new_n949), .ZN(G75));
  NOR2_X1   g764(.A1(new_n319), .A2(G952), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n276), .B1(new_n896), .B2(new_n911), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n954), .A2(new_n308), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n295), .B(new_n296), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT55), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT56), .B1(new_n958), .B2(KEYINPUT121), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(KEYINPUT121), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n952), .B1(new_n955), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT56), .B1(new_n953), .B2(new_n285), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT120), .ZN(new_n963));
  OR3_X1    g777(.A1(new_n962), .A2(new_n963), .A3(new_n958), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n962), .B2(new_n958), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(G51));
  XOR2_X1   g780(.A(new_n828), .B(KEYINPUT57), .Z(new_n967));
  INV_X1    g781(.A(new_n913), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n912), .B1(new_n896), .B2(new_n911), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n614), .B2(new_n613), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n954), .A2(new_n827), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n951), .B1(new_n971), .B2(new_n972), .ZN(G54));
  NAND2_X1  g787(.A1(KEYINPUT58), .A2(G475), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n953), .A2(new_n536), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n536), .B1(new_n953), .B2(new_n975), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n976), .A2(new_n977), .A3(new_n951), .ZN(G60));
  NAND2_X1  g792(.A1(G478), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT59), .Z(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n660), .B1(new_n918), .B2(new_n981), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n660), .B(new_n981), .C1(new_n968), .C2(new_n969), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n952), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n982), .A2(new_n984), .ZN(G63));
  NAND2_X1  g799(.A1(G217), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT122), .Z(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT60), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(new_n896), .B2(new_n911), .ZN(new_n989));
  INV_X1    g803(.A(new_n450), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n952), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT123), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT123), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n993), .B(new_n952), .C1(new_n989), .C2(new_n990), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n681), .A2(new_n685), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n989), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n992), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT61), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT124), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n997), .A2(KEYINPUT61), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1001), .B1(new_n1002), .B2(new_n991), .ZN(new_n1003));
  OR2_X1    g817(.A1(new_n989), .A2(new_n990), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n999), .B1(new_n989), .B2(new_n996), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1004), .A2(new_n1005), .A3(KEYINPUT124), .A4(new_n952), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1000), .A2(new_n1007), .ZN(G66));
  OAI21_X1  g822(.A(G953), .B1(new_n321), .B2(new_n201), .ZN(new_n1009));
  INV_X1    g823(.A(new_n319), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1009), .B1(new_n902), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(G898), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n295), .B1(new_n1012), .B2(new_n1010), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(KEYINPUT125), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1011), .B(new_n1014), .ZN(G69));
  AOI21_X1  g829(.A(new_n319), .B1(G227), .B2(G900), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(KEYINPUT127), .ZN(new_n1017));
  OR2_X1    g831(.A1(new_n1016), .A2(KEYINPUT127), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n349), .B1(new_n356), .B2(KEYINPUT30), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n521), .B1(new_n412), .B2(new_n518), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1010), .A2(G900), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n837), .A2(new_n846), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n835), .A2(new_n836), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1025), .A2(new_n454), .A3(new_n788), .ZN(new_n1026));
  AND3_X1   g840(.A1(new_n802), .A2(new_n809), .A3(new_n879), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1023), .B1(new_n1029), .B2(new_n319), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1021), .B(KEYINPUT126), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1031), .ZN(new_n1032));
  OAI22_X1  g846(.A1(new_n873), .A2(new_n875), .B1(new_n669), .B2(new_n760), .ZN(new_n1033));
  NAND4_X1  g847(.A1(new_n706), .A2(new_n454), .A3(new_n798), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(KEYINPUT62), .B1(new_n726), .B2(new_n879), .ZN(new_n1035));
  AND3_X1   g849(.A1(new_n726), .A2(KEYINPUT62), .A3(new_n879), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n1024), .B(new_n1034), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1032), .B1(new_n1037), .B2(new_n319), .ZN(new_n1038));
  OAI211_X1 g852(.A(new_n1017), .B(new_n1018), .C1(new_n1030), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1037), .A2(new_n319), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1040), .A2(new_n1031), .ZN(new_n1041));
  OAI211_X1 g855(.A(new_n1022), .B(new_n1021), .C1(new_n1028), .C2(new_n1010), .ZN(new_n1042));
  NAND4_X1  g856(.A1(new_n1041), .A2(KEYINPUT127), .A3(new_n1016), .A4(new_n1042), .ZN(new_n1043));
  AND2_X1   g857(.A1(new_n1039), .A2(new_n1043), .ZN(G72));
  NAND3_X1  g858(.A1(new_n357), .A2(new_n359), .A3(new_n374), .ZN(new_n1045));
  NAND4_X1  g859(.A1(new_n1024), .A2(new_n902), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1046));
  NAND2_X1  g860(.A1(G472), .A2(G902), .ZN(new_n1047));
  XOR2_X1   g861(.A(new_n1047), .B(KEYINPUT63), .Z(new_n1048));
  AOI21_X1  g862(.A(new_n1045), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g863(.A(new_n365), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1048), .B1(new_n1050), .B2(new_n398), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n952), .B1(new_n917), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n857), .A2(new_n870), .A3(new_n877), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1048), .B1(new_n1037), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n374), .B1(new_n357), .B2(new_n359), .ZN(new_n1055));
  AOI211_X1 g869(.A(new_n1049), .B(new_n1052), .C1(new_n1054), .C2(new_n1055), .ZN(G57));
endmodule


