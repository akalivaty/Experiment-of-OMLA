//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(KEYINPUT3), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n462), .A2(G137), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n460), .A2(new_n461), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(new_n463), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(KEYINPUT69), .A3(new_n468), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT66), .ZN(new_n474));
  OR2_X1    g049(.A1(new_n473), .A2(KEYINPUT66), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n465), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n474), .B(new_n475), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n479), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(KEYINPUT67), .B1(new_n479), .B2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n471), .B(new_n472), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT70), .Z(G160));
  NAND3_X1  g058(.A1(new_n462), .A2(G2105), .A3(new_n465), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT71), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n462), .A2(new_n486), .A3(G2105), .A4(new_n465), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n490));
  OR2_X1    g065(.A1(new_n463), .A2(G112), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n490), .A2(G136), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  NAND4_X1  g071(.A1(new_n462), .A2(G138), .A3(new_n463), .A4(new_n465), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(new_n463), .A3(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n477), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n462), .A2(G126), .A3(G2105), .A4(new_n465), .ZN(new_n504));
  OR2_X1    g079(.A1(G102), .A2(G2105), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n505), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  AND2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT72), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT72), .A2(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT6), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n513), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT73), .B(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n522), .B1(new_n516), .B2(new_n518), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n513), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n528));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(KEYINPUT72), .A2(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n521), .A2(new_n524), .A3(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND2_X1  g110(.A1(new_n519), .A2(G89), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT6), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n530), .B2(new_n531), .ZN(new_n538));
  OAI211_X1 g113(.A(G51), .B(G543), .C1(new_n538), .C2(new_n517), .ZN(new_n539));
  INV_X1    g114(.A(new_n512), .ZN(new_n540));
  NAND2_X1  g115(.A1(KEYINPUT5), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g117(.A1(G63), .A2(G651), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT7), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n546), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n542), .A2(new_n543), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n536), .A2(new_n539), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT74), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n536), .A2(new_n551), .A3(new_n539), .A4(new_n548), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n550), .A2(new_n552), .ZN(G168));
  XNOR2_X1  g128(.A(KEYINPUT75), .B(G90), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n519), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n523), .A2(G52), .ZN(new_n556));
  NAND2_X1  g131(.A1(G77), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G64), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n513), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(new_n532), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n555), .A2(new_n556), .A3(new_n560), .ZN(G301));
  INV_X1    g136(.A(G301), .ZN(G171));
  XOR2_X1   g137(.A(KEYINPUT77), .B(G81), .Z(new_n563));
  NAND2_X1  g138(.A1(new_n519), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g139(.A(KEYINPUT76), .B(G43), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n523), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G68), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G56), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n513), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(new_n532), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n564), .A2(new_n566), .A3(G860), .A4(new_n570), .ZN(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND4_X1  g149(.A1(G319), .A2(G483), .A3(G661), .A4(new_n574), .ZN(G188));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  XNOR2_X1  g151(.A(KEYINPUT78), .B(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n513), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(G91), .A2(new_n519), .B1(new_n578), .B2(G651), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT9), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n523), .A2(new_n580), .A3(G53), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n580), .B1(new_n523), .B2(G53), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(G299));
  AND2_X1   g159(.A1(new_n550), .A2(new_n552), .ZN(G286));
  INV_X1    g160(.A(G74), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n529), .B1(new_n513), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n519), .B2(G87), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n523), .A2(G49), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n588), .A2(KEYINPUT79), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(KEYINPUT79), .B1(new_n588), .B2(new_n589), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(new_n523), .A2(G48), .ZN(new_n593));
  OAI211_X1 g168(.A(G86), .B(new_n542), .C1(new_n538), .C2(new_n517), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n540), .B2(new_n541), .ZN(new_n596));
  AND2_X1   g171(.A1(G73), .A2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n532), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n593), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G60), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n513), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(new_n532), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT81), .ZN(new_n606));
  AOI22_X1  g181(.A1(G47), .A2(new_n523), .B1(new_n519), .B2(G85), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n523), .A2(G54), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G66), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n513), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G651), .ZN(new_n614));
  AND2_X1   g189(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g190(.A(G92), .B(new_n542), .C1(new_n538), .C2(new_n517), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(KEYINPUT82), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT10), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n519), .A2(new_n619), .A3(G92), .ZN(new_n620));
  AND3_X1   g195(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n618), .B1(new_n617), .B2(new_n620), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n609), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n609), .B1(new_n624), .B2(G868), .ZN(G321));
  NOR2_X1   g201(.A1(G299), .A2(G868), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g203(.A(new_n627), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n624), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND3_X1  g206(.A1(new_n564), .A2(new_n566), .A3(new_n570), .ZN(new_n632));
  INV_X1    g207(.A(G868), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n623), .A2(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(new_n633), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n488), .A2(G123), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT84), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n490), .A2(G135), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n463), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n639), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n643), .A2(G2096), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n467), .A2(new_n463), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n646), .A2(new_n477), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT12), .Z(new_n648));
  XOR2_X1   g223(.A(KEYINPUT83), .B(G2100), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT13), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n648), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n644), .A2(new_n645), .A3(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT85), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2430), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(KEYINPUT14), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XOR2_X1   g236(.A(G1341), .B(G1348), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n659), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2443), .B(G2446), .Z(new_n665));
  OAI21_X1  g240(.A(G14), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n665), .B2(new_n664), .ZN(G401));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT17), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT87), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2084), .B(G2090), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(new_n670), .B2(new_n668), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n671), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n672), .B2(new_n674), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT88), .Z(new_n677));
  OR3_X1    g252(.A1(new_n669), .A2(new_n670), .A3(new_n673), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n670), .A2(new_n668), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n679), .A2(new_n673), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT86), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT18), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n677), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2096), .B(G2100), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT89), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n687), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n694), .A2(new_n691), .A3(new_n687), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n692), .B1(new_n691), .B2(new_n687), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1981), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT91), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n700), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n703), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n704), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n704), .B2(new_n708), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(G229));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NOR2_X1   g289(.A1(G164), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G27), .B2(new_n714), .ZN(new_n716));
  INV_X1    g291(.A(G2078), .ZN(new_n717));
  INV_X1    g292(.A(G1961), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n719), .A2(G5), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G301), .B2(G16), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n716), .A2(new_n717), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT30), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n723), .A2(G28), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n714), .B1(new_n723), .B2(G28), .ZN(new_n725));
  AND2_X1   g300(.A1(KEYINPUT31), .A2(G11), .ZN(new_n726));
  NOR2_X1   g301(.A1(KEYINPUT31), .A2(G11), .ZN(new_n727));
  OAI22_X1  g302(.A1(new_n724), .A2(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(G16), .A2(G19), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n632), .B2(new_n719), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT97), .B(G1341), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n722), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(G115), .A2(G2104), .ZN(new_n734));
  INV_X1    g309(.A(G127), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n477), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT25), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n736), .A2(G2105), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n490), .A2(G139), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n741), .A2(new_n742), .A3(KEYINPUT100), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(KEYINPUT100), .B1(new_n741), .B2(new_n742), .ZN(new_n745));
  OAI21_X1  g320(.A(G29), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G33), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(G29), .B2(new_n747), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n733), .B1(new_n714), .B2(new_n643), .C1(G2072), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(G2072), .ZN(new_n750));
  NAND2_X1  g325(.A1(G162), .A2(G29), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G29), .B2(G35), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT29), .B(G2090), .Z(new_n753));
  OAI21_X1  g328(.A(new_n750), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT101), .ZN(new_n756));
  INV_X1    g331(.A(G105), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n646), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n467), .A2(KEYINPUT101), .A3(G105), .A4(new_n463), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n490), .A2(G141), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT26), .Z(new_n763));
  NAND3_X1  g338(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  AND3_X1   g339(.A1(new_n485), .A2(G129), .A3(new_n487), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(new_n714), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n714), .B2(G32), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT27), .B(G1996), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR4_X1   g345(.A1(new_n749), .A2(new_n754), .A3(new_n755), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n768), .A2(new_n769), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT102), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n714), .A2(G26), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT28), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT99), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n485), .A2(new_n487), .ZN(new_n777));
  INV_X1    g352(.A(G128), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n485), .A2(KEYINPUT99), .A3(G128), .A4(new_n487), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n782));
  INV_X1    g357(.A(G116), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G2105), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n490), .A2(G140), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT98), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n490), .A2(KEYINPUT98), .A3(G140), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n781), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n775), .B1(new_n791), .B2(new_n714), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n773), .B1(G2067), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n719), .A2(G21), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G168), .B2(new_n719), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G1966), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT103), .Z(new_n797));
  OAI22_X1  g372(.A1(new_n716), .A2(new_n717), .B1(new_n718), .B2(new_n721), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n719), .A2(G20), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT104), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT23), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G299), .B2(G16), .ZN(new_n802));
  INV_X1    g377(.A(G1956), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n795), .A2(G1966), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n730), .A2(new_n731), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n798), .A2(new_n804), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n771), .A2(new_n793), .A3(new_n797), .A4(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(KEYINPUT24), .A2(G34), .ZN(new_n809));
  NAND2_X1  g384(.A1(KEYINPUT24), .A2(G34), .ZN(new_n810));
  AOI21_X1  g385(.A(G29), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G160), .B2(G29), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G2084), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n719), .A2(G4), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n624), .B2(new_n719), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(G1348), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(G1348), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n816), .B(new_n817), .C1(G2067), .C2(new_n792), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n808), .A2(new_n813), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n714), .A2(G25), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n462), .A2(G131), .A3(new_n463), .A4(new_n465), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT92), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n485), .A2(G119), .A3(new_n487), .ZN(new_n823));
  OR2_X1    g398(.A1(G95), .A2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n824), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT93), .Z(new_n826));
  NAND3_X1  g401(.A1(new_n822), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT94), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT94), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n822), .A2(new_n829), .A3(new_n823), .A4(new_n826), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n820), .B1(new_n832), .B2(new_n714), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT95), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT35), .B(G1991), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n719), .A2(G6), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n599), .B(KEYINPUT80), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n838), .B2(new_n719), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT32), .B(G1981), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n719), .A2(G22), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(G166), .B2(new_n719), .ZN(new_n844));
  INV_X1    g419(.A(G1971), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n719), .A2(G23), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n588), .A2(new_n589), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n847), .B1(new_n849), .B2(new_n719), .ZN(new_n850));
  XNOR2_X1  g425(.A(KEYINPUT33), .B(G1976), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n841), .A2(new_n842), .A3(new_n846), .A4(new_n852), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(KEYINPUT34), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(KEYINPUT34), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT96), .ZN(new_n856));
  INV_X1    g431(.A(G290), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G16), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(G16), .B2(G24), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n856), .B1(new_n859), .B2(new_n705), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(new_n705), .B2(new_n859), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n836), .A2(new_n854), .A3(new_n855), .A4(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT36), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n819), .A2(new_n864), .A3(new_n865), .ZN(G311));
  NAND3_X1  g441(.A1(new_n819), .A2(new_n864), .A3(new_n865), .ZN(G150));
  NOR2_X1   g442(.A1(new_n623), .A2(new_n630), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT38), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n519), .A2(G93), .ZN(new_n870));
  NAND2_X1  g445(.A1(G80), .A2(G543), .ZN(new_n871));
  INV_X1    g446(.A(G67), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n513), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n532), .ZN(new_n874));
  OAI211_X1 g449(.A(G55), .B(G543), .C1(new_n538), .C2(new_n517), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n870), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n632), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n869), .B(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(KEYINPUT39), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(KEYINPUT39), .ZN(new_n880));
  XNOR2_X1  g455(.A(KEYINPUT105), .B(G860), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n881), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n876), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(KEYINPUT37), .Z(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(G145));
  NAND2_X1  g461(.A1(new_n490), .A2(G142), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n463), .A2(G118), .ZN(new_n888));
  OAI21_X1  g463(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n889));
  INV_X1    g464(.A(G130), .ZN(new_n890));
  OAI221_X1 g465(.A(new_n887), .B1(new_n888), .B2(new_n889), .C1(new_n777), .C2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n648), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n741), .A2(new_n742), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n765), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n894), .A2(new_n897), .A3(new_n898), .A4(new_n743), .ZN(new_n899));
  OAI22_X1  g474(.A1(new_n744), .A2(new_n745), .B1(new_n764), .B2(new_n765), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n828), .A2(KEYINPUT106), .A3(new_n830), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT106), .B1(new_n828), .B2(new_n830), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n899), .A2(new_n900), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n902), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n790), .B(new_n509), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n909), .B1(new_n905), .B2(new_n908), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n893), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n909), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n903), .A2(new_n901), .A3(new_n904), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n907), .B1(new_n906), .B2(new_n902), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n892), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n912), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(G160), .B(new_n495), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(new_n643), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n922), .A2(new_n912), .A3(new_n919), .A4(new_n918), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(G37), .B1(new_n920), .B2(new_n923), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n930), .A2(KEYINPUT108), .A3(new_n926), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n929), .A2(KEYINPUT40), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT40), .B1(new_n929), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(G395));
  NAND2_X1  g509(.A1(new_n876), .A2(new_n633), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n632), .A2(new_n876), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n632), .A2(new_n876), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT109), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(new_n635), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n941));
  INV_X1    g516(.A(G299), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n623), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g518(.A(G299), .B(new_n615), .C1(new_n621), .C2(new_n622), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n941), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n940), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT41), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n943), .A2(new_n950), .A3(new_n944), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n944), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n616), .A2(KEYINPUT82), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n619), .B1(new_n519), .B2(G92), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT10), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n617), .A2(new_n620), .A3(new_n618), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(G299), .B1(new_n958), .B2(new_n615), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT110), .B1(new_n953), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n946), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n952), .B1(new_n961), .B2(KEYINPUT41), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n949), .B1(new_n940), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(G305), .A2(G303), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n838), .A2(G166), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(G290), .A2(new_n849), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n606), .A2(new_n848), .A3(new_n607), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n964), .A2(new_n965), .A3(new_n967), .A4(new_n968), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT42), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n963), .B(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n935), .B1(new_n974), .B2(new_n633), .ZN(G295));
  OAI21_X1  g550(.A(new_n935), .B1(new_n974), .B2(new_n633), .ZN(G331));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n977));
  NAND2_X1  g552(.A1(G168), .A2(G171), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n550), .A2(new_n552), .A3(G301), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n938), .A3(new_n979), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n550), .A2(new_n552), .A3(G301), .ZN(new_n981));
  AOI21_X1  g556(.A(G301), .B1(new_n550), .B2(new_n552), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n877), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n943), .A2(new_n944), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(KEYINPUT41), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n972), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n950), .B1(new_n980), .B2(new_n983), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n961), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n977), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n984), .A2(KEYINPUT41), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n948), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n992), .A2(KEYINPUT112), .A3(new_n972), .A4(new_n986), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n995));
  INV_X1    g570(.A(new_n984), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n948), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n962), .B2(new_n996), .ZN(new_n998));
  INV_X1    g573(.A(new_n972), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT41), .B1(new_n945), .B2(new_n947), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n996), .B1(new_n1001), .B2(new_n951), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n961), .A2(new_n984), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n995), .B(new_n999), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n994), .B(new_n925), .C1(new_n1000), .C2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT43), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1008));
  AOI21_X1  g583(.A(G37), .B1(new_n1008), .B2(new_n972), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1007), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(KEYINPUT43), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT43), .B1(new_n990), .B2(new_n993), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1014), .B(new_n925), .C1(new_n1000), .C2(new_n1005), .ZN(new_n1015));
  AOI211_X1 g590(.A(new_n1012), .B(KEYINPUT44), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n972), .B(new_n997), .C1(new_n962), .C2(new_n996), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n925), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT111), .B1(new_n1008), .B2(new_n972), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1018), .B1(new_n1019), .B2(new_n1004), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT43), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1015), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT113), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1011), .B1(new_n1016), .B2(new_n1024), .ZN(G397));
  INV_X1    g600(.A(KEYINPUT127), .ZN(new_n1026));
  XOR2_X1   g601(.A(new_n766), .B(G1996), .Z(new_n1027));
  INV_X1    g602(.A(G1384), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n501), .B1(new_n497), .B2(KEYINPUT4), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1028), .B1(new_n1029), .B2(new_n507), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n471), .A2(new_n472), .ZN(new_n1033));
  OAI21_X1  g608(.A(G40), .B1(new_n480), .B2(new_n481), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1027), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n1037));
  INV_X1    g612(.A(G2067), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1038), .B1(new_n781), .B2(new_n789), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n781), .A2(new_n789), .A3(new_n1038), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1037), .B1(new_n1042), .B2(new_n1035), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1041), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1037), .B(new_n1035), .C1(new_n1044), .C2(new_n1039), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1036), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(KEYINPUT115), .B(new_n1036), .C1(new_n1043), .C2(new_n1046), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n832), .A2(new_n835), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n832), .A2(new_n835), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1035), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1049), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n857), .A2(new_n705), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G290), .A2(G1986), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1035), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1966), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1032), .ZN(new_n1060));
  INV_X1    g635(.A(G40), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n475), .A2(new_n474), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n465), .A2(new_n476), .A3(G125), .ZN(new_n1063));
  OAI21_X1  g638(.A(G2105), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT67), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n479), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1061), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n466), .A2(KEYINPUT69), .A3(new_n468), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT69), .B1(new_n466), .B2(new_n468), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1031), .A2(G1384), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n1029), .B2(new_n507), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1068), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1059), .B1(new_n1060), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1034), .A2(new_n1033), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT50), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1077), .B(new_n1028), .C1(new_n1029), .C2(new_n507), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1030), .A2(KEYINPUT50), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT120), .B(G2084), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1075), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G8), .ZN(new_n1083));
  NOR2_X1   g658(.A1(G168), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT51), .B1(new_n1084), .B2(KEYINPUT125), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1082), .A2(G8), .ZN(new_n1087));
  NAND2_X1  g662(.A1(G286), .A2(G8), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1083), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT125), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1090), .A2(new_n1093), .A3(new_n1084), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1085), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT62), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n599), .A2(G1981), .ZN(new_n1097));
  INV_X1    g672(.A(G1981), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n593), .A2(new_n1098), .A3(new_n594), .A4(new_n598), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT49), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1384), .B1(new_n503), .B2(new_n508), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1102), .A2(new_n1104), .A3(G8), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1097), .A2(KEYINPUT49), .A3(new_n1099), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1097), .A2(KEYINPUT119), .A3(KEYINPUT49), .A4(new_n1099), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n588), .A2(G1976), .A3(new_n589), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT118), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(G8), .A3(new_n1104), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1105), .A2(new_n1110), .B1(new_n1113), .B2(KEYINPUT52), .ZN(new_n1114));
  INV_X1    g689(.A(G1976), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT52), .B1(G288), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1083), .B1(new_n1076), .B2(new_n1103), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(new_n1112), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n509), .A2(new_n1119), .A3(new_n1072), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1073), .A2(KEYINPUT116), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1076), .A2(new_n1120), .A3(new_n1032), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n845), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT117), .B(G2090), .Z(new_n1124));
  NAND4_X1  g699(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .A4(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1083), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(G303), .A2(G8), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT55), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1114), .B(new_n1118), .C1(new_n1126), .C2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT53), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n1122), .B2(G2078), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1060), .A2(new_n1074), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1133), .A2(KEYINPUT53), .A3(new_n717), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1079), .A2(new_n1071), .A3(new_n1068), .A4(new_n1078), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n718), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1132), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(G171), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1135), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1139), .A2(new_n1124), .B1(new_n1122), .B2(new_n845), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1140), .A2(new_n1083), .A3(new_n1128), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1130), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1143), .B(new_n1085), .C1(new_n1089), .C2(new_n1094), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1096), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1110), .A2(new_n1117), .A3(new_n1102), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1113), .A2(KEYINPUT52), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1146), .A2(new_n1118), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1128), .B1(new_n1140), .B2(new_n1083), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1129), .B1(new_n1152), .B2(G8), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1146), .A2(new_n1147), .A3(new_n1118), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT121), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1090), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1141), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1151), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1090), .A2(G168), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1149), .A2(new_n1148), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT63), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1158), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1146), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1115), .B1(new_n590), .B2(new_n591), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1099), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1167), .A2(new_n1117), .B1(new_n1141), .B2(new_n1148), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1145), .A2(new_n1164), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n1170));
  XOR2_X1   g745(.A(G299), .B(KEYINPUT57), .Z(new_n1171));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1172), .B1(new_n1135), .B2(new_n803), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1135), .A2(new_n1172), .A3(new_n803), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1032), .A2(new_n1121), .ZN(new_n1177));
  XNOR2_X1  g752(.A(KEYINPUT56), .B(G2072), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1177), .A2(new_n1076), .A3(new_n1120), .A4(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1171), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1175), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1171), .B(new_n1179), .C1(new_n1181), .C2(new_n1173), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1170), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1184));
  AND4_X1   g759(.A1(new_n1038), .A2(new_n1103), .A3(new_n1071), .A4(new_n1068), .ZN(new_n1185));
  INV_X1    g760(.A(G1348), .ZN(new_n1186));
  AOI22_X1  g761(.A1(KEYINPUT123), .A2(new_n1185), .B1(new_n1135), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1188), .B1(new_n1104), .B2(G2067), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1187), .A2(KEYINPUT60), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(KEYINPUT60), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1190), .B1(new_n1191), .B2(new_n623), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1193), .A2(KEYINPUT60), .A3(new_n624), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1104), .ZN(new_n1196));
  XNOR2_X1  g771(.A(KEYINPUT58), .B(G1341), .ZN(new_n1197));
  OAI22_X1  g772(.A1(new_n1122), .A2(G1996), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n632), .A2(KEYINPUT124), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT59), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1179), .B1(new_n1181), .B2(new_n1173), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1171), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1204), .A2(KEYINPUT61), .A3(new_n1182), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1184), .A2(new_n1195), .A3(new_n1201), .A4(new_n1205), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1193), .A2(new_n623), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1182), .B1(new_n1207), .B2(new_n1180), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n1130), .A2(new_n1141), .ZN(new_n1210));
  AND2_X1   g785(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1211));
  XNOR2_X1  g786(.A(G301), .B(KEYINPUT54), .ZN(new_n1212));
  AND2_X1   g787(.A1(new_n1177), .A2(new_n1120), .ZN(new_n1213));
  NOR3_X1   g788(.A1(new_n1131), .A2(new_n1061), .A3(G2078), .ZN(new_n1214));
  AND3_X1   g789(.A1(new_n1071), .A2(new_n1064), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1212), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1216));
  AOI22_X1  g791(.A1(new_n1211), .A2(new_n1216), .B1(new_n1137), .B2(new_n1212), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1210), .A2(new_n1095), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1209), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1058), .B1(new_n1169), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1060), .A2(new_n1076), .ZN(new_n1222));
  NOR2_X1   g797(.A1(new_n1222), .A2(G1996), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n1223), .B(KEYINPUT46), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1044), .A2(new_n1039), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1222), .B1(new_n1225), .B2(new_n766), .ZN(new_n1226));
  NOR2_X1   g801(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  XNOR2_X1  g802(.A(new_n1227), .B(KEYINPUT47), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1035), .A2(new_n1056), .ZN(new_n1229));
  XNOR2_X1  g804(.A(new_n1229), .B(KEYINPUT48), .ZN(new_n1230));
  AOI21_X1  g805(.A(new_n1228), .B1(new_n1054), .B2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g806(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1232));
  INV_X1    g807(.A(KEYINPUT126), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n1232), .A2(new_n1233), .A3(new_n1041), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1234), .A2(new_n1035), .ZN(new_n1235));
  AOI21_X1  g810(.A(new_n1233), .B1(new_n1232), .B2(new_n1041), .ZN(new_n1236));
  OAI21_X1  g811(.A(new_n1231), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g812(.A(new_n1026), .B1(new_n1221), .B2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g813(.A1(new_n1145), .A2(new_n1164), .A3(new_n1168), .ZN(new_n1239));
  AOI21_X1  g814(.A(new_n1218), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1240));
  OAI211_X1 g815(.A(new_n1054), .B(new_n1057), .C1(new_n1239), .C2(new_n1240), .ZN(new_n1241));
  INV_X1    g816(.A(new_n1236), .ZN(new_n1242));
  NAND3_X1  g817(.A1(new_n1242), .A2(new_n1035), .A3(new_n1234), .ZN(new_n1243));
  NAND4_X1  g818(.A1(new_n1241), .A2(KEYINPUT127), .A3(new_n1243), .A4(new_n1231), .ZN(new_n1244));
  NAND2_X1  g819(.A1(new_n1238), .A2(new_n1244), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g820(.A1(new_n930), .A2(KEYINPUT108), .A3(new_n926), .ZN(new_n1247));
  AOI21_X1  g821(.A(KEYINPUT108), .B1(new_n930), .B2(new_n926), .ZN(new_n1248));
  NOR2_X1   g822(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g823(.A(G319), .ZN(new_n1250));
  NOR3_X1   g824(.A1(G227), .A2(G401), .A3(new_n1250), .ZN(new_n1251));
  NAND3_X1  g825(.A1(new_n1022), .A2(new_n712), .A3(new_n1251), .ZN(new_n1252));
  NOR2_X1   g826(.A1(new_n1249), .A2(new_n1252), .ZN(G308));
  OR2_X1    g827(.A1(new_n1249), .A2(new_n1252), .ZN(G225));
endmodule


