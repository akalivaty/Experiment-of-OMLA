//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n189));
  AOI21_X1  g003(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT88), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G214), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT88), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT18), .A2(G131), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT89), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n198), .A2(KEYINPUT89), .A3(new_n200), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n194), .A2(new_n196), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(new_n200), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT78), .B(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G140), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT77), .A3(G125), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT77), .ZN(new_n212));
  INV_X1    g026(.A(G125), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G140), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n210), .A2(G125), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(G140), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n207), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT90), .B1(new_n205), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT89), .B1(new_n198), .B2(new_n200), .ZN(new_n223));
  AOI211_X1 g037(.A(new_n202), .B(new_n199), .C1(new_n191), .C2(new_n197), .ZN(new_n224));
  OAI211_X1 g038(.A(KEYINPUT90), .B(new_n221), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n209), .A2(KEYINPUT16), .A3(new_n211), .A4(new_n214), .ZN(new_n227));
  OR3_X1    g041(.A1(new_n208), .A2(KEYINPUT16), .A3(G140), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(G146), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(G146), .B1(new_n227), .B2(new_n228), .ZN(new_n231));
  OR2_X1    g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n206), .A2(KEYINPUT17), .A3(G131), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n206), .B(G131), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(KEYINPUT17), .ZN(new_n235));
  OAI22_X1  g049(.A1(new_n222), .A2(new_n226), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G113), .B(G122), .ZN(new_n237));
  INV_X1    g051(.A(G104), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n236), .A2(KEYINPUT94), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT94), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n232), .A2(new_n235), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n221), .B1(new_n223), .B2(new_n224), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT90), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n243), .B1(new_n246), .B2(new_n225), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n242), .B1(new_n247), .B2(new_n239), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n236), .A2(new_n240), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n187), .B(new_n241), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G475), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT19), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n217), .A2(new_n218), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n214), .A2(new_n211), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(G140), .B2(new_n208), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n219), .B(new_n253), .C1(new_n255), .C2(new_n252), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT91), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n257), .A3(new_n229), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n258), .A2(new_n234), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n229), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT91), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n246), .A2(new_n225), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT92), .B1(new_n262), .B2(new_n239), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n234), .A3(new_n258), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(new_n222), .B2(new_n226), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT92), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(new_n240), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n247), .A2(new_n239), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n263), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT20), .ZN(new_n270));
  INV_X1    g084(.A(G475), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n187), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n272), .B(KEYINPUT93), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n269), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n270), .B1(new_n269), .B2(new_n273), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n251), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  XOR2_X1   g091(.A(KEYINPUT95), .B(KEYINPUT13), .Z(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(G128), .A3(new_n193), .ZN(new_n279));
  XNOR2_X1  g093(.A(G128), .B(G143), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n279), .B(G134), .C1(new_n278), .C2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G134), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(G116), .B(G122), .ZN(new_n285));
  INV_X1    g099(.A(G107), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n282), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  OR2_X1    g102(.A1(new_n288), .A2(KEYINPUT96), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(KEYINPUT96), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n280), .B(new_n283), .ZN(new_n291));
  INV_X1    g105(.A(G116), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(KEYINPUT14), .A3(G122), .ZN(new_n293));
  INV_X1    g107(.A(new_n285), .ZN(new_n294));
  OAI211_X1 g108(.A(G107), .B(new_n293), .C1(new_n294), .C2(KEYINPUT14), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n291), .B(new_n295), .C1(G107), .C2(new_n294), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n289), .A2(new_n290), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT9), .B(G234), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n298), .B(KEYINPUT82), .ZN(new_n299));
  INV_X1    g113(.A(G953), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT75), .B(G217), .Z(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(KEYINPUT97), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n297), .B(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT98), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n187), .ZN(new_n307));
  INV_X1    g121(.A(G478), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(KEYINPUT15), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n307), .B(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n277), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(G234), .A2(G237), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n313), .A2(G902), .A3(G953), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT21), .B(G898), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g130(.A1(KEYINPUT99), .A2(G952), .ZN(new_n317));
  NOR2_X1   g131(.A1(KEYINPUT99), .A2(G952), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n300), .B(new_n313), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT100), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n312), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G214), .B1(G237), .B2(G902), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G210), .B1(G237), .B2(G902), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT65), .B1(new_n219), .B2(G143), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT65), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n193), .A3(G146), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n219), .A2(G143), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT64), .ZN(new_n333));
  OR3_X1    g147(.A1(new_n193), .A2(KEYINPUT64), .A3(G146), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT0), .ZN(new_n335));
  INV_X1    g149(.A(G128), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n331), .A2(new_n333), .A3(new_n334), .A4(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n337), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n193), .A2(G146), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n332), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n335), .A2(new_n336), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n208), .B1(new_n338), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT87), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n336), .A2(KEYINPUT1), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n331), .A2(new_n333), .A3(new_n334), .A4(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n193), .A2(G146), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT1), .ZN(new_n349));
  OAI21_X1  g163(.A(G128), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n341), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n208), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n344), .A2(KEYINPUT87), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G224), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n355), .B1(new_n356), .B2(G953), .ZN(new_n357));
  OAI211_X1 g171(.A(G224), .B(new_n300), .C1(new_n353), .C2(new_n354), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(G110), .B(G122), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT5), .ZN(new_n362));
  INV_X1    g176(.A(G119), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(G116), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(G116), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n292), .A2(G119), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(G113), .B(new_n364), .C1(new_n367), .C2(new_n362), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n368), .A2(KEYINPUT85), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT3), .B1(new_n238), .B2(G107), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(new_n286), .A3(G104), .ZN(new_n372));
  INV_X1    g186(.A(G101), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n238), .A2(G107), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n370), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n238), .A2(G107), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n286), .A2(G104), .ZN(new_n377));
  OAI21_X1  g191(.A(G101), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n368), .A2(KEYINPUT85), .ZN(new_n381));
  XOR2_X1   g195(.A(KEYINPUT2), .B(G113), .Z(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n365), .A3(new_n366), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n369), .A2(new_n380), .A3(new_n381), .A4(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT2), .B(G113), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n367), .A2(new_n385), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n383), .A2(KEYINPUT68), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT68), .B1(new_n383), .B2(new_n386), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n370), .A2(new_n372), .A3(new_n374), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G101), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT4), .A3(new_n375), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(KEYINPUT4), .B2(new_n391), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n384), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT86), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n361), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n384), .B(KEYINPUT86), .C1(new_n389), .C2(new_n393), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n384), .B(new_n361), .C1(new_n389), .C2(new_n393), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT6), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n396), .A2(KEYINPUT6), .A3(new_n397), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n360), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  XOR2_X1   g217(.A(new_n361), .B(KEYINPUT8), .Z(new_n404));
  NAND2_X1  g218(.A1(new_n368), .A2(new_n383), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n380), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n369), .A2(new_n381), .A3(new_n383), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n406), .B1(new_n407), .B2(new_n380), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT7), .B1(new_n356), .B2(G953), .ZN(new_n409));
  INV_X1    g223(.A(new_n352), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n409), .B1(new_n410), .B2(new_n344), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n399), .A2(new_n408), .A3(new_n411), .ZN(new_n412));
  OR3_X1    g226(.A1(new_n353), .A2(new_n354), .A3(new_n409), .ZN(new_n413));
  AOI21_X1  g227(.A(G902), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n327), .B1(new_n403), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n402), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n396), .A2(new_n397), .B1(KEYINPUT6), .B2(new_n399), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n359), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n326), .A3(new_n414), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n325), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G469), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT11), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(KEYINPUT66), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n283), .A2(G137), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(KEYINPUT66), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT66), .ZN(new_n428));
  INV_X1    g242(.A(G137), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n428), .A2(new_n429), .A3(KEYINPUT11), .A4(G134), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n283), .A2(G137), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n427), .A2(new_n432), .A3(G131), .ZN(new_n433));
  INV_X1    g247(.A(G131), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n429), .A2(G134), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n424), .B2(new_n425), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n428), .A2(KEYINPUT11), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n428), .A2(KEYINPUT11), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n429), .A2(G134), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n434), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  OR2_X1    g255(.A1(new_n433), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n331), .A2(new_n333), .A3(new_n334), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n350), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n379), .B1(new_n444), .B2(new_n347), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n347), .A2(new_n351), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(new_n380), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n442), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT12), .B1(new_n442), .B2(KEYINPUT84), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI221_X1 g264(.A(new_n442), .B1(KEYINPUT84), .B2(KEYINPUT12), .C1(new_n445), .C2(new_n447), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n445), .A2(KEYINPUT10), .ZN(new_n453));
  INV_X1    g267(.A(new_n442), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT70), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n446), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n347), .A2(KEYINPUT70), .A3(new_n351), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n456), .A2(KEYINPUT10), .A3(new_n380), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n338), .A2(new_n343), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n460), .B(new_n392), .C1(KEYINPUT4), .C2(new_n391), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n453), .A2(new_n454), .A3(new_n458), .A4(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G110), .B(G140), .ZN(new_n463));
  INV_X1    g277(.A(G227), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(G953), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n463), .B(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n452), .A2(new_n462), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  OAI22_X1  g283(.A1(new_n393), .A2(new_n459), .B1(new_n445), .B2(KEYINPUT10), .ZN(new_n470));
  INV_X1    g284(.A(new_n457), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n380), .A2(KEYINPUT10), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT70), .B1(new_n347), .B2(new_n351), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n442), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n467), .B1(new_n475), .B2(new_n462), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n422), .B(new_n187), .C1(new_n469), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(G469), .A2(G902), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(new_n462), .A3(new_n467), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n470), .A2(new_n474), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n480), .A2(new_n454), .B1(new_n450), .B2(new_n451), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n466), .B(KEYINPUT83), .Z(new_n482));
  OAI211_X1 g296(.A(G469), .B(new_n479), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n477), .A2(new_n478), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G221), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n299), .B2(new_n187), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n323), .A2(new_n421), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G472), .ZN(new_n490));
  INV_X1    g304(.A(new_n389), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n436), .A2(new_n434), .A3(new_n440), .ZN(new_n492));
  OAI21_X1  g306(.A(G131), .B1(new_n425), .B2(new_n435), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT69), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT69), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n492), .A2(new_n496), .A3(new_n493), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n495), .A2(new_n456), .A3(new_n457), .A4(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n338), .B(new_n343), .C1(new_n433), .C2(new_n441), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(KEYINPUT30), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT67), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n446), .A2(new_n492), .A3(new_n493), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI211_X1 g319(.A(KEYINPUT67), .B(KEYINPUT30), .C1(new_n499), .C2(new_n502), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n491), .B(new_n500), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n188), .A2(G210), .ZN(new_n508));
  XOR2_X1   g322(.A(new_n508), .B(KEYINPUT27), .Z(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT26), .B(G101), .ZN(new_n510));
  XOR2_X1   g324(.A(new_n509), .B(new_n510), .Z(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n498), .A2(new_n389), .A3(new_n499), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n507), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n498), .A2(KEYINPUT28), .A3(new_n389), .A4(new_n499), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n491), .A2(new_n503), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n514), .B1(new_n519), .B2(new_n512), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT29), .ZN(new_n521));
  AOI21_X1  g335(.A(G902), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n516), .B(KEYINPUT73), .Z(new_n523));
  AOI21_X1  g337(.A(new_n389), .B1(new_n498), .B2(new_n499), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n524), .A2(KEYINPUT72), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n513), .B1(new_n524), .B2(KEYINPUT72), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT28), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n523), .A2(KEYINPUT29), .A3(new_n511), .A4(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n490), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(G472), .A2(G902), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n507), .A2(new_n511), .A3(new_n513), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT31), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n507), .A2(KEYINPUT31), .A3(new_n511), .A4(new_n513), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n517), .A2(new_n518), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n511), .B1(new_n536), .B2(new_n516), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT71), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT71), .ZN(new_n540));
  AOI211_X1 g354(.A(new_n540), .B(new_n537), .C1(new_n533), .C2(new_n534), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n530), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT32), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n529), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n535), .A2(new_n538), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n540), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n535), .A2(KEYINPUT71), .A3(new_n538), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n548), .A2(KEYINPUT74), .A3(KEYINPUT32), .A4(new_n530), .ZN(new_n549));
  OAI211_X1 g363(.A(KEYINPUT32), .B(new_n530), .C1(new_n539), .C2(new_n541), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT74), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n544), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n301), .B1(G234), .B2(new_n187), .ZN(new_n554));
  XNOR2_X1  g368(.A(G119), .B(G128), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT76), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT24), .B(G110), .Z(new_n557));
  NAND3_X1  g371(.A1(new_n336), .A2(KEYINPUT23), .A3(G119), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n363), .A2(G128), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n363), .A2(G128), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n558), .B(new_n559), .C1(new_n560), .C2(KEYINPUT23), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n556), .A2(new_n557), .B1(G110), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n230), .B2(new_n231), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT79), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g379(.A(KEYINPUT79), .B(new_n562), .C1(new_n230), .C2(new_n231), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT80), .B(G110), .ZN(new_n568));
  OAI22_X1  g382(.A1(new_n556), .A2(new_n557), .B1(new_n561), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n220), .A3(new_n229), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT22), .B(G137), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n300), .A2(G221), .A3(G234), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n571), .B(new_n572), .Z(new_n573));
  AND3_X1   g387(.A1(new_n567), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n573), .B1(new_n567), .B2(new_n570), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n576), .A2(KEYINPUT25), .A3(new_n187), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT25), .B1(new_n576), .B2(new_n187), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n554), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n554), .A2(G902), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n553), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT81), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT81), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n553), .A2(new_n585), .A3(new_n582), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n489), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(new_n373), .ZN(G3));
  NAND4_X1  g402(.A1(new_n582), .A2(new_n321), .A3(new_n421), .A4(new_n488), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n187), .B1(new_n539), .B2(new_n541), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G472), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n542), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n304), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n297), .B(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n596), .B1(new_n304), .B2(new_n597), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n595), .A2(new_n598), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n308), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n305), .A2(new_n308), .A3(new_n187), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n602), .B1(new_n308), .B2(new_n187), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n276), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n593), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT34), .B(G104), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G6));
  OAI211_X1 g422(.A(new_n310), .B(new_n251), .C1(new_n275), .C2(new_n274), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n593), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT35), .B(G107), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G9));
  AND3_X1   g426(.A1(new_n323), .A2(new_n421), .A3(new_n488), .ZN(new_n613));
  INV_X1    g427(.A(new_n592), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n567), .A2(new_n570), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT36), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n573), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n615), .B(new_n617), .Z(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n580), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n579), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n613), .A2(new_n614), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT37), .B(G110), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G12));
  XNOR2_X1  g437(.A(new_n319), .B(KEYINPUT102), .ZN(new_n624));
  INV_X1    g438(.A(G900), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n314), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n609), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n620), .A2(new_n421), .A3(new_n488), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n553), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G128), .ZN(G30));
  XOR2_X1   g445(.A(new_n627), .B(KEYINPUT39), .Z(new_n632));
  NAND2_X1  g446(.A1(new_n488), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT40), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n416), .A2(new_n420), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT38), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR4_X1   g451(.A1(new_n634), .A2(new_n637), .A3(new_n325), .A4(new_n620), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n549), .A2(new_n552), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n507), .A2(new_n513), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n511), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(G902), .ZN(new_n643));
  OR3_X1    g457(.A1(new_n525), .A2(new_n526), .A3(new_n511), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n490), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n542), .B2(new_n543), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n638), .A2(new_n310), .A3(new_n647), .A4(new_n276), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G143), .ZN(G45));
  INV_X1    g463(.A(new_n627), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n276), .A2(new_n604), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n553), .A2(new_n629), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(KEYINPUT103), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n553), .A2(new_n655), .A3(new_n629), .A4(new_n652), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT104), .B(G146), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G48));
  NAND2_X1  g473(.A1(new_n462), .A2(new_n467), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n476), .B1(new_n452), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(G469), .B1(new_n662), .B2(G902), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n663), .A2(new_n487), .A3(new_n477), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT105), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n663), .A2(new_n487), .A3(new_n477), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n421), .A2(new_n321), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n605), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n553), .A2(new_n582), .A3(new_n669), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  NOR2_X1   g488(.A1(new_n609), .A2(new_n670), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n553), .A2(new_n675), .A3(new_n582), .A4(new_n669), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G116), .ZN(G18));
  NAND2_X1  g491(.A1(new_n421), .A2(new_n664), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n579), .B2(new_n619), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n323), .A2(new_n553), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  AOI21_X1  g495(.A(G902), .B1(new_n546), .B2(new_n547), .ZN(new_n682));
  OAI21_X1  g496(.A(KEYINPUT106), .B1(new_n682), .B2(new_n490), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n590), .A2(new_n684), .A3(G472), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n665), .A2(new_n321), .A3(new_n668), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n276), .A2(new_n310), .A3(new_n421), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n535), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n511), .B1(new_n523), .B2(new_n527), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n530), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n686), .A2(new_n582), .A3(new_n689), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G122), .ZN(G24));
  NOR2_X1   g508(.A1(new_n651), .A2(new_n678), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n686), .A2(new_n620), .A3(new_n692), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G125), .ZN(G27));
  AND3_X1   g511(.A1(new_n416), .A2(new_n420), .A3(new_n324), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n699));
  INV_X1    g513(.A(new_n476), .ZN(new_n700));
  AOI211_X1 g514(.A(G469), .B(G902), .C1(new_n700), .C2(new_n468), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n483), .A2(new_n478), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n699), .B(new_n487), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n699), .B1(new_n484), .B2(new_n487), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n698), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n651), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n544), .A2(new_n550), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n582), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT42), .ZN(new_n710));
  INV_X1    g524(.A(new_n706), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n651), .A2(KEYINPUT42), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n553), .A2(new_n582), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT108), .B(G131), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G33));
  NAND4_X1  g530(.A1(new_n553), .A2(new_n628), .A3(new_n582), .A4(new_n711), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G134), .ZN(G36));
  NAND2_X1  g532(.A1(new_n277), .A2(new_n604), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n719), .B1(KEYINPUT109), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n721), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n592), .A3(new_n620), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n481), .A2(new_n482), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n475), .B2(new_n661), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n729), .A2(KEYINPUT45), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(KEYINPUT45), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(G469), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT46), .B1(new_n732), .B2(new_n478), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n701), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(KEYINPUT46), .A3(new_n478), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n486), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n698), .B(KEYINPUT110), .Z(new_n737));
  AND3_X1   g551(.A1(new_n736), .A2(new_n632), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n726), .A2(new_n727), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G137), .ZN(G39));
  XOR2_X1   g554(.A(new_n736), .B(KEYINPUT47), .Z(new_n741));
  INV_X1    g555(.A(new_n698), .ZN(new_n742));
  OR3_X1    g556(.A1(new_n651), .A2(new_n582), .A3(new_n742), .ZN(new_n743));
  OR3_X1    g557(.A1(new_n741), .A2(new_n553), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G140), .ZN(G42));
  NAND2_X1  g559(.A1(new_n663), .A2(new_n477), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n746), .B(KEYINPUT49), .Z(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(new_n324), .A3(new_n487), .A4(new_n582), .ZN(new_n748));
  NOR4_X1   g562(.A1(new_n647), .A2(new_n748), .A3(new_n636), .A4(new_n719), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT111), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n710), .A2(new_n713), .A3(new_n717), .ZN(new_n751));
  AND4_X1   g565(.A1(new_n672), .A2(new_n693), .A3(new_n676), .A4(new_n680), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n620), .A2(new_n698), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n704), .A2(new_n705), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n651), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n686), .A2(new_n692), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n488), .A2(new_n650), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n312), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n553), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n753), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n751), .A2(new_n752), .A3(new_n761), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n696), .A2(new_n630), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n688), .A2(new_n620), .A3(new_n757), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n647), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n657), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n762), .B1(KEYINPUT52), .B2(new_n766), .ZN(new_n767));
  XOR2_X1   g581(.A(new_n605), .B(KEYINPUT112), .Z(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n593), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT113), .B1(new_n587), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n586), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n585), .B1(new_n553), .B2(new_n582), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n613), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n769), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n621), .A2(new_n610), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n770), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n657), .A2(new_n763), .A3(new_n779), .A4(new_n765), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n767), .A2(new_n778), .A3(KEYINPUT53), .A4(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n766), .A2(KEYINPUT52), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n710), .A2(new_n713), .A3(new_n717), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n672), .A2(new_n693), .A3(new_n676), .A4(new_n680), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n784), .A2(new_n785), .A3(new_n760), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n783), .A2(new_n780), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n770), .A2(new_n776), .A3(new_n777), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n782), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n781), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT115), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n781), .A2(new_n789), .A3(new_n793), .A4(new_n790), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n781), .A2(new_n789), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT54), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n792), .A2(new_n797), .A3(new_n798), .A4(new_n794), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT51), .ZN(new_n804));
  INV_X1    g618(.A(new_n647), .ZN(new_n805));
  INV_X1    g619(.A(new_n319), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n742), .A2(new_n666), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n805), .A2(new_n806), .A3(new_n582), .A4(new_n807), .ZN(new_n808));
  OR3_X1    g622(.A1(new_n808), .A2(new_n276), .A3(new_n604), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n686), .A2(new_n692), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n620), .ZN(new_n811));
  INV_X1    g625(.A(new_n624), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n723), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n807), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n741), .B1(new_n487), .B2(new_n746), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n737), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n810), .A2(new_n582), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n813), .ZN(new_n818));
  OAI221_X1 g632(.A(new_n809), .B1(new_n811), .B2(new_n814), .C1(new_n816), .C2(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n636), .A2(new_n324), .A3(new_n666), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n817), .A2(new_n813), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n821), .B(new_n822), .Z(new_n823));
  OAI21_X1  g637(.A(new_n804), .B1(new_n819), .B2(new_n823), .ZN(new_n824));
  OR3_X1    g638(.A1(new_n819), .A2(new_n804), .A3(new_n823), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n708), .A2(new_n582), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n813), .A2(new_n826), .A3(new_n807), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n827), .B(KEYINPUT48), .Z(new_n828));
  OAI221_X1 g642(.A(new_n300), .B1(new_n803), .B2(KEYINPUT51), .C1(new_n317), .C2(new_n318), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  OAI221_X1 g644(.A(new_n830), .B1(new_n605), .B2(new_n808), .C1(new_n818), .C2(new_n678), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n802), .A2(new_n824), .A3(new_n825), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(G952), .A2(G953), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n750), .B1(new_n833), .B2(new_n834), .ZN(G75));
  XOR2_X1   g649(.A(new_n359), .B(KEYINPUT55), .Z(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n796), .A2(G210), .A3(G902), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n837), .B1(new_n839), .B2(KEYINPUT56), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT56), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(new_n841), .A3(new_n836), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n401), .A2(new_n402), .ZN(new_n844));
  XOR2_X1   g658(.A(new_n844), .B(KEYINPUT118), .Z(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT119), .Z(new_n846));
  NOR2_X1   g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n846), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n840), .B2(new_n842), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n300), .A2(G952), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(G51));
  NAND2_X1  g665(.A1(new_n791), .A2(KEYINPUT120), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n781), .A2(new_n789), .A3(new_n853), .A4(new_n790), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n797), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n796), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n855), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n478), .B(KEYINPUT57), .Z(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n861), .B1(new_n476), .B2(new_n469), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n796), .A2(G902), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n863), .A2(new_n732), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n850), .B1(new_n862), .B2(new_n864), .ZN(G54));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n863), .A2(new_n866), .A3(new_n271), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n867), .A2(new_n269), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n269), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n868), .A2(new_n869), .A3(new_n850), .ZN(G60));
  AND2_X1   g684(.A1(new_n599), .A2(new_n600), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n308), .A2(new_n187), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT59), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n859), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n850), .B1(new_n876), .B2(KEYINPUT122), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n872), .B1(new_n802), .B2(new_n874), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n859), .A2(new_n879), .A3(new_n875), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(G63));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n882));
  NAND2_X1  g696(.A1(G217), .A2(G902), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT60), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n796), .A2(new_n618), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(G952), .B2(new_n300), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n576), .B1(new_n796), .B2(new_n885), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n882), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n887), .B1(new_n888), .B2(KEYINPUT123), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n888), .A2(KEYINPUT123), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n882), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n890), .B2(new_n892), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n889), .B1(new_n894), .B2(new_n895), .ZN(G66));
  INV_X1    g710(.A(new_n315), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n300), .B1(new_n897), .B2(G224), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n778), .A2(new_n752), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n899), .B2(new_n300), .ZN(new_n900));
  INV_X1    g714(.A(G898), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n845), .B1(new_n901), .B2(G953), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n900), .B(new_n902), .ZN(G69));
  OAI21_X1  g717(.A(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n253), .B1(new_n255), .B2(new_n252), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n907), .A2(new_n464), .A3(new_n300), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n744), .A2(new_n739), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n657), .A2(new_n763), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n736), .A2(new_n632), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n688), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n826), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n909), .A2(new_n910), .A3(new_n751), .A4(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(G953), .B1(new_n914), .B2(new_n906), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n768), .A2(new_n609), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n742), .A2(new_n633), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n916), .B(new_n917), .C1(new_n772), .C2(new_n771), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n744), .A2(new_n739), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n910), .A2(new_n648), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n919), .A2(new_n922), .A3(new_n907), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n908), .B1(new_n915), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n464), .B1(new_n907), .B2(KEYINPUT125), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n925), .A2(G900), .ZN(new_n926));
  OAI22_X1  g740(.A1(new_n924), .A2(KEYINPUT125), .B1(new_n300), .B2(new_n926), .ZN(G72));
  NAND2_X1  g741(.A1(G472), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT63), .Z(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(new_n914), .B2(new_n899), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n514), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n931), .B2(new_n930), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n796), .A2(new_n514), .A3(new_n641), .A4(new_n929), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n919), .A2(new_n922), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n929), .B1(new_n935), .B2(new_n899), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n850), .B1(new_n936), .B2(new_n642), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n933), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT127), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n933), .A2(new_n940), .A3(new_n934), .A4(new_n937), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(G57));
endmodule


