//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  OR2_X1    g000(.A1(KEYINPUT66), .A2(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT66), .A2(G119), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(G116), .A3(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n196));
  AND2_X1   g010(.A1(KEYINPUT66), .A2(G119), .ZN(new_n197));
  NOR2_X1   g011(.A1(KEYINPUT66), .A2(G119), .ZN(new_n198));
  INV_X1    g012(.A(G116), .ZN(new_n199));
  NOR3_X1   g013(.A1(new_n197), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n196), .B1(new_n200), .B2(new_n191), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n189), .A2(KEYINPUT67), .A3(new_n192), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n195), .B1(new_n203), .B2(new_n194), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G104), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G101), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n206), .A2(new_n209), .A3(new_n213), .A4(new_n210), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(KEYINPUT4), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT4), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n211), .A2(new_n216), .A3(G101), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT82), .B1(new_n204), .B2(new_n218), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n189), .A2(KEYINPUT67), .A3(new_n192), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT67), .B1(new_n189), .B2(new_n192), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n194), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n195), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n215), .A2(new_n217), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT82), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n219), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n201), .A2(new_n202), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n189), .A2(new_n229), .ZN(new_n231));
  INV_X1    g045(.A(G113), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n195), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n205), .A2(G107), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n208), .A2(G104), .ZN(new_n236));
  OAI21_X1  g050(.A(G101), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n214), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n234), .A2(KEYINPUT84), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n230), .A2(new_n233), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(new_n223), .A3(new_n239), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT84), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n228), .A2(new_n240), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G110), .B(G122), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT85), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n228), .A2(new_n246), .A3(new_n240), .A4(new_n244), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n248), .A2(new_n249), .A3(KEYINPUT6), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(KEYINPUT6), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n234), .A2(KEYINPUT84), .A3(new_n239), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT84), .B1(new_n234), .B2(new_n239), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n246), .B1(new_n255), .B2(new_n228), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n245), .A2(new_n258), .A3(new_n247), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT85), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n251), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G143), .ZN(new_n263));
  INV_X1    g077(.A(G143), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G146), .ZN(new_n265));
  OR2_X1    g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n263), .A2(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n263), .A2(new_n265), .A3(new_n267), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G125), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT1), .B1(new_n264), .B2(G146), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G128), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n263), .A2(new_n265), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT1), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n263), .A2(new_n265), .A3(new_n277), .A4(G128), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G125), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n272), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G953), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G224), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n282), .A2(G224), .A3(new_n284), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n261), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G210), .B1(G237), .B2(G902), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT7), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n286), .A2(new_n287), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n283), .A2(new_n292), .A3(new_n285), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n246), .B(KEYINPUT8), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n189), .A2(KEYINPUT5), .A3(new_n192), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n195), .B1(new_n233), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n297), .B1(new_n299), .B2(new_n238), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(new_n238), .B2(new_n234), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(G902), .B1(new_n302), .B2(new_n250), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n290), .A2(new_n291), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n291), .ZN(new_n305));
  OAI211_X1 g119(.A(KEYINPUT85), .B(new_n259), .C1(new_n252), .C2(new_n256), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n288), .B1(new_n306), .B2(new_n251), .ZN(new_n307));
  INV_X1    g121(.A(new_n303), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n304), .A2(new_n309), .A3(KEYINPUT86), .ZN(new_n310));
  OAI21_X1  g124(.A(G214), .B1(G237), .B2(G902), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT86), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n290), .A2(new_n312), .A3(new_n291), .A4(new_n303), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(G475), .A2(G902), .ZN(new_n315));
  XNOR2_X1  g129(.A(G113), .B(G122), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(new_n205), .ZN(new_n317));
  NOR2_X1   g131(.A1(KEYINPUT68), .A2(G953), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G237), .ZN(new_n320));
  NAND2_X1  g134(.A1(KEYINPUT68), .A2(G953), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n319), .A2(G214), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n264), .ZN(new_n323));
  AND2_X1   g137(.A1(KEYINPUT68), .A2(G953), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(new_n318), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n325), .A2(G143), .A3(G214), .A4(new_n320), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(KEYINPUT18), .A3(G131), .ZN(new_n328));
  NAND2_X1  g142(.A1(KEYINPUT18), .A2(G131), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n323), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n280), .A2(G140), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G146), .ZN(new_n335));
  XNOR2_X1  g149(.A(G125), .B(G140), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n262), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n337), .A3(KEYINPUT87), .ZN(new_n338));
  OR3_X1    g152(.A1(new_n336), .A2(KEYINPUT87), .A3(new_n262), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n328), .A2(new_n330), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n327), .A2(G131), .ZN(new_n341));
  INV_X1    g155(.A(G131), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n342), .B1(new_n323), .B2(new_n326), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n341), .A2(KEYINPUT17), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(KEYINPUT17), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n336), .A2(KEYINPUT16), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n332), .A2(KEYINPUT16), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(G146), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(G146), .B1(new_n346), .B2(new_n347), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n317), .B(new_n340), .C1(new_n344), .C2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT19), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n334), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n336), .A2(KEYINPUT19), .ZN(new_n357));
  AOI21_X1  g171(.A(G146), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n349), .B1(KEYINPUT88), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n334), .A2(new_n355), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n336), .A2(KEYINPUT19), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n262), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT88), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n359), .B(new_n364), .C1(new_n343), .C2(new_n341), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n317), .B1(new_n365), .B2(new_n340), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n315), .B1(new_n354), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT89), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT20), .ZN(new_n369));
  INV_X1    g183(.A(new_n315), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n341), .A2(new_n343), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n358), .A2(KEYINPUT88), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n364), .A2(new_n372), .A3(new_n348), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n340), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n317), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n370), .B1(new_n376), .B2(new_n353), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT20), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT89), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n378), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n369), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n340), .B1(new_n344), .B2(new_n352), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n375), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT90), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n383), .A2(new_n384), .A3(new_n353), .ZN(new_n385));
  INV_X1    g199(.A(G902), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(new_n383), .B2(new_n384), .ZN(new_n387));
  OAI21_X1  g201(.A(G475), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n381), .A2(new_n388), .ZN(new_n389));
  AOI211_X1 g203(.A(new_n386), .B(new_n325), .C1(G234), .C2(G237), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT21), .B(G898), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G952), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n393), .A2(KEYINPUT94), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(KEYINPUT94), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n284), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(G234), .B2(G237), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  XOR2_X1   g213(.A(new_n399), .B(KEYINPUT95), .Z(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT9), .B(G234), .ZN(new_n402));
  INV_X1    g216(.A(G217), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n402), .A2(new_n403), .A3(G953), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT91), .ZN(new_n406));
  INV_X1    g220(.A(G122), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G116), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n199), .A2(G122), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(G107), .ZN(new_n411));
  XNOR2_X1  g225(.A(G116), .B(G122), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(new_n208), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n406), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G128), .B(G143), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n264), .A2(G128), .ZN(new_n417));
  OAI21_X1  g231(.A(G134), .B1(new_n417), .B2(KEYINPUT13), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n415), .B(G134), .C1(KEYINPUT13), .C2(new_n417), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n410), .A2(G107), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n412), .A2(new_n208), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT91), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n414), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT92), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n199), .A2(KEYINPUT14), .A3(G122), .ZN(new_n427));
  OAI211_X1 g241(.A(G107), .B(new_n427), .C1(new_n410), .C2(KEYINPUT14), .ZN(new_n428));
  INV_X1    g242(.A(G134), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n416), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n415), .A2(G134), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n428), .A2(new_n430), .A3(new_n423), .A4(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n425), .A2(new_n426), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n426), .B1(new_n425), .B2(new_n432), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n405), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n425), .A2(new_n432), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT92), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n425), .A2(new_n426), .A3(new_n432), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n404), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(KEYINPUT93), .A3(new_n386), .ZN(new_n441));
  INV_X1    g255(.A(G478), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(KEYINPUT15), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n441), .B(new_n443), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n389), .A2(new_n401), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G221), .B1(new_n402), .B2(G902), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT10), .ZN(new_n448));
  INV_X1    g262(.A(new_n278), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT79), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n273), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(KEYINPUT79), .B(KEYINPUT1), .C1(new_n264), .C2(G146), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(G128), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n449), .B1(new_n453), .B2(new_n275), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT80), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n454), .A2(new_n455), .A3(new_n238), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n452), .A2(G128), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT79), .B1(new_n263), .B2(KEYINPUT1), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n275), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n278), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT80), .B1(new_n460), .B2(new_n239), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n448), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n448), .B1(new_n276), .B2(new_n278), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n239), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n218), .B2(new_n270), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT64), .B1(new_n429), .B2(G137), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n467), .A2(KEYINPUT11), .B1(new_n429), .B2(G137), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT11), .ZN(new_n469));
  OAI211_X1 g283(.A(KEYINPUT64), .B(new_n469), .C1(new_n429), .C2(G137), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n342), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n342), .B1(new_n468), .B2(new_n470), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n462), .A2(new_n466), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n474), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n455), .B1(new_n454), .B2(new_n238), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n460), .A2(KEYINPUT80), .A3(new_n239), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT10), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n476), .B1(new_n479), .B2(new_n465), .ZN(new_n480));
  XOR2_X1   g294(.A(G110), .B(G140), .Z(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT78), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n325), .A2(G227), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n482), .B(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n475), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n479), .A2(new_n476), .A3(new_n465), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n456), .A2(new_n461), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n239), .A2(new_n279), .ZN(new_n488));
  OAI211_X1 g302(.A(KEYINPUT12), .B(new_n476), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT12), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n488), .B1(new_n477), .B2(new_n478), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n490), .B1(new_n491), .B2(new_n474), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n486), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(G469), .B(new_n485), .C1(new_n493), .C2(new_n484), .ZN(new_n494));
  INV_X1    g308(.A(G469), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(new_n386), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT81), .ZN(new_n499));
  INV_X1    g313(.A(new_n484), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n499), .B1(new_n486), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n489), .A2(new_n492), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n475), .A2(KEYINPUT81), .A3(new_n484), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n480), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n500), .B1(new_n505), .B2(new_n486), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n495), .A3(new_n386), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n447), .B1(new_n498), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n445), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n314), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n403), .B1(G234), .B2(new_n386), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  XOR2_X1   g327(.A(KEYINPUT24), .B(G110), .Z(new_n514));
  NAND3_X1  g328(.A1(new_n187), .A2(G128), .A3(new_n188), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT73), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n190), .A2(G128), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n516), .B1(new_n515), .B2(new_n518), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n514), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT74), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(KEYINPUT74), .B(new_n514), .C1(new_n519), .C2(new_n520), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n351), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n515), .A2(KEYINPUT23), .ZN(new_n527));
  INV_X1    g341(.A(G128), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n528), .B1(new_n197), .B2(new_n198), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT75), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT75), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n531), .B(new_n528), .C1(new_n197), .C2(new_n198), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n527), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n517), .A2(KEYINPUT23), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT76), .B1(new_n535), .B2(G110), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT76), .ZN(new_n537));
  INV_X1    g351(.A(G110), .ZN(new_n538));
  AOI211_X1 g352(.A(new_n537), .B(new_n538), .C1(new_n533), .C2(new_n534), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n525), .B(new_n526), .C1(new_n536), .C2(new_n539), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n348), .A2(new_n337), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT77), .ZN(new_n542));
  AOI22_X1  g356(.A1(KEYINPUT23), .A2(new_n515), .B1(new_n529), .B2(KEYINPUT75), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n543), .A2(new_n532), .B1(KEYINPUT23), .B2(new_n517), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n542), .B1(new_n544), .B2(new_n538), .ZN(new_n545));
  OR3_X1    g359(.A1(new_n519), .A2(new_n520), .A3(new_n514), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n533), .A2(new_n542), .A3(new_n538), .A4(new_n534), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n541), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n325), .A2(G221), .A3(G234), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT22), .B(G137), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n540), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n552), .B1(new_n540), .B2(new_n549), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(KEYINPUT25), .A3(new_n386), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n540), .A2(new_n549), .ZN(new_n557));
  INV_X1    g371(.A(new_n552), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n540), .A2(new_n549), .A3(new_n552), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n386), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT25), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n513), .B1(new_n556), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n512), .A2(G902), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n555), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n467), .A2(KEYINPUT11), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n429), .A2(G137), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n470), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G131), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n270), .B1(new_n572), .B2(new_n471), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT65), .B1(new_n429), .B2(G137), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n570), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n429), .A2(KEYINPUT65), .A3(G137), .ZN(new_n576));
  OAI21_X1  g390(.A(G131), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n279), .A2(new_n471), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n224), .B1(new_n573), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n271), .B1(new_n472), .B2(new_n473), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n279), .A2(new_n471), .A3(new_n577), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n204), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT28), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT28), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT69), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n582), .A2(KEYINPUT69), .A3(new_n585), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n325), .A2(G210), .A3(new_n320), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT27), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT26), .B(G101), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n582), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT30), .B1(new_n578), .B2(new_n573), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT30), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n580), .A2(new_n599), .A3(new_n581), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n597), .B1(new_n601), .B2(new_n224), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT31), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n603), .A3(new_n594), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n578), .A2(new_n573), .A3(KEYINPUT30), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n599), .B1(new_n580), .B2(new_n581), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n224), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(new_n594), .A3(new_n582), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT31), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n596), .A2(new_n604), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(G472), .A2(G902), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT70), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT71), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT32), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT71), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n610), .A2(new_n617), .A3(new_n613), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n584), .A2(new_n588), .A3(new_n594), .A4(new_n589), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(KEYINPUT72), .B2(KEYINPUT29), .ZN(new_n621));
  AOI22_X1  g435(.A1(KEYINPUT28), .A2(new_n583), .B1(new_n586), .B2(new_n587), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT72), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n622), .A2(new_n623), .A3(new_n594), .A4(new_n589), .ZN(new_n624));
  INV_X1    g438(.A(new_n602), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n595), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n621), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n590), .A2(new_n595), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n628), .B2(KEYINPUT29), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n590), .A2(new_n595), .B1(new_n608), .B2(KEYINPUT31), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n612), .B1(new_n631), .B2(new_n604), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n630), .A2(G472), .B1(new_n632), .B2(KEYINPUT32), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n568), .B1(new_n619), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n511), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT96), .B(G101), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G3));
  INV_X1    g451(.A(KEYINPUT33), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n440), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n435), .A2(new_n439), .A3(KEYINPUT33), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n442), .A2(G902), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n440), .A2(new_n386), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT97), .B(G478), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n642), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n643), .B1(new_n642), .B2(new_n646), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n389), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT99), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n642), .A2(new_n646), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT98), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n653), .A2(new_n647), .B1(new_n381), .B2(new_n388), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n311), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n304), .B2(new_n309), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n657), .A2(new_n400), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n615), .A2(new_n618), .ZN(new_n661));
  INV_X1    g475(.A(G472), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n610), .B2(new_n386), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n567), .A3(new_n509), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT34), .B(G104), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n369), .A2(new_n379), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n669), .B1(new_n369), .B2(new_n379), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n380), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n444), .A2(new_n388), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n659), .A2(new_n674), .A3(new_n400), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n665), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT35), .B(G107), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  AND2_X1   g492(.A1(new_n615), .A2(new_n618), .ZN(new_n679));
  INV_X1    g493(.A(new_n663), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT25), .B1(new_n555), .B2(new_n386), .ZN(new_n681));
  NOR4_X1   g495(.A1(new_n553), .A2(new_n554), .A3(new_n562), .A4(G902), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n512), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n558), .A2(KEYINPUT36), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n557), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n565), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n679), .A2(new_n680), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT101), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n511), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT37), .B(G110), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G12));
  NAND2_X1  g506(.A1(new_n556), .A2(new_n563), .ZN(new_n693));
  AOI22_X1  g507(.A1(new_n693), .A2(new_n512), .B1(new_n565), .B2(new_n685), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n619), .B2(new_n633), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n509), .A3(new_n659), .ZN(new_n696));
  INV_X1    g510(.A(G900), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n390), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n398), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n672), .A2(new_n673), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n672), .A2(new_n673), .A3(KEYINPUT102), .A4(new_n699), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n696), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n528), .ZN(G30));
  NAND2_X1  g520(.A1(new_n310), .A2(new_n313), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT38), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n699), .B(KEYINPUT39), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n509), .A2(new_n709), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n625), .A2(new_n594), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n583), .A2(new_n594), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(G902), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n662), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n716), .B1(new_n632), .B2(KEYINPUT32), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n619), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n389), .A2(new_n444), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n687), .A2(new_n719), .A3(new_n658), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n711), .A2(new_n712), .A3(new_n718), .A4(new_n720), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n708), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT103), .B(G143), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G45));
  NAND2_X1  g538(.A1(new_n654), .A2(new_n699), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n695), .A2(new_n509), .A3(new_n726), .A4(new_n659), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G146), .ZN(G48));
  NAND2_X1  g542(.A1(new_n619), .A2(new_n633), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n507), .A2(new_n386), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G469), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n731), .A2(new_n446), .A3(new_n508), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n729), .A2(new_n567), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n660), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT41), .B(G113), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  NOR2_X1   g550(.A1(new_n675), .A2(new_n733), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT104), .B(G116), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G18));
  NAND4_X1  g553(.A1(new_n695), .A2(new_n659), .A3(new_n445), .A4(new_n732), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  AOI21_X1  g555(.A(G902), .B1(new_n631), .B2(new_n604), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n614), .B1(new_n742), .B2(new_n662), .ZN(new_n743));
  NOR4_X1   g557(.A1(new_n743), .A2(new_n564), .A3(new_n566), .A4(new_n401), .ZN(new_n744));
  INV_X1    g558(.A(new_n719), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(new_n659), .A3(new_n745), .A4(new_n732), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  OAI21_X1  g561(.A(KEYINPUT105), .B1(new_n694), .B2(new_n743), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n663), .A2(new_n632), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n687), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(new_n659), .A3(new_n726), .A4(new_n732), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G125), .ZN(G27));
  AOI21_X1  g568(.A(new_n658), .B1(new_n310), .B2(new_n313), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n756));
  AOI211_X1 g570(.A(G469), .B(G902), .C1(new_n504), .C2(new_n506), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n494), .A2(new_n497), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n498), .A2(new_n508), .A3(KEYINPUT106), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n759), .A2(new_n446), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT107), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n759), .A2(new_n760), .A3(new_n446), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n755), .A2(new_n762), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(new_n767), .A3(new_n634), .A4(new_n726), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n755), .A2(new_n762), .A3(new_n634), .A4(new_n765), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT108), .B1(new_n769), .B2(new_n725), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT42), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n614), .A2(new_n616), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n568), .B1(new_n633), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n766), .A2(KEYINPUT42), .A3(new_n726), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G131), .ZN(G33));
  NAND2_X1  g591(.A1(new_n704), .A2(KEYINPUT109), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n702), .A2(new_n779), .A3(new_n703), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n766), .A2(new_n634), .A3(new_n778), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G134), .ZN(G36));
  OAI21_X1  g596(.A(new_n485), .B1(new_n493), .B2(new_n484), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n495), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n785), .B1(new_n784), .B2(new_n783), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT110), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n497), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(KEYINPUT46), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n508), .B1(new_n791), .B2(KEYINPUT46), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n446), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n709), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n389), .B1(new_n647), .B2(new_n653), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT43), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n664), .A2(new_n694), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT44), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n755), .B1(new_n800), .B2(new_n801), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(KEYINPUT111), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(KEYINPUT111), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n796), .B(new_n802), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G137), .ZN(G39));
  INV_X1    g621(.A(new_n755), .ZN(new_n808));
  OR4_X1    g622(.A1(new_n729), .A2(new_n808), .A3(new_n567), .A4(new_n725), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT47), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n794), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g625(.A(KEYINPUT47), .B(new_n446), .C1(new_n792), .C2(new_n793), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n809), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(new_n331), .ZN(G42));
  AND2_X1   g628(.A1(new_n731), .A2(new_n508), .ZN(new_n815));
  XOR2_X1   g629(.A(new_n815), .B(KEYINPUT49), .Z(new_n816));
  INV_X1    g630(.A(new_n797), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n816), .A2(new_n718), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n567), .A2(new_n311), .A3(new_n446), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n819), .B(KEYINPUT112), .Z(new_n820));
  NAND3_X1  g634(.A1(new_n818), .A2(new_n708), .A3(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n683), .A2(new_n686), .A3(new_n699), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n619), .B2(new_n717), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(new_n761), .A3(new_n659), .A4(new_n745), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI211_X1 g641(.A(new_n658), .B(new_n719), .C1(new_n304), .C2(new_n309), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(KEYINPUT113), .A3(new_n761), .A4(new_n824), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n753), .B(new_n727), .C1(new_n704), .C2(new_n696), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n822), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT115), .ZN(new_n833));
  INV_X1    g647(.A(new_n831), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n827), .A2(new_n829), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(KEYINPUT52), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n837), .B(new_n822), .C1(new_n830), .C2(new_n831), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n833), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n740), .B(new_n746), .C1(new_n660), .C2(new_n733), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n444), .A2(new_n381), .A3(new_n388), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n401), .B1(new_n650), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n664), .A3(new_n567), .A4(new_n509), .ZN(new_n843));
  OAI22_X1  g657(.A1(new_n843), .A2(new_n314), .B1(new_n675), .B2(new_n733), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n725), .B1(new_n748), .B2(new_n751), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(new_n755), .A3(new_n762), .A4(new_n765), .ZN(new_n847));
  INV_X1    g661(.A(new_n444), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n388), .A2(new_n672), .A3(new_n848), .A4(new_n699), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n755), .A2(new_n509), .A3(new_n695), .A4(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n511), .B1(new_n689), .B2(new_n634), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n845), .A2(new_n781), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n853), .B1(new_n772), .B2(new_n775), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n839), .A2(new_n854), .A3(KEYINPUT53), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n781), .A2(new_n845), .A3(new_n852), .A4(new_n851), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n857), .B1(new_n830), .B2(new_n831), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n836), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n856), .A2(new_n859), .A3(new_n776), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n855), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n798), .A2(new_n397), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n755), .A2(new_n732), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n752), .ZN(new_n869));
  OR4_X1    g683(.A1(new_n568), .A2(new_n867), .A3(new_n398), .A4(new_n718), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n653), .A2(new_n381), .A3(new_n388), .A4(new_n647), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n567), .A2(new_n749), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n866), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n708), .A3(new_n658), .A4(new_n732), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT50), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n876), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n872), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n811), .A2(new_n812), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n815), .A2(new_n447), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n755), .B(new_n874), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT51), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n879), .A2(new_n882), .A3(KEYINPUT51), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n868), .A2(new_n774), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT48), .Z(new_n888));
  AOI21_X1  g702(.A(new_n870), .B1(new_n651), .B2(new_n656), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n874), .A2(new_n659), .A3(new_n732), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n396), .B(KEYINPUT117), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n888), .A2(new_n889), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n885), .A2(new_n886), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n854), .A2(KEYINPUT53), .A3(new_n859), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(KEYINPUT116), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n839), .A2(new_n854), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT116), .B1(new_n897), .B2(new_n861), .ZN(new_n898));
  INV_X1    g712(.A(new_n894), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI211_X1 g714(.A(new_n865), .B(new_n893), .C1(new_n900), .C2(KEYINPUT54), .ZN(new_n901));
  NOR2_X1   g715(.A1(G952), .A2(G953), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n821), .B1(new_n901), .B2(new_n902), .ZN(G75));
  NOR2_X1   g717(.A1(new_n325), .A2(G952), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n386), .B1(new_n855), .B2(new_n862), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT56), .B1(new_n906), .B2(G210), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n261), .B(new_n289), .ZN(new_n908));
  XNOR2_X1  g722(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n908), .B(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n905), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(G210), .ZN(new_n912));
  AOI211_X1 g726(.A(new_n912), .B(new_n386), .C1(new_n855), .C2(new_n862), .ZN(new_n913));
  INV_X1    g727(.A(new_n910), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(KEYINPUT56), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT119), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n907), .A2(new_n910), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n914), .B1(new_n913), .B2(KEYINPUT56), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT119), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .A4(new_n905), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n916), .A2(new_n920), .ZN(G51));
  NAND2_X1  g735(.A1(new_n855), .A2(new_n862), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n923), .A2(KEYINPUT120), .A3(new_n864), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n925), .A3(KEYINPUT54), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n496), .B(KEYINPUT57), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n507), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n788), .A2(new_n789), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n906), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n904), .B1(new_n929), .B2(new_n931), .ZN(G54));
  AND3_X1   g746(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n376), .A2(new_n353), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n905), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n934), .B2(new_n933), .ZN(G60));
  INV_X1    g750(.A(new_n639), .ZN(new_n937));
  INV_X1    g751(.A(new_n640), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n838), .A2(new_n836), .ZN(new_n940));
  INV_X1    g754(.A(new_n705), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n835), .A2(new_n941), .A3(new_n727), .A4(new_n753), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n837), .B1(new_n942), .B2(new_n822), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n856), .A2(new_n776), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n861), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT116), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n895), .B1(new_n948), .B2(new_n894), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n864), .B1(new_n949), .B2(new_n863), .ZN(new_n950));
  NAND2_X1  g764(.A1(G478), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT59), .Z(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n939), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n937), .A2(new_n938), .A3(new_n952), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n924), .A2(new_n926), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n905), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n954), .A2(new_n957), .ZN(G63));
  NAND2_X1  g772(.A1(G217), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT60), .Z(new_n960));
  NAND2_X1  g774(.A1(new_n922), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n553), .B2(new_n554), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n922), .A2(new_n685), .A3(new_n960), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n905), .A3(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n962), .A2(KEYINPUT61), .A3(new_n905), .A4(new_n963), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(G66));
  NAND2_X1  g782(.A1(new_n845), .A2(new_n852), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n325), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT121), .Z(new_n971));
  INV_X1    g785(.A(G224), .ZN(new_n972));
  OAI21_X1  g786(.A(G953), .B1(new_n391), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT122), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n306), .B(new_n251), .C1(G898), .C2(new_n325), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  NOR2_X1   g791(.A1(new_n360), .A2(new_n361), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n601), .B(new_n978), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT123), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n722), .A2(new_n834), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n981), .A2(KEYINPUT62), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT124), .ZN(new_n983));
  INV_X1    g797(.A(new_n634), .ZN(new_n984));
  AOI211_X1 g798(.A(new_n710), .B(new_n984), .C1(new_n650), .C2(new_n841), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n755), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n806), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n813), .B1(KEYINPUT62), .B2(new_n981), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n983), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n325), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n980), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n979), .B1(G900), .B2(new_n991), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n796), .A2(new_n828), .A3(new_n774), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n781), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n995), .A2(new_n813), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT125), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n806), .A2(new_n997), .A3(new_n834), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n997), .B1(new_n806), .B2(new_n834), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n776), .B(new_n996), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n993), .B1(new_n1000), .B2(new_n991), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n992), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n325), .B1(G227), .B2(G900), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1003), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n992), .A2(new_n1001), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1004), .A2(new_n1006), .ZN(G72));
  XNOR2_X1  g821(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1008));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1010), .B1(new_n989), .B2(new_n969), .ZN(new_n1011));
  INV_X1    g825(.A(new_n713), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n904), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1010), .B1(new_n1000), .B2(new_n969), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1014), .A2(new_n595), .A3(new_n602), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n626), .B(KEYINPUT127), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n608), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n900), .A2(new_n1010), .A3(new_n1017), .ZN(new_n1018));
  AND3_X1   g832(.A1(new_n1013), .A2(new_n1015), .A3(new_n1018), .ZN(G57));
endmodule


