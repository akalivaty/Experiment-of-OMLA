//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT24), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G183gat), .ZN(new_n211));
  INV_X1    g010(.A(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT24), .A3(new_n207), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n205), .A2(new_n210), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT25), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT64), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n215), .A2(new_n216), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n216), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n206), .A2(new_n203), .A3(KEYINPUT26), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n203), .A2(KEYINPUT26), .ZN(new_n225));
  NOR3_X1   g024(.A1(new_n224), .A2(new_n225), .A3(new_n208), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT27), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT27), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G183gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n229), .A3(new_n212), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT28), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(KEYINPUT65), .A3(new_n231), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n228), .A2(G183gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n211), .A2(KEYINPUT27), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT66), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n227), .A2(new_n229), .A3(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n231), .A2(G190gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT67), .B1(new_n236), .B2(new_n243), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n230), .A2(KEYINPUT65), .A3(new_n231), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT65), .B1(new_n230), .B2(new_n231), .ZN(new_n246));
  OAI211_X1 g045(.A(KEYINPUT67), .B(new_n243), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n226), .B1(new_n244), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT68), .ZN(new_n250));
  INV_X1    g049(.A(new_n226), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n243), .B1(new_n245), .B2(new_n246), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n251), .B1(new_n254), .B2(new_n247), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n223), .B1(new_n250), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n202), .B1(new_n258), .B2(KEYINPUT29), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n249), .A2(KEYINPUT71), .A3(new_n217), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n261));
  INV_X1    g060(.A(new_n217), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n255), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n264));
  INV_X1    g063(.A(new_n202), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n260), .A2(new_n263), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n260), .A2(new_n263), .A3(new_n265), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT72), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n259), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(G197gat), .A2(G204gat), .ZN(new_n270));
  AND2_X1   g069(.A1(G197gat), .A2(G204gat), .ZN(new_n271));
  AND2_X1   g070(.A1(G211gat), .A2(G218gat), .ZN(new_n272));
  OAI22_X1  g071(.A1(new_n270), .A2(new_n271), .B1(new_n272), .B2(KEYINPUT22), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n273), .A2(KEYINPUT70), .ZN(new_n274));
  NOR2_X1   g073(.A1(G211gat), .A2(G218gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n274), .A2(new_n277), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n269), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT73), .ZN(new_n282));
  INV_X1    g081(.A(new_n222), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n220), .B1(new_n219), .B2(new_n221), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n254), .A2(new_n247), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n256), .B1(new_n286), .B2(new_n226), .ZN(new_n287));
  AOI211_X1 g086(.A(KEYINPUT68), .B(new_n251), .C1(new_n254), .C2(new_n247), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n285), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n260), .A2(new_n263), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n265), .A2(KEYINPUT29), .ZN(new_n291));
  OAI22_X1  g090(.A1(new_n202), .A2(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n280), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n269), .A2(new_n295), .A3(new_n280), .ZN(new_n296));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n297), .B(new_n298), .Z(new_n299));
  NAND4_X1  g098(.A1(new_n282), .A2(new_n294), .A3(new_n296), .A4(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT30), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n296), .A2(new_n294), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n303), .A2(KEYINPUT30), .A3(new_n282), .A4(new_n299), .ZN(new_n304));
  INV_X1    g103(.A(new_n299), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n296), .A2(new_n294), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n295), .B1(new_n269), .B2(new_n280), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n302), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G120gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G113gat), .ZN(new_n312));
  INV_X1    g111(.A(G113gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G120gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n318));
  INV_X1    g117(.A(G127gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G134gat), .ZN(new_n322));
  INV_X1    g121(.A(G134gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n318), .A2(new_n323), .A3(new_n320), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n289), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G227gat), .ZN(new_n327));
  INV_X1    g126(.A(G233gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n322), .A2(new_n324), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n285), .B(new_n330), .C1(new_n287), .C2(new_n288), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n326), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT33), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(G15gat), .B(G43gat), .Z(new_n335));
  XNOR2_X1  g134(.A(G71gat), .B(G99gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n326), .A2(new_n331), .ZN(new_n339));
  INV_X1    g138(.A(new_n329), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT34), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT34), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(new_n343), .A3(new_n340), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n338), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n332), .A2(KEYINPUT32), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n337), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(new_n332), .B2(new_n333), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n343), .B1(new_n339), .B2(new_n340), .ZN(new_n350));
  AOI211_X1 g149(.A(KEYINPUT34), .B(new_n329), .C1(new_n326), .C2(new_n331), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n345), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n354));
  XNOR2_X1  g153(.A(G141gat), .B(G148gat), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT2), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(G155gat), .B2(G162gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT74), .ZN(new_n358));
  AND2_X1   g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359));
  OAI22_X1  g158(.A1(new_n355), .A2(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n360), .A2(new_n362), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(KEYINPUT29), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT78), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(new_n368), .B2(KEYINPUT29), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n280), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G228gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n280), .B2(KEYINPUT29), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n377), .B1(new_n363), .B2(new_n364), .ZN(new_n378));
  OR2_X1    g177(.A1(new_n360), .A2(new_n362), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n360), .A2(new_n362), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(KEYINPUT75), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n374), .B1(new_n376), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n373), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G22gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n379), .A2(new_n380), .ZN(new_n386));
  OR2_X1    g185(.A1(new_n277), .A2(new_n273), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT29), .B1(new_n277), .B2(new_n273), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n367), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT77), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  OR3_X1    g189(.A1(new_n386), .A2(new_n389), .A3(KEYINPUT77), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n390), .B(new_n391), .C1(new_n369), .C2(new_n293), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n374), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n384), .A2(new_n385), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n385), .B1(new_n384), .B2(new_n393), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n354), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n396), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n398), .A2(KEYINPUT79), .A3(new_n394), .ZN(new_n399));
  XNOR2_X1  g198(.A(G78gat), .B(G106gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT31), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(G50gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n397), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n354), .B(new_n402), .C1(new_n395), .C2(new_n396), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n347), .B1(new_n345), .B2(new_n352), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n353), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n325), .A2(KEYINPUT4), .A3(new_n386), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT4), .B1(new_n325), .B2(new_n386), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n375), .B1(new_n378), .B2(new_n381), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n322), .B(new_n324), .C1(new_n365), .C2(new_n367), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G225gat), .A2(G233gat), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n411), .A2(new_n415), .A3(KEYINPUT5), .A4(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n416), .ZN(new_n418));
  NOR4_X1   g217(.A1(new_n414), .A2(new_n409), .A3(new_n410), .A4(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT5), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n330), .A2(new_n382), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n421), .B1(new_n365), .B2(new_n330), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n420), .B1(new_n422), .B2(new_n418), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n417), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G1gat), .B(G29gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT0), .ZN(new_n426));
  XNOR2_X1  g225(.A(G57gat), .B(G85gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  NAND2_X1  g227(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430));
  INV_X1    g229(.A(new_n428), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n431), .B(new_n417), .C1(new_n419), .C2(new_n423), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  OR3_X1    g232(.A1(new_n424), .A2(new_n430), .A3(new_n428), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n310), .A2(new_n408), .A3(KEYINPUT35), .A4(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT35), .ZN(new_n438));
  INV_X1    g237(.A(new_n406), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n345), .A2(new_n347), .A3(new_n352), .ZN(new_n440));
  INV_X1    g239(.A(new_n352), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n346), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n302), .A2(new_n436), .A3(new_n304), .A4(new_n308), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n438), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n437), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n411), .A2(new_n415), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n418), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n450), .B(KEYINPUT39), .C1(new_n418), .C2(new_n422), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n451), .B(new_n428), .C1(KEYINPUT39), .C2(new_n450), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT40), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n432), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n454), .B1(new_n453), .B2(new_n452), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n309), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT38), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n306), .A2(new_n307), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT81), .B(KEYINPUT37), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n299), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT37), .B1(new_n306), .B2(new_n307), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n457), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n282), .A2(new_n294), .A3(new_n296), .A4(new_n459), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n269), .A2(new_n293), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT37), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n465), .B1(new_n292), .B2(new_n280), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT38), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(new_n305), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n468), .A2(new_n435), .A3(new_n300), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n456), .B(new_n439), .C1(new_n462), .C2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT36), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(new_n353), .B2(new_n407), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n443), .A2(KEYINPUT36), .A3(new_n440), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n445), .A2(new_n406), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n470), .B1(KEYINPUT80), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n445), .A2(new_n406), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n472), .A2(new_n473), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT80), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n448), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G50gat), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT85), .B1(new_n480), .B2(G43gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(KEYINPUT15), .ZN(new_n482));
  XOR2_X1   g281(.A(G43gat), .B(G50gat), .Z(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n485));
  INV_X1    g284(.A(G29gat), .ZN(new_n486));
  INV_X1    g285(.A(G36gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT83), .B1(G29gat), .B2(G36gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(KEYINPUT14), .A3(new_n489), .ZN(new_n490));
  OAI221_X1 g289(.A(new_n490), .B1(KEYINPUT14), .B2(new_n489), .C1(new_n486), .C2(new_n487), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n484), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT15), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n483), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT84), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n495), .A2(new_n496), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(KEYINPUT17), .A3(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G15gat), .B(G22gat), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n503), .A2(G1gat), .ZN(new_n504));
  AOI21_X1  g303(.A(G8gat), .B1(new_n504), .B2(KEYINPUT86), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT16), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n503), .B1(new_n506), .B2(G1gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(new_n505), .B(new_n508), .Z(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(new_n498), .B2(new_n500), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n502), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n501), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n509), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT18), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n515), .B(new_n510), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n514), .B(KEYINPUT13), .Z(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n517), .A2(new_n518), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n519), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G169gat), .B(G197gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(KEYINPUT12), .Z(new_n531));
  OR2_X1    g330(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n525), .A2(new_n531), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n479), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT88), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT89), .ZN(new_n543));
  INV_X1    g342(.A(G57gat), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n542), .B(G64gat), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(G64gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT88), .ZN(new_n547));
  INV_X1    g346(.A(G64gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(G57gat), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n545), .B(new_n547), .C1(new_n543), .C2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT90), .ZN(new_n551));
  NOR2_X1   g350(.A1(G71gat), .A2(G78gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT9), .ZN(new_n553));
  NAND2_X1  g352(.A1(G71gat), .A2(G78gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n551), .B1(new_n550), .B2(new_n555), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n552), .B1(KEYINPUT87), .B2(new_n554), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(KEYINPUT87), .B2(new_n554), .ZN(new_n561));
  NOR2_X1   g360(.A1(KEYINPUT87), .A2(KEYINPUT9), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n562), .B1(new_n546), .B2(new_n549), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT91), .B1(new_n559), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n555), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT90), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n564), .B1(new_n568), .B2(new_n556), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT91), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n565), .A2(new_n566), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G231gat), .A2(G233gat), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n576), .B(KEYINPUT92), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n565), .A2(new_n571), .A3(new_n566), .A4(new_n573), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n578), .B1(new_n575), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n541), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n575), .A2(new_n579), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n577), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n540), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n565), .A2(new_n571), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n509), .B1(new_n587), .B2(KEYINPUT21), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n582), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n589), .B1(new_n582), .B2(new_n586), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n539), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n582), .A2(new_n586), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(new_n588), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n582), .A2(new_n586), .A3(new_n589), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(new_n538), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n592), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n592), .B2(new_n596), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n537), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n590), .A2(new_n591), .A3(new_n539), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n538), .B1(new_n594), .B2(new_n595), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n597), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n592), .A2(new_n596), .A3(new_n598), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(new_n536), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G134gat), .B(G162gat), .Z(new_n607));
  AOI21_X1  g406(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  INV_X1    g409(.A(G85gat), .ZN(new_n611));
  INV_X1    g410(.A(G92gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(KEYINPUT8), .A2(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(G85gat), .A3(G92gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT7), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G99gat), .B(G106gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT99), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n621), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n623), .A2(new_n615), .A3(new_n618), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT100), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(new_n624), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n502), .A2(new_n512), .A3(new_n626), .A4(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AOI22_X1  g430(.A1(new_n626), .A2(new_n629), .B1(new_n499), .B2(new_n501), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT41), .ZN(new_n633));
  INV_X1    g432(.A(G232gat), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n633), .A2(new_n634), .A3(new_n328), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT101), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n629), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n627), .A2(new_n628), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n515), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n640));
  INV_X1    g439(.A(new_n635), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n631), .B1(new_n636), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G190gat), .B(G218gat), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n609), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n636), .A2(new_n642), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n630), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n644), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n650), .B1(new_n646), .B2(new_n649), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n643), .A2(new_n645), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n649), .A2(KEYINPUT102), .A3(new_n654), .ZN(new_n655));
  OR3_X1    g454(.A1(new_n648), .A2(KEYINPUT102), .A3(new_n644), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(new_n656), .A3(new_n609), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G230gat), .A2(G233gat), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT104), .B1(new_n627), .B2(new_n569), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(new_n587), .B2(new_n627), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n565), .A2(new_n625), .A3(KEYINPUT104), .A4(new_n571), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT10), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n626), .A2(new_n629), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n665), .A2(KEYINPUT10), .A3(new_n587), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n660), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(G120gat), .B(G148gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(G176gat), .B(G204gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n668), .B(new_n669), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n662), .A2(new_n663), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n671), .A2(new_n660), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n667), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n660), .B(KEYINPUT105), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n664), .B2(new_n666), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n672), .ZN(new_n678));
  INV_X1    g477(.A(new_n670), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n674), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  AOI211_X1 g479(.A(KEYINPUT106), .B(new_n670), .C1(new_n677), .C2(new_n672), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n673), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n601), .A2(new_n606), .A3(new_n659), .A4(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n535), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n435), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G1gat), .ZN(G1324gat));
  AND4_X1   g487(.A1(new_n534), .A2(new_n479), .A3(new_n309), .A4(new_n685), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(G8gat), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n691), .B1(new_n692), .B2(new_n689), .ZN(new_n693));
  MUX2_X1   g492(.A(new_n691), .B(new_n693), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g493(.A(G15gat), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n353), .A2(new_n407), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n686), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n472), .A2(new_n473), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT107), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n686), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n697), .B1(new_n700), .B2(new_n695), .ZN(G1326gat));
  XNOR2_X1  g500(.A(KEYINPUT43), .B(G22gat), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n535), .A2(new_n406), .A3(new_n685), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT108), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n704), .A2(KEYINPUT108), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n707), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(new_n705), .A3(new_n702), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(G1327gat));
  NAND2_X1  g510(.A1(new_n601), .A2(new_n606), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n713), .A2(new_n659), .A3(new_n682), .ZN(new_n714));
  AND4_X1   g513(.A1(new_n486), .A2(new_n535), .A3(new_n435), .A4(new_n714), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n715), .A2(KEYINPUT45), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n435), .A2(new_n300), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(new_n460), .B2(new_n467), .ZN(new_n719));
  INV_X1    g518(.A(new_n461), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n463), .A2(new_n305), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT38), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n406), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n698), .B1(new_n723), .B2(new_n456), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n445), .A2(KEYINPUT110), .A3(new_n406), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT110), .B1(new_n445), .B2(new_n406), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n447), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n717), .B1(new_n728), .B2(new_n659), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n659), .A2(new_n717), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n479), .A2(new_n730), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n599), .A2(new_n600), .A3(new_n537), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n536), .B1(new_n604), .B2(new_n605), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n601), .A2(new_n606), .A3(KEYINPUT109), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n534), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n738), .A2(new_n739), .A3(new_n682), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n732), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G29gat), .B1(new_n741), .B2(new_n436), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n715), .A2(KEYINPUT45), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n716), .A2(new_n742), .A3(new_n743), .ZN(G1328gat));
  OAI21_X1  g543(.A(G36gat), .B1(new_n741), .B2(new_n310), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n535), .A2(new_n487), .A3(new_n309), .A4(new_n714), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT46), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n746), .A2(KEYINPUT46), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(G1329gat));
  INV_X1    g548(.A(new_n696), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(G43gat), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n479), .A2(new_n534), .A3(new_n714), .A4(new_n751), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n752), .A2(KEYINPUT111), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(KEYINPUT111), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n729), .A2(new_n731), .A3(new_n698), .A4(new_n740), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(G43gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n755), .A2(KEYINPUT47), .A3(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n729), .A2(new_n731), .A3(new_n699), .A4(new_n740), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n753), .A2(new_n754), .B1(new_n759), .B2(G43gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(KEYINPUT47), .B2(new_n760), .ZN(G1330gat));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n729), .A2(new_n731), .A3(new_n406), .A4(new_n740), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(G50gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n406), .A2(new_n480), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT112), .Z(new_n766));
  AND4_X1   g565(.A1(new_n534), .A2(new_n479), .A3(new_n714), .A4(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n763), .B2(G50gat), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT48), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n764), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI221_X4 g569(.A(new_n767), .B1(new_n762), .B2(KEYINPUT48), .C1(new_n763), .C2(G50gat), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(G1331gat));
  INV_X1    g571(.A(new_n726), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n445), .A2(KEYINPUT110), .A3(new_n406), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n470), .A2(new_n773), .A3(new_n477), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n448), .ZN(new_n776));
  NOR4_X1   g575(.A1(new_n712), .A2(new_n534), .A3(new_n658), .A4(new_n683), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n436), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(new_n544), .ZN(G1332gat));
  NOR2_X1   g579(.A1(new_n778), .A2(new_n310), .ZN(new_n781));
  NOR2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  AND2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(G1333gat));
  NAND4_X1  g584(.A1(new_n776), .A2(G71gat), .A3(new_n699), .A4(new_n777), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n778), .A2(new_n750), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(KEYINPUT114), .ZN(new_n788));
  INV_X1    g587(.A(G71gat), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n787), .B2(KEYINPUT114), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n786), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT50), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n793), .B(new_n786), .C1(new_n788), .C2(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1334gat));
  NOR2_X1   g594(.A1(new_n778), .A2(new_n439), .ZN(new_n796));
  XNOR2_X1  g595(.A(KEYINPUT115), .B(G78gat), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n796), .B(new_n797), .ZN(G1335gat));
  NOR3_X1   g597(.A1(new_n713), .A2(new_n534), .A3(new_n683), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n732), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G85gat), .B1(new_n800), .B2(new_n436), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n659), .B1(new_n775), .B2(new_n448), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n713), .A2(new_n534), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n802), .A2(KEYINPUT51), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT51), .B1(new_n802), .B2(new_n803), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n683), .A2(new_n436), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(new_n611), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n801), .A2(new_n808), .ZN(G1336gat));
  NAND4_X1  g608(.A1(new_n729), .A2(new_n731), .A3(new_n309), .A4(new_n799), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G92gat), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n309), .A2(new_n612), .A3(new_n682), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT116), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n804), .B2(new_n805), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g615(.A(new_n699), .ZN(new_n817));
  OAI21_X1  g616(.A(G99gat), .B1(new_n800), .B2(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n750), .A2(new_n683), .A3(G99gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n806), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(G1338gat));
  NAND4_X1  g620(.A1(new_n729), .A2(new_n731), .A3(new_n406), .A4(new_n799), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G106gat), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n439), .A2(new_n683), .A3(G106gat), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n804), .B2(new_n805), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(KEYINPUT117), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n827), .A3(KEYINPUT53), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n823), .B(new_n825), .C1(KEYINPUT117), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(G1339gat));
  NAND2_X1  g630(.A1(new_n520), .A2(new_n522), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n514), .B1(new_n513), .B2(new_n516), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n530), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n682), .A2(new_n532), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT10), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n671), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n666), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n842), .A3(new_n675), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n843), .A2(new_n667), .A3(KEYINPUT54), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n845), .B(new_n676), .C1(new_n664), .C2(new_n666), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n679), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n839), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n843), .A2(KEYINPUT54), .A3(new_n667), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n849), .A2(KEYINPUT55), .A3(new_n679), .A4(new_n846), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n673), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n838), .B1(new_n739), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n532), .A2(new_n837), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n853), .B1(new_n653), .B2(new_n657), .ZN(new_n854));
  INV_X1    g653(.A(new_n851), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n852), .A2(new_n659), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n736), .B2(new_n737), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n685), .A2(new_n739), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n750), .A2(new_n436), .A3(new_n406), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n310), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n739), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(new_n313), .ZN(G1340gat));
  NOR2_X1   g663(.A1(new_n862), .A2(new_n683), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(new_n311), .ZN(G1341gat));
  OAI21_X1  g665(.A(new_n319), .B1(new_n862), .B2(new_n712), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n738), .A2(G127gat), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT119), .B1(new_n862), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n862), .A2(KEYINPUT119), .A3(new_n868), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(G1342gat));
  NAND2_X1  g671(.A1(new_n310), .A2(new_n658), .ZN(new_n873));
  XNOR2_X1  g672(.A(KEYINPUT69), .B(G134gat), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n861), .A3(new_n875), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n876), .A2(KEYINPUT120), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(KEYINPUT120), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n877), .A2(KEYINPUT56), .A3(new_n878), .ZN(new_n882));
  OAI21_X1  g681(.A(G134gat), .B1(new_n862), .B2(new_n659), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(G1343gat));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n684), .A2(new_n534), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n885), .B(new_n406), .C1(new_n857), .C2(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n698), .A2(new_n436), .A3(new_n309), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n851), .A2(KEYINPUT121), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n848), .A2(new_n850), .A3(new_n890), .A4(new_n673), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n889), .A2(new_n534), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n658), .B1(new_n892), .B2(new_n838), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n854), .A2(new_n855), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n712), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n439), .B1(new_n895), .B2(new_n859), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n887), .B(new_n888), .C1(new_n896), .C2(new_n885), .ZN(new_n897));
  OAI21_X1  g696(.A(G141gat), .B1(new_n897), .B2(new_n739), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n439), .B1(new_n858), .B2(new_n859), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n699), .A2(new_n436), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n739), .A2(G141gat), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n901), .A2(new_n310), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n900), .A2(new_n905), .A3(KEYINPUT58), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT58), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n898), .B(new_n904), .C1(new_n899), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1344gat));
  NAND2_X1  g708(.A1(new_n901), .A2(new_n902), .ZN(new_n910));
  OR4_X1    g709(.A1(G148gat), .A2(new_n910), .A3(new_n309), .A4(new_n683), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n897), .A2(new_n683), .ZN(new_n912));
  INV_X1    g711(.A(G148gat), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n912), .A2(KEYINPUT59), .A3(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n915));
  OAI211_X1 g714(.A(KEYINPUT57), .B(new_n406), .C1(new_n857), .C2(new_n886), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n916), .B1(new_n896), .B2(KEYINPUT57), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n917), .A2(new_n310), .A3(new_n477), .A4(new_n807), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n915), .B1(new_n918), .B2(G148gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n911), .B1(new_n914), .B2(new_n919), .ZN(G1345gat));
  OR4_X1    g719(.A1(G155gat), .A2(new_n910), .A3(new_n309), .A4(new_n712), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n736), .A2(new_n737), .ZN(new_n922));
  OAI21_X1  g721(.A(G155gat), .B1(new_n897), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1346gat));
  OAI21_X1  g723(.A(G162gat), .B1(new_n897), .B2(new_n659), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n873), .A2(G162gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n910), .B2(new_n926), .ZN(G1347gat));
  NAND2_X1  g726(.A1(new_n309), .A2(new_n436), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n928), .A2(new_n444), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n860), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n534), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n932), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT123), .B1(new_n932), .B2(G169gat), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n933), .A2(new_n934), .B1(G169gat), .B2(new_n932), .ZN(G1348gat));
  NAND2_X1  g734(.A1(new_n931), .A2(new_n682), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(G176gat), .ZN(G1349gat));
  NAND4_X1  g736(.A1(new_n931), .A2(new_n239), .A3(new_n241), .A4(new_n713), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n939));
  OAI21_X1  g738(.A(G183gat), .B1(new_n930), .B2(new_n922), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT60), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT60), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n938), .A2(new_n940), .A3(new_n939), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1350gat));
  OAI211_X1 g744(.A(KEYINPUT61), .B(G190gat), .C1(new_n930), .C2(new_n659), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n930), .A2(new_n659), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(new_n212), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n948), .A2(KEYINPUT125), .A3(new_n212), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT125), .B1(new_n948), .B2(new_n212), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n946), .B(new_n949), .C1(new_n950), .C2(new_n951), .ZN(G1351gat));
  NOR2_X1   g751(.A1(new_n699), .A2(new_n928), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n901), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n534), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n953), .B(KEYINPUT126), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(new_n917), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n534), .A2(G197gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n682), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G204gat), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n683), .A2(G204gat), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n901), .A2(new_n953), .A3(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT62), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n962), .A2(new_n965), .ZN(G1353gat));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n967));
  OAI21_X1  g766(.A(G211gat), .B1(new_n967), .B2(KEYINPUT63), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n699), .A2(new_n712), .A3(new_n928), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n917), .B2(new_n969), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n967), .A2(KEYINPUT63), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n970), .B(new_n971), .ZN(new_n972));
  OR3_X1    g771(.A1(new_n954), .A2(G211gat), .A3(new_n712), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1354gat));
  AOI21_X1  g773(.A(G218gat), .B1(new_n955), .B2(new_n658), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n658), .A2(G218gat), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n958), .B2(new_n976), .ZN(G1355gat));
endmodule


