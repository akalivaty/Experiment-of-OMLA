//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n590, new_n591, new_n594, new_n596, new_n597, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  NAND2_X1  g033(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g036(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n460), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n460), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT65), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n474), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n466), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n463), .A2(G136), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n476), .B1(new_n461), .B2(new_n462), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n476), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  AND3_X1   g060(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n487));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G114), .C2(new_n476), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n470), .B2(new_n473), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n463), .B2(G138), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n491), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT67), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT65), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT65), .B1(new_n471), .B2(new_n472), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n493), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n476), .B1(new_n486), .B2(new_n487), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT4), .B1(new_n503), .B2(new_n492), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(new_n491), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  NAND2_X1  g084(.A1(KEYINPUT68), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n510), .B(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(G543), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n515), .A2(new_n521), .ZN(G166));
  AND2_X1   g097(.A1(new_n512), .A2(new_n516), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n525), .B(new_n527), .C1(new_n520), .C2(new_n528), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n524), .A2(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  AOI22_X1  g106(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n514), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n517), .A2(new_n534), .B1(new_n535), .B2(new_n520), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  AOI22_X1  g112(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n514), .ZN(new_n539));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  INV_X1    g115(.A(G43), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n517), .A2(new_n540), .B1(new_n541), .B2(new_n520), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT69), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  INV_X1    g124(.A(new_n520), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n550), .A2(KEYINPUT70), .A3(G53), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT9), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n514), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n523), .A2(G91), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(G299));
  INV_X1    g131(.A(G171), .ZN(G301));
  INV_X1    g132(.A(G166), .ZN(G303));
  NAND2_X1  g133(.A1(new_n523), .A2(G87), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n550), .A2(G49), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(G288));
  AOI22_X1  g137(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(new_n514), .ZN(new_n564));
  INV_X1    g139(.A(G86), .ZN(new_n565));
  INV_X1    g140(.A(G48), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n517), .A2(new_n565), .B1(new_n566), .B2(new_n520), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n564), .A2(new_n567), .ZN(G305));
  AOI22_X1  g143(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT71), .ZN(new_n570));
  OR3_X1    g145(.A1(new_n569), .A2(new_n570), .A3(new_n514), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n569), .B2(new_n514), .ZN(new_n572));
  XNOR2_X1  g147(.A(KEYINPUT72), .B(G85), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n523), .A2(new_n573), .B1(G47), .B2(new_n550), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(G301), .A2(G868), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n512), .A2(G92), .A3(new_n516), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT73), .Z(new_n578));
  INV_X1    g153(.A(KEYINPUT10), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n550), .A2(G54), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n582), .B2(new_n514), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT74), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n577), .B(KEYINPUT73), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT10), .ZN(new_n586));
  AND3_X1   g161(.A1(new_n580), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n576), .B1(new_n587), .B2(G868), .ZN(G284));
  OAI21_X1  g163(.A(new_n576), .B1(new_n587), .B2(G868), .ZN(G321));
  NAND2_X1  g164(.A1(G286), .A2(G868), .ZN(new_n590));
  INV_X1    g165(.A(G299), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(G868), .ZN(G297));
  OAI21_X1  g167(.A(new_n590), .B1(new_n591), .B2(G868), .ZN(G280));
  INV_X1    g168(.A(G559), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n587), .B1(new_n594), .B2(G860), .ZN(G148));
  NAND2_X1  g170(.A1(new_n587), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G868), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g173(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g174(.A1(new_n474), .A2(new_n465), .ZN(new_n600));
  XOR2_X1   g175(.A(new_n600), .B(KEYINPUT76), .Z(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT75), .B(KEYINPUT12), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XOR2_X1   g178(.A(KEYINPUT77), .B(KEYINPUT13), .Z(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G2100), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  OAI21_X1  g183(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n609));
  INV_X1    g184(.A(G111), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G2105), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n480), .A2(G123), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT78), .ZN(new_n613));
  AOI211_X1 g188(.A(new_n611), .B(new_n613), .C1(G135), .C2(new_n463), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2096), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n607), .A2(new_n608), .A3(new_n615), .ZN(G156));
  XNOR2_X1  g191(.A(KEYINPUT15), .B(G2435), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT79), .B(G2438), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(G2427), .B(G2430), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n621), .A2(KEYINPUT14), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(G2451), .B(G2454), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(G1341), .B(G1348), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n623), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  AND2_X1   g205(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(G14), .B1(new_n628), .B2(new_n630), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n631), .A2(new_n632), .ZN(G401));
  XNOR2_X1  g208(.A(G2072), .B(G2078), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT17), .Z(new_n635));
  XNOR2_X1  g210(.A(G2067), .B(G2678), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2084), .B(G2090), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT80), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n634), .A2(new_n636), .ZN(new_n641));
  NOR3_X1   g216(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT82), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n635), .A2(new_n637), .A3(new_n640), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT83), .Z(new_n645));
  NAND3_X1  g220(.A1(new_n640), .A2(new_n636), .A3(new_n634), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT81), .B(KEYINPUT18), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n643), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2096), .B(G2100), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(G227));
  XNOR2_X1  g226(.A(G1971), .B(G1976), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT19), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  XOR2_X1   g230(.A(G1961), .B(G1966), .Z(new_n656));
  AND2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT20), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n655), .A2(new_n656), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n654), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n654), .B2(new_n660), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G1981), .ZN(new_n664));
  INV_X1    g239(.A(G1986), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT85), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT84), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  OR3_X1    g248(.A1(new_n668), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n673), .B1(new_n668), .B2(new_n669), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(G229));
  NOR2_X1   g251(.A1(G4), .A2(G16), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n587), .B2(G16), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT91), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n679), .A2(G1348), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(G1348), .ZN(new_n681));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NOR2_X1   g257(.A1(G286), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT96), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(KEYINPUT96), .B1(G16), .B2(G21), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n687), .A2(G1966), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT97), .ZN(new_n689));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G26), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT28), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n463), .A2(G140), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n480), .A2(G128), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n476), .A2(G116), .ZN(new_n695));
  OAI21_X1  g270(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n693), .B(new_n694), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n692), .B1(new_n697), .B2(G29), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G2067), .ZN(new_n699));
  INV_X1    g274(.A(new_n687), .ZN(new_n700));
  INV_X1    g275(.A(G1966), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n690), .A2(G35), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G162), .B2(new_n690), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT29), .Z(new_n705));
  INV_X1    g280(.A(G2090), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G171), .A2(new_n682), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G5), .B2(new_n682), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G16), .A2(G19), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n543), .B2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT92), .B(G1341), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n710), .A2(G1961), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  INV_X1    g290(.A(G11), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(KEYINPUT31), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(KEYINPUT31), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT30), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n719), .A2(G28), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n690), .B1(new_n719), .B2(G28), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n717), .B(new_n718), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n614), .B2(G29), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n707), .A2(new_n714), .A3(new_n715), .A4(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT24), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n690), .B1(new_n725), .B2(G34), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n725), .B2(G34), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G160), .B2(G29), .ZN(new_n728));
  AOI211_X1 g303(.A(new_n702), .B(new_n724), .C1(G2084), .C2(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n680), .A2(new_n681), .A3(new_n689), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n463), .A2(G139), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT25), .Z(new_n733));
  AOI22_X1  g308(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n731), .B(new_n733), .C1(new_n734), .C2(new_n476), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT93), .ZN(new_n736));
  MUX2_X1   g311(.A(G33), .B(new_n736), .S(G29), .Z(new_n737));
  XOR2_X1   g312(.A(KEYINPUT94), .B(G2072), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n690), .A2(G32), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT26), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n743), .A2(new_n744), .B1(G105), .B2(new_n465), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n463), .A2(G141), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n480), .A2(G129), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n740), .B1(new_n749), .B2(new_n690), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT95), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n682), .A2(G20), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT23), .Z(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G299), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1956), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  AOI211_X1 g334(.A(new_n754), .B(new_n759), .C1(new_n706), .C2(new_n705), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n690), .A2(G27), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G164), .B2(new_n690), .ZN(new_n762));
  INV_X1    g337(.A(G2078), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G1961), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n709), .A2(new_n765), .B1(new_n750), .B2(new_n752), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G2084), .B2(new_n728), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT98), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n739), .A2(new_n760), .A3(new_n764), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n730), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n682), .A2(G23), .ZN(new_n772));
  INV_X1    g347(.A(G288), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n682), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(KEYINPUT87), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(KEYINPUT87), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT33), .B(G1976), .Z(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n775), .A2(new_n778), .A3(new_n776), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n682), .A2(G22), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G166), .B2(new_n682), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G1971), .Z(new_n784));
  NOR2_X1   g359(.A1(G6), .A2(G16), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n564), .A2(new_n567), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(G16), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT32), .B(G1981), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n780), .A2(new_n781), .A3(new_n784), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(KEYINPUT34), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n463), .A2(G131), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n480), .A2(G119), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n476), .A2(G107), .ZN(new_n795));
  OAI21_X1  g370(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n793), .B(new_n794), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G25), .B(new_n797), .S(G29), .Z(new_n798));
  XOR2_X1   g373(.A(KEYINPUT35), .B(G1991), .Z(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(new_n800), .ZN(new_n801));
  MUX2_X1   g376(.A(G24), .B(G290), .S(G16), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(new_n665), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT86), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI221_X1 g380(.A(new_n805), .B1(new_n804), .B2(new_n803), .C1(new_n790), .C2(KEYINPUT34), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(KEYINPUT88), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(KEYINPUT88), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n792), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT36), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT89), .B(KEYINPUT36), .Z(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT90), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n811), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n809), .A2(new_n813), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT90), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n771), .B1(new_n816), .B2(new_n818), .ZN(G311));
  INV_X1    g394(.A(new_n818), .ZN(new_n820));
  OAI22_X1  g395(.A1(new_n817), .A2(KEYINPUT90), .B1(new_n810), .B2(new_n809), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n770), .B1(new_n820), .B2(new_n821), .ZN(G150));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n584), .A3(new_n586), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n823), .A2(new_n594), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(G93), .ZN(new_n827));
  INV_X1    g402(.A(G55), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n517), .A2(new_n827), .B1(new_n828), .B2(new_n520), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT100), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(new_n514), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n539), .B2(new_n542), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n831), .A2(new_n543), .A3(new_n833), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n826), .B(new_n837), .Z(new_n838));
  INV_X1    g413(.A(KEYINPUT39), .ZN(new_n839));
  AOI21_X1  g414(.A(G860), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n834), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(G145));
  XNOR2_X1  g419(.A(new_n477), .B(G162), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n614), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n480), .A2(G130), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n476), .A2(G118), .ZN(new_n848));
  OAI21_X1  g423(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(G142), .B2(new_n463), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n797), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n603), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT102), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n498), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n505), .A2(KEYINPUT101), .A3(new_n491), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n697), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n736), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n749), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n854), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n854), .A2(new_n861), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n846), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(KEYINPUT103), .B(G37), .Z(new_n865));
  OR2_X1    g440(.A1(new_n863), .A2(new_n846), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n861), .A2(new_n853), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n864), .B(new_n865), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g444(.A(G868), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n834), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n596), .B(new_n837), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n587), .A2(G299), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n823), .A2(new_n874), .A3(new_n591), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n874), .B1(new_n823), .B2(new_n591), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n872), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT105), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n876), .A2(new_n878), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n876), .A2(new_n885), .A3(KEYINPUT41), .A4(new_n878), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n878), .A2(KEYINPUT41), .A3(new_n873), .A4(new_n875), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT106), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n872), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n881), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(G290), .B(new_n773), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n892), .A2(KEYINPUT107), .ZN(new_n893));
  XNOR2_X1  g468(.A(G305), .B(G166), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n894), .B1(new_n892), .B2(KEYINPUT107), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n894), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n896), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(KEYINPUT108), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n900), .B(KEYINPUT42), .Z(new_n901));
  XNOR2_X1  g476(.A(new_n891), .B(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n871), .B1(new_n902), .B2(new_n870), .ZN(G295));
  OAI21_X1  g478(.A(new_n871), .B1(new_n902), .B2(new_n870), .ZN(G331));
  XNOR2_X1  g479(.A(G286), .B(G171), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n837), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n835), .B2(new_n836), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n907), .A2(KEYINPUT109), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n837), .A2(KEYINPUT109), .A3(new_n906), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n889), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n907), .A2(new_n908), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n882), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n915), .B2(new_n898), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n899), .A3(new_n914), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT43), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n917), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n913), .B1(new_n884), .B2(new_n887), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n879), .B1(new_n909), .B2(new_n910), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n898), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n865), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n919), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT44), .B1(new_n918), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n924), .B1(new_n916), .B2(new_n917), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n919), .A2(new_n923), .A3(KEYINPUT43), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n930), .ZN(G397));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(new_n858), .B2(G1384), .ZN(new_n933));
  OAI211_X1 g508(.A(G40), .B(new_n466), .C1(new_n475), .C2(new_n476), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G1996), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT46), .ZN(new_n938));
  INV_X1    g513(.A(new_n935), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n697), .B(G2067), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT110), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n941), .A2(new_n749), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n938), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT125), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n943), .A2(KEYINPUT125), .ZN(new_n947));
  OR3_X1    g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n748), .B(new_n936), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n941), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n797), .A2(new_n800), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n697), .A2(G2067), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n939), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n797), .B(new_n799), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n951), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(G290), .A2(G1986), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n935), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n957), .A2(new_n935), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n955), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n948), .A2(new_n949), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n498), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n934), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(KEYINPUT112), .B(G8), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(G305), .A2(G1981), .ZN(new_n970));
  XNOR2_X1  g545(.A(KEYINPUT113), .B(G1981), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n786), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT49), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT114), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n977));
  AOI211_X1 g552(.A(new_n977), .B(KEYINPUT49), .C1(new_n970), .C2(new_n973), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n969), .B1(new_n974), .B2(new_n975), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n981), .A2(G1976), .A3(G288), .ZN(new_n982));
  INV_X1    g557(.A(new_n973), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n969), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G8), .ZN(new_n985));
  INV_X1    g560(.A(new_n934), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n932), .A2(G1384), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n856), .A2(new_n857), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(G1384), .B1(new_n499), .B2(new_n507), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n986), .B(new_n988), .C1(new_n989), .C2(KEYINPUT45), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n991), .A2(G1971), .ZN(new_n992));
  AOI21_X1  g567(.A(G1384), .B1(new_n505), .B2(new_n491), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT111), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n989), .B2(new_n994), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n488), .A2(new_n490), .ZN(new_n997));
  AOI211_X1 g572(.A(KEYINPUT67), .B(new_n997), .C1(new_n502), .C2(new_n504), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n506), .B1(new_n505), .B2(new_n491), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n965), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n934), .B1(new_n996), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n706), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n985), .B1(new_n992), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G303), .A2(G8), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT55), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1976), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT52), .B1(G288), .B2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n969), .B(new_n1010), .C1(new_n1009), .C2(G288), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n969), .B1(new_n1009), .B2(G288), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT52), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1011), .B(new_n1013), .C1(new_n979), .C2(new_n980), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n984), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT63), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1014), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n991), .A2(G1971), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n508), .A2(new_n994), .A3(new_n965), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n934), .B1(KEYINPUT50), .B2(new_n966), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(G2090), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1018), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1006), .B1(new_n1023), .B2(new_n968), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1017), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G2084), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1002), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n934), .B1(new_n932), .B2(new_n966), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1966), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n968), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G168), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1016), .B1(new_n1025), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1016), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1035), .B(new_n1017), .C1(new_n1007), .C2(new_n1004), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1015), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(G168), .A2(new_n968), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1032), .A2(KEYINPUT51), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1030), .B1(new_n1002), .B2(new_n1026), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT120), .B1(new_n1040), .B2(new_n985), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1038), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n1043));
  AOI211_X1 g618(.A(G2084), .B(new_n934), .C1(new_n996), .C2(new_n1001), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1043), .B(G8), .C1(new_n1044), .C2(new_n1030), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(new_n1042), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n1032), .B2(G286), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1039), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT62), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n996), .A2(new_n1001), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n986), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n765), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1028), .A2(KEYINPUT53), .A3(new_n763), .A4(new_n1029), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT122), .B(new_n1055), .C1(new_n990), .C2(G2078), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n988), .A2(new_n986), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1000), .A2(new_n932), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(new_n763), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT122), .B1(new_n1060), .B2(new_n1055), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1053), .B(new_n1054), .C1(new_n1057), .C2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(G171), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1025), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1050), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1049), .A2(KEYINPUT62), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1037), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n989), .A2(KEYINPUT45), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n988), .A2(new_n986), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT56), .B(G2072), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1068), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(G1956), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1073));
  NAND2_X1  g648(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n1074));
  NOR2_X1   g649(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(G299), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1078), .A2(new_n1079), .B1(G91), .B2(new_n523), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .A4(new_n554), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1077), .A2(new_n1083), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1072), .A2(new_n1073), .A3(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1002), .A2(G1348), .ZN(new_n1086));
  INV_X1    g661(.A(new_n967), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1087), .A2(G2067), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n587), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT116), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1021), .A2(new_n758), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1058), .A2(new_n1059), .A3(new_n1070), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1095), .A3(new_n1084), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1085), .B1(new_n1090), .B2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(KEYINPUT60), .B(new_n1088), .C1(new_n1002), .C2(G1348), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1098), .A2(KEYINPUT118), .A3(new_n823), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n823), .B1(new_n1098), .B2(KEYINPUT118), .ZN(new_n1100));
  OAI22_X1  g675(.A1(new_n1099), .A2(new_n1100), .B1(KEYINPUT118), .B2(new_n1098), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n1102), .A2(KEYINPUT60), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1073), .B1(new_n991), .B2(new_n1070), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1077), .A2(new_n1083), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1096), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1107), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1105), .B1(new_n1110), .B2(new_n1085), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n990), .B2(G1996), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1058), .A2(new_n1059), .A3(KEYINPUT117), .A4(new_n936), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT58), .B(G1341), .Z(new_n1115));
  NAND2_X1  g690(.A1(new_n1087), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n543), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1118), .B1(new_n1117), .B2(new_n543), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1109), .B(new_n1111), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  AOI211_X1 g697(.A(KEYINPUT119), .B(new_n1097), .C1(new_n1104), .C2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1098), .A2(KEYINPUT118), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1098), .A2(KEYINPUT118), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n587), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1098), .A2(KEYINPUT118), .A3(new_n823), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1127), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1102), .A2(KEYINPUT60), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1125), .B(new_n1126), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1097), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1124), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1123), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1058), .A2(KEYINPUT53), .A3(new_n933), .A4(new_n763), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1053), .B(new_n1138), .C1(new_n1057), .C2(new_n1061), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1139), .A2(G171), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1055), .B1(new_n990), .B2(G2078), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1143), .A2(new_n1056), .B1(new_n765), .B2(new_n1052), .ZN(new_n1144));
  AOI21_X1  g719(.A(G301), .B1(new_n1144), .B2(new_n1054), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1137), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1062), .B2(G171), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1137), .B1(new_n1139), .B2(G171), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1144), .A2(KEYINPUT123), .A3(G301), .A4(new_n1054), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1017), .A2(new_n1024), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1146), .A2(new_n1151), .A3(new_n1049), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT124), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1063), .B1(G171), .B2(new_n1139), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1025), .B1(new_n1155), .B2(new_n1137), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(new_n1151), .A4(new_n1049), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1154), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1067), .B1(new_n1136), .B2(new_n1159), .ZN(new_n1160));
  AND2_X1   g735(.A1(G290), .A2(G1986), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n957), .A2(new_n958), .A3(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1162), .A2(new_n939), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n964), .B1(new_n1160), .B2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g739(.A(G319), .B1(new_n631), .B2(new_n632), .ZN(new_n1166));
  NOR2_X1   g740(.A1(G227), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g741(.A1(new_n674), .A2(new_n675), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g744(.A1(new_n674), .A2(new_n675), .A3(KEYINPUT127), .A4(new_n1167), .ZN(new_n1171));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g746(.A(new_n1172), .B(new_n868), .C1(new_n928), .C2(new_n929), .ZN(G225));
  INV_X1    g747(.A(G225), .ZN(G308));
endmodule


