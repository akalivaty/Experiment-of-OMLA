

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U556 ( .A1(G164), .A2(G1384), .ZN(n715) );
  NOR2_X2 U557 ( .A1(G2104), .A2(n530), .ZN(n903) );
  OR2_X2 U558 ( .A1(n676), .A2(n674), .ZN(n658) );
  NOR2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XNOR2_X1 U560 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n524) );
  NOR2_X1 U561 ( .A1(G168), .A2(n652), .ZN(n654) );
  NAND2_X1 U562 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U563 ( .A1(G543), .A2(n539), .ZN(n540) );
  XNOR2_X1 U564 ( .A(n590), .B(n589), .ZN(n776) );
  XNOR2_X1 U565 ( .A(KEYINPUT97), .B(KEYINPUT32), .ZN(n521) );
  XOR2_X1 U566 ( .A(KEYINPUT86), .B(n672), .Z(n522) );
  INV_X1 U567 ( .A(KEYINPUT94), .ZN(n653) );
  XNOR2_X1 U568 ( .A(n670), .B(n521), .ZN(n685) );
  INV_X1 U569 ( .A(KEYINPUT101), .ZN(n701) );
  AND2_X1 U570 ( .A1(n775), .A2(n587), .ZN(n591) );
  INV_X1 U571 ( .A(G2105), .ZN(n530) );
  INV_X1 U572 ( .A(KEYINPUT13), .ZN(n601) );
  INV_X1 U573 ( .A(KEYINPUT23), .ZN(n589) );
  XNOR2_X1 U574 ( .A(n583), .B(KEYINPUT66), .ZN(n775) );
  XNOR2_X1 U575 ( .A(n524), .B(n523), .ZN(n582) );
  INV_X1 U576 ( .A(n582), .ZN(n525) );
  INV_X2 U577 ( .A(n525), .ZN(n899) );
  NAND2_X1 U578 ( .A1(G138), .A2(n899), .ZN(n529) );
  INV_X1 U579 ( .A(G2104), .ZN(n526) );
  NOR2_X1 U580 ( .A1(n526), .A2(G2105), .ZN(n527) );
  XNOR2_X1 U581 ( .A(n527), .B(KEYINPUT64), .ZN(n588) );
  BUF_X2 U582 ( .A(n588), .Z(n900) );
  NAND2_X1 U583 ( .A1(G102), .A2(n900), .ZN(n528) );
  NAND2_X1 U584 ( .A1(n529), .A2(n528), .ZN(n534) );
  NAND2_X1 U585 ( .A1(G126), .A2(n903), .ZN(n532) );
  AND2_X1 U586 ( .A1(G2105), .A2(G2104), .ZN(n904) );
  NAND2_X1 U587 ( .A1(G114), .A2(n904), .ZN(n531) );
  NAND2_X1 U588 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X2 U589 ( .A1(n534), .A2(n533), .ZN(G164) );
  NOR2_X2 U590 ( .A1(G651), .A2(G543), .ZN(n809) );
  NAND2_X1 U591 ( .A1(n809), .A2(G89), .ZN(n535) );
  XNOR2_X1 U592 ( .A(n535), .B(KEYINPUT4), .ZN(n537) );
  XOR2_X1 U593 ( .A(KEYINPUT0), .B(G543), .Z(n566) );
  INV_X1 U594 ( .A(G651), .ZN(n539) );
  NOR2_X2 U595 ( .A1(n566), .A2(n539), .ZN(n810) );
  NAND2_X1 U596 ( .A1(G76), .A2(n810), .ZN(n536) );
  NAND2_X1 U597 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U598 ( .A(n538), .B(KEYINPUT5), .ZN(n545) );
  XOR2_X2 U599 ( .A(KEYINPUT1), .B(n540), .Z(n805) );
  NAND2_X1 U600 ( .A1(G63), .A2(n805), .ZN(n542) );
  NOR2_X2 U601 ( .A1(G651), .A2(n566), .ZN(n806) );
  NAND2_X1 U602 ( .A1(G51), .A2(n806), .ZN(n541) );
  NAND2_X1 U603 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U604 ( .A(KEYINPUT6), .B(n543), .Z(n544) );
  NAND2_X1 U605 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U606 ( .A(n546), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U607 ( .A1(G64), .A2(n805), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G52), .A2(n806), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G90), .A2(n809), .ZN(n550) );
  NAND2_X1 U611 ( .A1(G77), .A2(n810), .ZN(n549) );
  NAND2_X1 U612 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U613 ( .A(KEYINPUT67), .B(n551), .ZN(n552) );
  XNOR2_X1 U614 ( .A(KEYINPUT9), .B(n552), .ZN(n553) );
  NOR2_X1 U615 ( .A1(n554), .A2(n553), .ZN(G171) );
  INV_X1 U616 ( .A(G171), .ZN(G301) );
  XOR2_X1 U617 ( .A(G168), .B(KEYINPUT8), .Z(n555) );
  XNOR2_X1 U618 ( .A(KEYINPUT70), .B(n555), .ZN(G286) );
  NAND2_X1 U619 ( .A1(G88), .A2(n809), .ZN(n557) );
  NAND2_X1 U620 ( .A1(G75), .A2(n810), .ZN(n556) );
  NAND2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U622 ( .A1(G62), .A2(n805), .ZN(n558) );
  XNOR2_X1 U623 ( .A(KEYINPUT75), .B(n558), .ZN(n559) );
  NOR2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U625 ( .A1(n806), .A2(G50), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n562), .A2(n561), .ZN(G303) );
  NAND2_X1 U627 ( .A1(G49), .A2(n806), .ZN(n564) );
  NAND2_X1 U628 ( .A1(G74), .A2(G651), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U630 ( .A1(n805), .A2(n565), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n566), .A2(G87), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(G288) );
  NAND2_X1 U633 ( .A1(G61), .A2(n805), .ZN(n570) );
  NAND2_X1 U634 ( .A1(G48), .A2(n806), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n810), .A2(G73), .ZN(n571) );
  XOR2_X1 U637 ( .A(KEYINPUT2), .B(n571), .Z(n572) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n809), .A2(G86), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(G305) );
  NAND2_X1 U641 ( .A1(G60), .A2(n805), .ZN(n577) );
  NAND2_X1 U642 ( .A1(G47), .A2(n806), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U644 ( .A1(G85), .A2(n809), .ZN(n579) );
  NAND2_X1 U645 ( .A1(G72), .A2(n810), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  OR2_X1 U647 ( .A1(n581), .A2(n580), .ZN(G290) );
  NAND2_X1 U648 ( .A1(G137), .A2(n582), .ZN(n583) );
  INV_X1 U649 ( .A(G40), .ZN(n586) );
  NAND2_X1 U650 ( .A1(G125), .A2(n903), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G113), .A2(n904), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n778) );
  NOR2_X1 U653 ( .A1(n586), .A2(n778), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n588), .A2(G101), .ZN(n590) );
  NAND2_X1 U655 ( .A1(n591), .A2(n776), .ZN(n714) );
  XNOR2_X1 U656 ( .A(n714), .B(KEYINPUT85), .ZN(n592) );
  NAND2_X1 U657 ( .A1(n715), .A2(n592), .ZN(n649) );
  NAND2_X1 U658 ( .A1(n649), .A2(G1341), .ZN(n593) );
  XNOR2_X1 U659 ( .A(n593), .B(KEYINPUT92), .ZN(n605) );
  NAND2_X1 U660 ( .A1(G56), .A2(n805), .ZN(n594) );
  XNOR2_X1 U661 ( .A(n594), .B(KEYINPUT14), .ZN(n597) );
  NAND2_X1 U662 ( .A1(G43), .A2(n806), .ZN(n595) );
  XOR2_X1 U663 ( .A(KEYINPUT69), .B(n595), .Z(n596) );
  NAND2_X1 U664 ( .A1(n597), .A2(n596), .ZN(n604) );
  NAND2_X1 U665 ( .A1(G68), .A2(n810), .ZN(n600) );
  NAND2_X1 U666 ( .A1(n809), .A2(G81), .ZN(n598) );
  XNOR2_X1 U667 ( .A(n598), .B(KEYINPUT12), .ZN(n599) );
  NAND2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n602) );
  XNOR2_X1 U669 ( .A(n602), .B(n601), .ZN(n603) );
  NOR2_X1 U670 ( .A1(n604), .A2(n603), .ZN(n1020) );
  NAND2_X1 U671 ( .A1(n605), .A2(n1020), .ZN(n608) );
  INV_X2 U672 ( .A(n649), .ZN(n642) );
  NAND2_X1 U673 ( .A1(G1996), .A2(n642), .ZN(n606) );
  XOR2_X1 U674 ( .A(n606), .B(KEYINPUT26), .Z(n607) );
  NOR2_X1 U675 ( .A1(n608), .A2(n607), .ZN(n619) );
  NAND2_X1 U676 ( .A1(G66), .A2(n805), .ZN(n610) );
  NAND2_X1 U677 ( .A1(G54), .A2(n806), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U679 ( .A1(G92), .A2(n809), .ZN(n612) );
  NAND2_X1 U680 ( .A1(G79), .A2(n810), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U682 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U683 ( .A(KEYINPUT15), .B(n615), .ZN(n916) );
  NOR2_X1 U684 ( .A1(n642), .A2(G1348), .ZN(n617) );
  BUF_X2 U685 ( .A(n649), .Z(n662) );
  NOR2_X1 U686 ( .A1(G2067), .A2(n662), .ZN(n616) );
  NOR2_X1 U687 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U688 ( .A1(n916), .A2(n620), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n619), .A2(n618), .ZN(n622) );
  OR2_X1 U690 ( .A1(n620), .A2(n916), .ZN(n621) );
  NAND2_X1 U691 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U692 ( .A(n623), .B(KEYINPUT93), .ZN(n634) );
  NAND2_X1 U693 ( .A1(n642), .A2(G2072), .ZN(n624) );
  XNOR2_X1 U694 ( .A(n624), .B(KEYINPUT27), .ZN(n626) );
  XNOR2_X1 U695 ( .A(G1956), .B(KEYINPUT89), .ZN(n980) );
  NOR2_X1 U696 ( .A1(n980), .A2(n642), .ZN(n625) );
  NOR2_X1 U697 ( .A1(n626), .A2(n625), .ZN(n635) );
  NAND2_X1 U698 ( .A1(G65), .A2(n805), .ZN(n628) );
  NAND2_X1 U699 ( .A1(G53), .A2(n806), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U701 ( .A1(G91), .A2(n809), .ZN(n630) );
  NAND2_X1 U702 ( .A1(G78), .A2(n810), .ZN(n629) );
  NAND2_X1 U703 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U704 ( .A1(n632), .A2(n631), .ZN(n1024) );
  NAND2_X1 U705 ( .A1(n635), .A2(n1024), .ZN(n633) );
  NAND2_X1 U706 ( .A1(n634), .A2(n633), .ZN(n640) );
  NOR2_X1 U707 ( .A1(n635), .A2(n1024), .ZN(n638) );
  XNOR2_X1 U708 ( .A(KEYINPUT28), .B(KEYINPUT91), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n636), .B(KEYINPUT90), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n638), .B(n637), .ZN(n639) );
  NAND2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U712 ( .A(n641), .B(KEYINPUT29), .ZN(n676) );
  NOR2_X1 U713 ( .A1(n642), .A2(G1961), .ZN(n643) );
  XOR2_X1 U714 ( .A(KEYINPUT87), .B(n643), .Z(n645) );
  XOR2_X1 U715 ( .A(G2078), .B(KEYINPUT25), .Z(n963) );
  NOR2_X1 U716 ( .A1(n963), .A2(n662), .ZN(n644) );
  NOR2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n647) );
  NOR2_X1 U718 ( .A1(n647), .A2(G301), .ZN(n646) );
  XNOR2_X1 U719 ( .A(KEYINPUT88), .B(n646), .ZN(n674) );
  NAND2_X1 U720 ( .A1(n647), .A2(G301), .ZN(n648) );
  XOR2_X1 U721 ( .A(KEYINPUT95), .B(n648), .Z(n656) );
  NAND2_X1 U722 ( .A1(n649), .A2(G8), .ZN(n661) );
  NOR2_X1 U723 ( .A1(G1966), .A2(n661), .ZN(n673) );
  NOR2_X1 U724 ( .A1(G2084), .A2(n662), .ZN(n671) );
  NOR2_X1 U725 ( .A1(n673), .A2(n671), .ZN(n650) );
  NAND2_X1 U726 ( .A1(G8), .A2(n650), .ZN(n651) );
  XNOR2_X1 U727 ( .A(KEYINPUT30), .B(n651), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n654), .B(n653), .ZN(n655) );
  NAND2_X1 U729 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n657), .B(KEYINPUT31), .ZN(n678) );
  NAND2_X1 U731 ( .A1(n658), .A2(n678), .ZN(n660) );
  AND2_X1 U732 ( .A1(G286), .A2(G8), .ZN(n659) );
  NAND2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n669) );
  INV_X1 U734 ( .A(G8), .ZN(n667) );
  NOR2_X1 U735 ( .A1(G1971), .A2(n661), .ZN(n664) );
  NOR2_X1 U736 ( .A1(G2090), .A2(n662), .ZN(n663) );
  NOR2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U738 ( .A1(n665), .A2(G303), .ZN(n666) );
  OR2_X1 U739 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U740 ( .A1(G8), .A2(n671), .ZN(n672) );
  OR2_X1 U741 ( .A1(n522), .A2(n673), .ZN(n677) );
  OR2_X1 U742 ( .A1(n674), .A2(n677), .ZN(n675) );
  OR2_X1 U743 ( .A1(n676), .A2(n675), .ZN(n682) );
  INV_X1 U744 ( .A(n677), .ZN(n680) );
  INV_X1 U745 ( .A(n678), .ZN(n679) );
  NAND2_X1 U746 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U748 ( .A(n683), .B(KEYINPUT96), .ZN(n684) );
  NAND2_X1 U749 ( .A1(n685), .A2(n684), .ZN(n705) );
  NOR2_X1 U750 ( .A1(G1971), .A2(G303), .ZN(n686) );
  NOR2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n1021) );
  NOR2_X1 U752 ( .A1(n686), .A2(n1021), .ZN(n687) );
  NAND2_X1 U753 ( .A1(n705), .A2(n687), .ZN(n688) );
  XNOR2_X1 U754 ( .A(n688), .B(KEYINPUT98), .ZN(n689) );
  NAND2_X1 U755 ( .A1(G1976), .A2(G288), .ZN(n1023) );
  NAND2_X1 U756 ( .A1(n689), .A2(n1023), .ZN(n690) );
  XNOR2_X1 U757 ( .A(n690), .B(KEYINPUT99), .ZN(n691) );
  INV_X1 U758 ( .A(n661), .ZN(n693) );
  NAND2_X1 U759 ( .A1(n691), .A2(n693), .ZN(n692) );
  INV_X1 U760 ( .A(KEYINPUT33), .ZN(n695) );
  NAND2_X1 U761 ( .A1(n692), .A2(n695), .ZN(n700) );
  NAND2_X1 U762 ( .A1(n693), .A2(n1021), .ZN(n694) );
  NOR2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U764 ( .A(n696), .B(KEYINPUT100), .Z(n698) );
  XNOR2_X1 U765 ( .A(G1981), .B(G305), .ZN(n1014) );
  INV_X1 U766 ( .A(n1014), .ZN(n697) );
  AND2_X1 U767 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n702) );
  XNOR2_X1 U769 ( .A(n702), .B(n701), .ZN(n708) );
  NOR2_X1 U770 ( .A1(G2090), .A2(G303), .ZN(n703) );
  NAND2_X1 U771 ( .A1(G8), .A2(n703), .ZN(n704) );
  NAND2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U773 ( .A1(n706), .A2(n661), .ZN(n707) );
  NAND2_X1 U774 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U775 ( .A(n709), .B(KEYINPUT102), .ZN(n713) );
  NOR2_X1 U776 ( .A1(G1981), .A2(G305), .ZN(n710) );
  XOR2_X1 U777 ( .A(n710), .B(KEYINPUT24), .Z(n711) );
  NOR2_X1 U778 ( .A1(n661), .A2(n711), .ZN(n712) );
  NOR2_X1 U779 ( .A1(n713), .A2(n712), .ZN(n746) );
  NOR2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n760) );
  NAND2_X1 U781 ( .A1(G140), .A2(n899), .ZN(n717) );
  NAND2_X1 U782 ( .A1(G104), .A2(n900), .ZN(n716) );
  NAND2_X1 U783 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U784 ( .A(KEYINPUT34), .B(n718), .ZN(n724) );
  NAND2_X1 U785 ( .A1(n904), .A2(G116), .ZN(n719) );
  XOR2_X1 U786 ( .A(KEYINPUT79), .B(n719), .Z(n721) );
  NAND2_X1 U787 ( .A1(n903), .A2(G128), .ZN(n720) );
  NAND2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U789 ( .A(KEYINPUT35), .B(n722), .Z(n723) );
  NOR2_X1 U790 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U791 ( .A(KEYINPUT36), .B(n725), .Z(n913) );
  XOR2_X1 U792 ( .A(KEYINPUT37), .B(G2067), .Z(n757) );
  AND2_X1 U793 ( .A1(n913), .A2(n757), .ZN(n936) );
  NAND2_X1 U794 ( .A1(n760), .A2(n936), .ZN(n755) );
  NAND2_X1 U795 ( .A1(G129), .A2(n903), .ZN(n727) );
  NAND2_X1 U796 ( .A1(G117), .A2(n904), .ZN(n726) );
  NAND2_X1 U797 ( .A1(n727), .A2(n726), .ZN(n731) );
  NAND2_X1 U798 ( .A1(n900), .A2(G105), .ZN(n728) );
  XNOR2_X1 U799 ( .A(n728), .B(KEYINPUT83), .ZN(n729) );
  XNOR2_X1 U800 ( .A(n729), .B(KEYINPUT38), .ZN(n730) );
  NOR2_X1 U801 ( .A1(n731), .A2(n730), .ZN(n733) );
  NAND2_X1 U802 ( .A1(n899), .A2(G141), .ZN(n732) );
  NAND2_X1 U803 ( .A1(n733), .A2(n732), .ZN(n895) );
  AND2_X1 U804 ( .A1(n895), .A2(G1996), .ZN(n947) );
  NAND2_X1 U805 ( .A1(G119), .A2(n903), .ZN(n734) );
  XNOR2_X1 U806 ( .A(n734), .B(KEYINPUT80), .ZN(n741) );
  NAND2_X1 U807 ( .A1(G131), .A2(n899), .ZN(n736) );
  NAND2_X1 U808 ( .A1(G107), .A2(n904), .ZN(n735) );
  NAND2_X1 U809 ( .A1(n736), .A2(n735), .ZN(n739) );
  NAND2_X1 U810 ( .A1(G95), .A2(n900), .ZN(n737) );
  XNOR2_X1 U811 ( .A(KEYINPUT81), .B(n737), .ZN(n738) );
  NOR2_X1 U812 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U814 ( .A(KEYINPUT82), .B(n742), .ZN(n910) );
  AND2_X1 U815 ( .A1(G1991), .A2(n910), .ZN(n952) );
  OR2_X1 U816 ( .A1(n947), .A2(n952), .ZN(n743) );
  NAND2_X1 U817 ( .A1(n760), .A2(n743), .ZN(n749) );
  NAND2_X1 U818 ( .A1(n755), .A2(n749), .ZN(n744) );
  XNOR2_X1 U819 ( .A(n744), .B(KEYINPUT84), .ZN(n745) );
  NOR2_X1 U820 ( .A1(n746), .A2(n745), .ZN(n748) );
  XNOR2_X1 U821 ( .A(G1986), .B(G290), .ZN(n1030) );
  NAND2_X1 U822 ( .A1(n1030), .A2(n760), .ZN(n747) );
  NAND2_X1 U823 ( .A1(n748), .A2(n747), .ZN(n763) );
  NOR2_X1 U824 ( .A1(G1996), .A2(n895), .ZN(n933) );
  INV_X1 U825 ( .A(n749), .ZN(n752) );
  NOR2_X1 U826 ( .A1(G1991), .A2(n910), .ZN(n949) );
  NOR2_X1 U827 ( .A1(G1986), .A2(G290), .ZN(n750) );
  NOR2_X1 U828 ( .A1(n949), .A2(n750), .ZN(n751) );
  NOR2_X1 U829 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U830 ( .A1(n933), .A2(n753), .ZN(n754) );
  XNOR2_X1 U831 ( .A(n754), .B(KEYINPUT39), .ZN(n756) );
  NAND2_X1 U832 ( .A1(n756), .A2(n755), .ZN(n759) );
  NOR2_X1 U833 ( .A1(n913), .A2(n757), .ZN(n758) );
  XNOR2_X1 U834 ( .A(KEYINPUT103), .B(n758), .ZN(n937) );
  NAND2_X1 U835 ( .A1(n759), .A2(n937), .ZN(n761) );
  NAND2_X1 U836 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U837 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U838 ( .A(n764), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U839 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U840 ( .A(G2446), .B(G2430), .Z(n766) );
  XNOR2_X1 U841 ( .A(G2451), .B(KEYINPUT104), .ZN(n765) );
  XNOR2_X1 U842 ( .A(n766), .B(n765), .ZN(n767) );
  XOR2_X1 U843 ( .A(n767), .B(G2427), .Z(n769) );
  XNOR2_X1 U844 ( .A(G1348), .B(G1341), .ZN(n768) );
  XNOR2_X1 U845 ( .A(n769), .B(n768), .ZN(n773) );
  XOR2_X1 U846 ( .A(G2443), .B(G2435), .Z(n771) );
  XNOR2_X1 U847 ( .A(G2438), .B(G2454), .ZN(n770) );
  XNOR2_X1 U848 ( .A(n771), .B(n770), .ZN(n772) );
  XOR2_X1 U849 ( .A(n773), .B(n772), .Z(n774) );
  AND2_X1 U850 ( .A1(G14), .A2(n774), .ZN(G401) );
  AND2_X1 U851 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U852 ( .A(n1024), .ZN(G299) );
  INV_X1 U853 ( .A(G132), .ZN(G219) );
  INV_X1 U854 ( .A(G82), .ZN(G220) );
  INV_X1 U855 ( .A(G57), .ZN(G237) );
  NAND2_X1 U856 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U857 ( .A1(n778), .A2(n777), .ZN(G160) );
  NAND2_X1 U858 ( .A1(G7), .A2(G661), .ZN(n779) );
  XNOR2_X1 U859 ( .A(n779), .B(KEYINPUT68), .ZN(n780) );
  XOR2_X1 U860 ( .A(KEYINPUT10), .B(n780), .Z(n931) );
  NAND2_X1 U861 ( .A1(n931), .A2(G567), .ZN(n781) );
  XOR2_X1 U862 ( .A(KEYINPUT11), .B(n781), .Z(G234) );
  NAND2_X1 U863 ( .A1(n1020), .A2(G860), .ZN(G153) );
  NAND2_X1 U864 ( .A1(G868), .A2(G301), .ZN(n783) );
  INV_X1 U865 ( .A(G868), .ZN(n823) );
  NAND2_X1 U866 ( .A1(n916), .A2(n823), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n783), .A2(n782), .ZN(G284) );
  NAND2_X1 U868 ( .A1(G868), .A2(G286), .ZN(n785) );
  NAND2_X1 U869 ( .A1(G299), .A2(n823), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n785), .A2(n784), .ZN(G297) );
  INV_X1 U871 ( .A(G559), .ZN(n789) );
  NOR2_X1 U872 ( .A1(G860), .A2(n789), .ZN(n786) );
  XNOR2_X1 U873 ( .A(KEYINPUT71), .B(n786), .ZN(n787) );
  INV_X1 U874 ( .A(n916), .ZN(n1008) );
  NAND2_X1 U875 ( .A1(n787), .A2(n1008), .ZN(n788) );
  XNOR2_X1 U876 ( .A(n788), .B(KEYINPUT16), .ZN(G148) );
  AND2_X1 U877 ( .A1(n823), .A2(n1020), .ZN(n792) );
  NAND2_X1 U878 ( .A1(G868), .A2(n789), .ZN(n790) );
  NOR2_X1 U879 ( .A1(n790), .A2(n916), .ZN(n791) );
  NOR2_X1 U880 ( .A1(n792), .A2(n791), .ZN(G282) );
  NAND2_X1 U881 ( .A1(G123), .A2(n903), .ZN(n793) );
  XNOR2_X1 U882 ( .A(n793), .B(KEYINPUT18), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G111), .A2(n904), .ZN(n794) );
  XOR2_X1 U884 ( .A(KEYINPUT73), .B(n794), .Z(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n801) );
  NAND2_X1 U886 ( .A1(n899), .A2(G135), .ZN(n797) );
  XNOR2_X1 U887 ( .A(n797), .B(KEYINPUT72), .ZN(n799) );
  NAND2_X1 U888 ( .A1(G99), .A2(n900), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U890 ( .A1(n801), .A2(n800), .ZN(n946) );
  XNOR2_X1 U891 ( .A(G2096), .B(n946), .ZN(n802) );
  INV_X1 U892 ( .A(G2100), .ZN(n864) );
  NAND2_X1 U893 ( .A1(n802), .A2(n864), .ZN(G156) );
  XOR2_X1 U894 ( .A(n1020), .B(KEYINPUT74), .Z(n804) );
  NAND2_X1 U895 ( .A1(G559), .A2(n1008), .ZN(n803) );
  XNOR2_X1 U896 ( .A(n804), .B(n803), .ZN(n821) );
  NOR2_X1 U897 ( .A1(G860), .A2(n821), .ZN(n815) );
  NAND2_X1 U898 ( .A1(G67), .A2(n805), .ZN(n808) );
  NAND2_X1 U899 ( .A1(G55), .A2(n806), .ZN(n807) );
  NAND2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n814) );
  NAND2_X1 U901 ( .A1(G93), .A2(n809), .ZN(n812) );
  NAND2_X1 U902 ( .A1(G80), .A2(n810), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n812), .A2(n811), .ZN(n813) );
  OR2_X1 U904 ( .A1(n814), .A2(n813), .ZN(n824) );
  XOR2_X1 U905 ( .A(n815), .B(n824), .Z(G145) );
  INV_X1 U906 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U907 ( .A(KEYINPUT19), .B(G288), .ZN(n820) );
  XOR2_X1 U908 ( .A(n824), .B(G305), .Z(n816) );
  XOR2_X1 U909 ( .A(n816), .B(G166), .Z(n817) );
  XOR2_X1 U910 ( .A(G299), .B(n817), .Z(n818) );
  XNOR2_X1 U911 ( .A(n818), .B(G290), .ZN(n819) );
  XNOR2_X1 U912 ( .A(n820), .B(n819), .ZN(n917) );
  XOR2_X1 U913 ( .A(n917), .B(n821), .Z(n822) );
  NOR2_X1 U914 ( .A1(n823), .A2(n822), .ZN(n826) );
  NOR2_X1 U915 ( .A1(G868), .A2(n824), .ZN(n825) );
  NOR2_X1 U916 ( .A1(n826), .A2(n825), .ZN(G295) );
  NAND2_X1 U917 ( .A1(G2078), .A2(G2084), .ZN(n827) );
  XOR2_X1 U918 ( .A(KEYINPUT20), .B(n827), .Z(n828) );
  NAND2_X1 U919 ( .A1(n828), .A2(G2090), .ZN(n829) );
  XNOR2_X1 U920 ( .A(n829), .B(KEYINPUT76), .ZN(n830) );
  XNOR2_X1 U921 ( .A(KEYINPUT21), .B(n830), .ZN(n831) );
  NAND2_X1 U922 ( .A1(G2072), .A2(n831), .ZN(G158) );
  NAND2_X1 U923 ( .A1(G120), .A2(G108), .ZN(n832) );
  NOR2_X1 U924 ( .A1(G237), .A2(n832), .ZN(n833) );
  NAND2_X1 U925 ( .A1(G69), .A2(n833), .ZN(n849) );
  NAND2_X1 U926 ( .A1(G567), .A2(n849), .ZN(n834) );
  XNOR2_X1 U927 ( .A(n834), .B(KEYINPUT77), .ZN(n839) );
  NOR2_X1 U928 ( .A1(G220), .A2(G219), .ZN(n835) );
  XNOR2_X1 U929 ( .A(KEYINPUT22), .B(n835), .ZN(n836) );
  NAND2_X1 U930 ( .A1(n836), .A2(G96), .ZN(n837) );
  OR2_X1 U931 ( .A1(G218), .A2(n837), .ZN(n850) );
  AND2_X1 U932 ( .A1(G2106), .A2(n850), .ZN(n838) );
  NOR2_X1 U933 ( .A1(n839), .A2(n838), .ZN(G319) );
  NAND2_X1 U934 ( .A1(G661), .A2(G483), .ZN(n841) );
  INV_X1 U935 ( .A(G319), .ZN(n840) );
  NOR2_X1 U936 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U937 ( .A(n842), .B(KEYINPUT78), .ZN(n847) );
  NAND2_X1 U938 ( .A1(G36), .A2(n847), .ZN(G176) );
  NAND2_X1 U939 ( .A1(G2106), .A2(n931), .ZN(G217) );
  NAND2_X1 U940 ( .A1(G15), .A2(G2), .ZN(n844) );
  INV_X1 U941 ( .A(G661), .ZN(n843) );
  NOR2_X1 U942 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n845), .B(KEYINPUT105), .ZN(G259) );
  NAND2_X1 U944 ( .A1(G3), .A2(G1), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n846), .B(KEYINPUT106), .ZN(n848) );
  NAND2_X1 U946 ( .A1(n848), .A2(n847), .ZN(G188) );
  XNOR2_X1 U947 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U949 ( .A(G120), .ZN(G236) );
  INV_X1 U950 ( .A(G96), .ZN(G221) );
  NOR2_X1 U951 ( .A1(n850), .A2(n849), .ZN(G325) );
  INV_X1 U952 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U953 ( .A(G1956), .B(KEYINPUT41), .ZN(n860) );
  XOR2_X1 U954 ( .A(G1976), .B(G1961), .Z(n852) );
  XNOR2_X1 U955 ( .A(G1986), .B(G1971), .ZN(n851) );
  XNOR2_X1 U956 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U957 ( .A(G1966), .B(G1981), .Z(n854) );
  XNOR2_X1 U958 ( .A(G1996), .B(G1991), .ZN(n853) );
  XNOR2_X1 U959 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U960 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U961 ( .A(KEYINPUT110), .B(G2474), .ZN(n857) );
  XNOR2_X1 U962 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(G229) );
  XNOR2_X1 U964 ( .A(G2067), .B(G2084), .ZN(n861) );
  XNOR2_X1 U965 ( .A(n861), .B(KEYINPUT42), .ZN(n872) );
  XOR2_X1 U966 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n863) );
  XNOR2_X1 U967 ( .A(G2678), .B(G2096), .ZN(n862) );
  XNOR2_X1 U968 ( .A(n863), .B(n862), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n864), .B(G2078), .ZN(n866) );
  XNOR2_X1 U970 ( .A(G2090), .B(G2072), .ZN(n865) );
  XNOR2_X1 U971 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U972 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U973 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n869) );
  XNOR2_X1 U974 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U975 ( .A(n872), .B(n871), .ZN(G227) );
  NAND2_X1 U976 ( .A1(G124), .A2(n903), .ZN(n873) );
  XNOR2_X1 U977 ( .A(n873), .B(KEYINPUT44), .ZN(n876) );
  NAND2_X1 U978 ( .A1(G112), .A2(n904), .ZN(n874) );
  XOR2_X1 U979 ( .A(KEYINPUT111), .B(n874), .Z(n875) );
  NAND2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G136), .A2(n899), .ZN(n878) );
  NAND2_X1 U982 ( .A1(G100), .A2(n900), .ZN(n877) );
  NAND2_X1 U983 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U984 ( .A1(n880), .A2(n879), .ZN(G162) );
  NAND2_X1 U985 ( .A1(G118), .A2(n904), .ZN(n889) );
  XNOR2_X1 U986 ( .A(KEYINPUT113), .B(KEYINPUT45), .ZN(n884) );
  NAND2_X1 U987 ( .A1(G142), .A2(n899), .ZN(n882) );
  NAND2_X1 U988 ( .A1(G106), .A2(n900), .ZN(n881) );
  NAND2_X1 U989 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U990 ( .A(n884), .B(n883), .ZN(n887) );
  NAND2_X1 U991 ( .A1(n903), .A2(G130), .ZN(n885) );
  XOR2_X1 U992 ( .A(KEYINPUT112), .B(n885), .Z(n886) );
  NOR2_X1 U993 ( .A1(n887), .A2(n886), .ZN(n888) );
  NAND2_X1 U994 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U995 ( .A(n890), .B(G162), .ZN(n894) );
  XOR2_X1 U996 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n892) );
  XNOR2_X1 U997 ( .A(G160), .B(KEYINPUT114), .ZN(n891) );
  XNOR2_X1 U998 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U999 ( .A(n894), .B(n893), .Z(n897) );
  XOR2_X1 U1000 ( .A(G164), .B(n895), .Z(n896) );
  XNOR2_X1 U1001 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U1002 ( .A(n898), .B(n946), .Z(n912) );
  NAND2_X1 U1003 ( .A1(G139), .A2(n899), .ZN(n902) );
  NAND2_X1 U1004 ( .A1(G103), .A2(n900), .ZN(n901) );
  NAND2_X1 U1005 ( .A1(n902), .A2(n901), .ZN(n909) );
  NAND2_X1 U1006 ( .A1(G127), .A2(n903), .ZN(n906) );
  NAND2_X1 U1007 ( .A1(G115), .A2(n904), .ZN(n905) );
  NAND2_X1 U1008 ( .A1(n906), .A2(n905), .ZN(n907) );
  XOR2_X1 U1009 ( .A(KEYINPUT47), .B(n907), .Z(n908) );
  NOR2_X1 U1010 ( .A1(n909), .A2(n908), .ZN(n939) );
  XNOR2_X1 U1011 ( .A(n910), .B(n939), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(n912), .B(n911), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n915), .ZN(G395) );
  XOR2_X1 U1015 ( .A(n916), .B(n1020), .Z(n918) );
  XNOR2_X1 U1016 ( .A(n918), .B(n917), .ZN(n919) );
  XOR2_X1 U1017 ( .A(n919), .B(KEYINPUT116), .Z(n921) );
  XOR2_X1 U1018 ( .A(G301), .B(KEYINPUT115), .Z(n920) );
  XNOR2_X1 U1019 ( .A(n921), .B(n920), .ZN(n922) );
  XOR2_X1 U1020 ( .A(n922), .B(G286), .Z(n923) );
  NOR2_X1 U1021 ( .A1(G37), .A2(n923), .ZN(G397) );
  NOR2_X1 U1022 ( .A1(G229), .A2(G227), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(KEYINPUT49), .B(KEYINPUT117), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(n925), .B(n924), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n926), .A2(G319), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(G401), .A2(n927), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(KEYINPUT118), .B(n928), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(G395), .A2(G397), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(G225) );
  INV_X1 U1030 ( .A(G225), .ZN(G308) );
  INV_X1 U1031 ( .A(G69), .ZN(G235) );
  INV_X1 U1032 ( .A(n931), .ZN(G223) );
  XOR2_X1 U1033 ( .A(G2090), .B(G162), .Z(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1035 ( .A(n934), .B(KEYINPUT51), .ZN(n935) );
  NOR2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n938) );
  NAND2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n945) );
  XOR2_X1 U1038 ( .A(G2072), .B(n939), .Z(n941) );
  XOR2_X1 U1039 ( .A(G164), .B(G2078), .Z(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1041 ( .A(KEYINPUT50), .B(n942), .Z(n943) );
  XNOR2_X1 U1042 ( .A(KEYINPUT120), .B(n943), .ZN(n944) );
  NOR2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n955) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n951) );
  XOR2_X1 U1045 ( .A(G160), .B(G2084), .Z(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(KEYINPUT52), .B(n956), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(KEYINPUT121), .B(n957), .ZN(n958) );
  INV_X1 U1052 ( .A(KEYINPUT55), .ZN(n1004) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n1004), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n959), .A2(G29), .ZN(n1040) );
  XOR2_X1 U1055 ( .A(G25), .B(G1991), .Z(n960) );
  NAND2_X1 U1056 ( .A1(n960), .A2(G28), .ZN(n969) );
  XNOR2_X1 U1057 ( .A(G2067), .B(G26), .ZN(n962) );
  XNOR2_X1 U1058 ( .A(G33), .B(G2072), .ZN(n961) );
  NOR2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G1996), .B(G32), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(G27), .B(n963), .ZN(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(n970), .B(KEYINPUT123), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(n971), .B(KEYINPUT53), .ZN(n974) );
  XOR2_X1 U1067 ( .A(G2084), .B(G34), .Z(n972) );
  XNOR2_X1 U1068 ( .A(KEYINPUT54), .B(n972), .ZN(n973) );
  NAND2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(KEYINPUT122), .B(G2090), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(G35), .B(n975), .ZN(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1073 ( .A(KEYINPUT124), .B(n978), .Z(n1003) );
  OR2_X1 U1074 ( .A1(n1004), .A2(n1003), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(G11), .A2(n979), .ZN(n1038) );
  XNOR2_X1 U1076 ( .A(G20), .B(n980), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(G1981), .B(G6), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(G1341), .B(G19), .ZN(n981) );
  NOR2_X1 U1079 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n987) );
  XOR2_X1 U1081 ( .A(KEYINPUT59), .B(G1348), .Z(n985) );
  XNOR2_X1 U1082 ( .A(G4), .B(n985), .ZN(n986) );
  NOR2_X1 U1083 ( .A1(n987), .A2(n986), .ZN(n989) );
  XOR2_X1 U1084 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n988) );
  XNOR2_X1 U1085 ( .A(n989), .B(n988), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(G1961), .B(G5), .ZN(n991) );
  XNOR2_X1 U1087 ( .A(G1966), .B(G21), .ZN(n990) );
  NOR2_X1 U1088 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1089 ( .A1(n993), .A2(n992), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(G1971), .B(G22), .ZN(n995) );
  XNOR2_X1 U1091 ( .A(G23), .B(G1976), .ZN(n994) );
  NOR2_X1 U1092 ( .A1(n995), .A2(n994), .ZN(n997) );
  XOR2_X1 U1093 ( .A(G1986), .B(G24), .Z(n996) );
  NAND2_X1 U1094 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1095 ( .A(KEYINPUT58), .B(n998), .ZN(n999) );
  NOR2_X1 U1096 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1097 ( .A(KEYINPUT61), .B(n1001), .Z(n1002) );
  NOR2_X1 U1098 ( .A1(G16), .A2(n1002), .ZN(n1007) );
  NAND2_X1 U1099 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1100 ( .A1(G29), .A2(n1005), .ZN(n1006) );
  NOR2_X1 U1101 ( .A1(n1007), .A2(n1006), .ZN(n1036) );
  XNOR2_X1 U1102 ( .A(G16), .B(KEYINPUT56), .ZN(n1034) );
  XOR2_X1 U1103 ( .A(G301), .B(G1961), .Z(n1011) );
  XNOR2_X1 U1104 ( .A(G1348), .B(KEYINPUT125), .ZN(n1009) );
  XOR2_X1 U1105 ( .A(n1009), .B(n1008), .Z(n1010) );
  NAND2_X1 U1106 ( .A1(n1011), .A2(n1010), .ZN(n1019) );
  XOR2_X1 U1107 ( .A(G1971), .B(G303), .Z(n1012) );
  XNOR2_X1 U1108 ( .A(n1012), .B(KEYINPUT126), .ZN(n1017) );
  XOR2_X1 U1109 ( .A(G1966), .B(G168), .Z(n1013) );
  NOR2_X1 U1110 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1111 ( .A(KEYINPUT57), .B(n1015), .Z(n1016) );
  NAND2_X1 U1112 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1113 ( .A1(n1019), .A2(n1018), .ZN(n1032) );
  XNOR2_X1 U1114 ( .A(n1020), .B(G1341), .ZN(n1028) );
  INV_X1 U1115 ( .A(n1021), .ZN(n1022) );
  NAND2_X1 U1116 ( .A1(n1023), .A2(n1022), .ZN(n1026) );
  XOR2_X1 U1117 ( .A(G1956), .B(n1024), .Z(n1025) );
  NOR2_X1 U1118 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1119 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1120 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1121 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1122 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1123 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NOR2_X1 U1124 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1125 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNOR2_X1 U1126 ( .A(KEYINPUT62), .B(n1041), .ZN(G150) );
  INV_X1 U1127 ( .A(G150), .ZN(G311) );
endmodule

