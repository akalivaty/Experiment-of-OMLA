//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n550, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n591, new_n592, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1145, new_n1146, new_n1147;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT67), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT68), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT69), .Z(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT71), .B1(new_n469), .B2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(new_n465), .A3(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G101), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g050(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g053(.A(KEYINPUT70), .B(G125), .C1(new_n466), .C2(new_n467), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n475), .B1(new_n481), .B2(G2105), .ZN(G160));
  NOR2_X1   g057(.A1(new_n466), .A2(new_n467), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(new_n465), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  AND2_X1   g060(.A1(G112), .A2(G2105), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(G100), .B2(new_n465), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n469), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n483), .A2(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(G136), .B2(new_n489), .ZN(G162));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(new_n469), .ZN(new_n493));
  NAND2_X1  g068(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(G2105), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(KEYINPUT72), .A2(KEYINPUT4), .A3(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n493), .B2(new_n494), .ZN(new_n499));
  NAND2_X1  g074(.A1(G102), .A2(G2104), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n465), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(G138), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n497), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT73), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n516), .A2(new_n522), .ZN(G166));
  AND2_X1   g098(.A1(new_n513), .A2(new_n517), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n517), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n525), .A2(new_n527), .A3(new_n529), .A4(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  AOI22_X1  g107(.A1(new_n524), .A2(G90), .B1(new_n528), .B2(G52), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n515), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n535), .A2(new_n536), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n533), .B1(new_n538), .B2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n515), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n518), .A2(new_n544), .B1(new_n520), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(new_n550));
  XOR2_X1   g125(.A(new_n550), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(G188));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G53), .ZN(new_n556));
  OR3_X1    g131(.A1(new_n520), .A2(KEYINPUT9), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n520), .B2(new_n556), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n515), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n524), .A2(G91), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n559), .A2(new_n561), .A3(new_n562), .ZN(G299));
  INV_X1    g138(.A(G166), .ZN(G303));
  NAND2_X1  g139(.A1(new_n524), .A2(G87), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n528), .A2(G49), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(G288));
  AOI22_X1  g143(.A1(new_n524), .A2(G86), .B1(new_n528), .B2(G48), .ZN(new_n569));
  INV_X1    g144(.A(G61), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n510), .B2(new_n512), .ZN(new_n571));
  AND2_X1   g146(.A1(G73), .A2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(G305));
  AOI22_X1  g149(.A1(new_n524), .A2(G85), .B1(new_n528), .B2(G47), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n515), .B2(new_n576), .ZN(G290));
  NAND2_X1  g152(.A1(new_n524), .A2(G92), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT10), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n578), .B(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(new_n515), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n528), .A2(KEYINPUT77), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n528), .A2(KEYINPUT77), .ZN(new_n585));
  OAI21_X1  g160(.A(G54), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n580), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  MUX2_X1   g163(.A(G301), .B(new_n587), .S(new_n588), .Z(G284));
  MUX2_X1   g164(.A(G301), .B(new_n587), .S(new_n588), .Z(G321));
  NOR2_X1   g165(.A1(G286), .A2(new_n588), .ZN(new_n591));
  INV_X1    g166(.A(G299), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(new_n588), .ZN(G297));
  XNOR2_X1  g168(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g169(.A(new_n587), .ZN(new_n595));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G860), .ZN(G148));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G868), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n547), .A2(G868), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(KEYINPUT79), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(KEYINPUT79), .B2(new_n599), .ZN(G323));
  XNOR2_X1  g177(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g178(.A1(new_n470), .A2(new_n472), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n493), .A2(new_n494), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  INV_X1    g183(.A(G2100), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  MUX2_X1   g186(.A(G99), .B(G111), .S(G2105), .Z(new_n612));
  AOI22_X1  g187(.A1(new_n484), .A2(G123), .B1(G2104), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G135), .ZN(new_n614));
  INV_X1    g189(.A(new_n489), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(G2096), .Z(new_n617));
  NAND3_X1  g192(.A1(new_n610), .A2(new_n611), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT80), .ZN(G156));
  XOR2_X1   g194(.A(KEYINPUT15), .B(G2435), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2438), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n621), .A2(G2427), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(G2427), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G2430), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n622), .A2(G2430), .A3(new_n623), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n626), .A2(KEYINPUT14), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2451), .B(G2454), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n628), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT81), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n633), .A2(new_n634), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(G14), .A3(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT82), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT83), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n646), .A2(KEYINPUT17), .A3(new_n647), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n646), .B1(KEYINPUT17), .B2(new_n647), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(KEYINPUT84), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n645), .A2(new_n653), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n647), .B1(new_n655), .B2(KEYINPUT17), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n650), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2096), .B(G2100), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT85), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(G227));
  XNOR2_X1  g235(.A(G1956), .B(G2474), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT87), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1961), .B(G1966), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT20), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n662), .A2(new_n663), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n670), .A2(new_n667), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT88), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n664), .A2(new_n667), .A3(new_n670), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n676), .B(new_n679), .ZN(G229));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G32), .ZN(new_n682));
  NAND3_X1  g257(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT26), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n604), .A2(G105), .ZN(new_n685));
  AOI211_X1 g260(.A(new_n684), .B(new_n685), .C1(G129), .C2(new_n484), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n489), .A2(G141), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT97), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n682), .B1(new_n690), .B2(new_n681), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT27), .B(G1996), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G2078), .ZN(new_n694));
  NAND2_X1  g269(.A1(G164), .A2(G29), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G27), .B2(G29), .ZN(new_n696));
  AOI22_X1  g271(.A1(new_n691), .A2(new_n693), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(new_n694), .B2(new_n696), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT31), .B(G11), .Z(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT30), .B(G28), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n699), .B1(new_n681), .B2(new_n700), .ZN(new_n701));
  OAI221_X1 g276(.A(new_n701), .B1(new_n681), .B2(new_n616), .C1(new_n691), .C2(new_n693), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT95), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT25), .ZN(new_n705));
  NAND2_X1  g280(.A1(G115), .A2(G2104), .ZN(new_n706));
  INV_X1    g281(.A(G127), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n483), .B2(new_n707), .ZN(new_n708));
  AOI22_X1  g283(.A1(new_n708), .A2(G2105), .B1(new_n489), .B2(G139), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(G33), .B(new_n710), .S(G29), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G2072), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n698), .A2(new_n702), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT98), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G16), .B2(G21), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NOR2_X1   g291(.A1(G286), .A2(new_n716), .ZN(new_n717));
  MUX2_X1   g292(.A(new_n715), .B(new_n714), .S(new_n717), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT99), .ZN(new_n719));
  INV_X1    g294(.A(G1966), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n716), .A2(G5), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G171), .B2(new_n716), .ZN(new_n723));
  INV_X1    g298(.A(G1961), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(G160), .A2(G29), .ZN(new_n726));
  AND2_X1   g301(.A1(KEYINPUT24), .A2(G34), .ZN(new_n727));
  NOR2_X1   g302(.A1(KEYINPUT24), .A2(G34), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n681), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT96), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(G2084), .Z(new_n732));
  AND4_X1   g307(.A1(new_n713), .A2(new_n721), .A3(new_n725), .A4(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT100), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NOR2_X1   g311(.A1(G29), .A2(G35), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G162), .B2(G29), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT29), .Z(new_n739));
  INV_X1    g314(.A(G2090), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n595), .A2(G16), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G4), .B2(G16), .ZN(new_n742));
  INV_X1    g317(.A(G1348), .ZN(new_n743));
  OAI22_X1  g318(.A1(new_n739), .A2(new_n740), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n716), .A2(G20), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT23), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n592), .B2(new_n716), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(G1956), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n742), .B2(new_n743), .ZN(new_n749));
  NOR2_X1   g324(.A1(G16), .A2(G19), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n547), .B2(G16), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1341), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G1956), .B2(new_n747), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n681), .A2(G26), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT93), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT28), .ZN(new_n756));
  MUX2_X1   g331(.A(G104), .B(G116), .S(G2105), .Z(new_n757));
  AOI22_X1  g332(.A1(new_n484), .A2(G128), .B1(G2104), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G140), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n615), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G29), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n761), .A2(KEYINPUT92), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(KEYINPUT92), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n756), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT94), .B(G2067), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n749), .A2(new_n753), .A3(new_n766), .ZN(new_n767));
  AOI211_X1 g342(.A(new_n744), .B(new_n767), .C1(new_n740), .C2(new_n739), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n735), .A2(new_n736), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G6), .A2(G16), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n569), .A2(new_n573), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(G16), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT89), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT90), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT32), .B(G1981), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G23), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT91), .Z(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G288), .B2(new_n716), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT33), .B(G1976), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n780), .B(new_n781), .Z(new_n782));
  NOR2_X1   g357(.A1(G16), .A2(G22), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G166), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1971), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n776), .A2(new_n777), .A3(new_n782), .A4(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT34), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(KEYINPUT34), .ZN(new_n789));
  MUX2_X1   g364(.A(G95), .B(G107), .S(G2105), .Z(new_n790));
  AOI22_X1  g365(.A1(new_n484), .A2(G119), .B1(G2104), .B2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G131), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n615), .ZN(new_n793));
  MUX2_X1   g368(.A(G25), .B(new_n793), .S(G29), .Z(new_n794));
  XOR2_X1   g369(.A(KEYINPUT35), .B(G1991), .Z(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n794), .B(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G24), .B(G290), .S(G16), .Z(new_n798));
  AND2_X1   g373(.A1(new_n798), .A2(G1986), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(G1986), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n797), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n788), .A2(new_n789), .A3(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT36), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(KEYINPUT36), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n769), .B1(new_n803), .B2(new_n804), .ZN(G311));
  INV_X1    g380(.A(G311), .ZN(G150));
  AOI22_X1  g381(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(new_n515), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n524), .A2(G93), .B1(new_n528), .B2(G55), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G860), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT37), .Z(new_n812));
  INV_X1    g387(.A(new_n547), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(new_n810), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n547), .A2(new_n808), .A3(new_n809), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT38), .Z(new_n817));
  NOR2_X1   g392(.A1(new_n587), .A2(new_n596), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n821));
  INV_X1    g396(.A(G860), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n820), .B2(KEYINPUT39), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n812), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT101), .ZN(G145));
  XNOR2_X1  g400(.A(new_n760), .B(G164), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  OAI22_X1  g402(.A1(new_n827), .A2(new_n690), .B1(KEYINPUT102), .B2(new_n710), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n690), .B2(new_n827), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n607), .B(new_n793), .ZN(new_n830));
  MUX2_X1   g405(.A(G106), .B(G118), .S(G2105), .Z(new_n831));
  AOI22_X1  g406(.A1(new_n484), .A2(G130), .B1(G2104), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G142), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n615), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n830), .B(new_n834), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n829), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n710), .A2(KEYINPUT102), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  XOR2_X1   g414(.A(G162), .B(G160), .Z(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(new_n616), .Z(new_n841));
  OR3_X1    g416(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G37), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n841), .B1(new_n838), .B2(new_n839), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g421(.A1(new_n810), .A2(new_n588), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n587), .B(G299), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(KEYINPUT41), .ZN(new_n850));
  INV_X1    g425(.A(new_n816), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n598), .B(new_n851), .ZN(new_n852));
  MUX2_X1   g427(.A(new_n849), .B(new_n850), .S(new_n852), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n771), .B(G166), .ZN(new_n854));
  XNOR2_X1  g429(.A(G290), .B(G288), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n854), .B(new_n855), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT42), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n853), .A2(new_n857), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n858), .B1(new_n859), .B2(KEYINPUT103), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(KEYINPUT103), .B2(new_n859), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n847), .B1(new_n861), .B2(new_n588), .ZN(G295));
  OAI21_X1  g437(.A(new_n847), .B1(new_n861), .B2(new_n588), .ZN(G331));
  XNOR2_X1  g438(.A(G301), .B(G286), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n816), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n865), .A2(KEYINPUT106), .ZN(new_n866));
  XNOR2_X1  g441(.A(G301), .B(G168), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n851), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n868), .A3(KEYINPUT106), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n850), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n864), .A2(KEYINPUT105), .A3(new_n816), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n873), .A3(new_n868), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n870), .B1(new_n848), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n856), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n850), .ZN(new_n877));
  INV_X1    g452(.A(new_n856), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n866), .A2(new_n869), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n877), .B(new_n878), .C1(new_n879), .C2(new_n848), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(new_n843), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT43), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n877), .B1(new_n879), .B2(new_n848), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n856), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(new_n843), .A3(new_n880), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n882), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n881), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n884), .A2(KEYINPUT43), .A3(new_n843), .A4(new_n880), .ZN(new_n889));
  XOR2_X1   g464(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT107), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT107), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n886), .A2(new_n895), .A3(new_n892), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(G397));
  INV_X1    g472(.A(G40), .ZN(new_n898));
  AOI211_X1 g473(.A(new_n898), .B(new_n475), .C1(new_n481), .C2(G2105), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT45), .ZN(new_n900));
  INV_X1    g475(.A(G1384), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n506), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(G1996), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n904), .A2(KEYINPUT46), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(KEYINPUT46), .ZN(new_n906));
  INV_X1    g481(.A(new_n903), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n760), .B(G2067), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n907), .B1(new_n908), .B2(new_n689), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n904), .A2(new_n690), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT108), .ZN(new_n914));
  INV_X1    g489(.A(G1996), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n907), .B1(new_n916), .B2(new_n908), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n793), .B(new_n795), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n918), .B1(new_n903), .B2(new_n919), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n903), .A2(G1986), .A3(G290), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT48), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n912), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n793), .A2(new_n796), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n918), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n760), .A2(G2067), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n903), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT126), .ZN(new_n929));
  XNOR2_X1  g504(.A(G290), .B(G1986), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n920), .B1(new_n907), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(G8), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n902), .A2(new_n900), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n901), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n899), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n720), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT50), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(new_n506), .B2(new_n901), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n479), .A2(new_n480), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT70), .B1(new_n605), .B2(G125), .ZN(new_n940));
  OAI21_X1  g515(.A(G2105), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n475), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(G40), .A3(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n938), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n506), .A2(new_n937), .A3(new_n901), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n506), .A2(KEYINPUT109), .A3(new_n937), .A4(new_n901), .ZN(new_n948));
  XNOR2_X1  g523(.A(KEYINPUT116), .B(G2084), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n944), .A2(new_n947), .A3(new_n948), .A4(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n932), .B1(new_n936), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT124), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT51), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n936), .A2(new_n951), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(G8), .ZN(new_n956));
  NOR2_X1   g531(.A1(G168), .A2(new_n932), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n956), .A2(new_n953), .A3(KEYINPUT51), .A4(new_n958), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n952), .A2(G286), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT62), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G1981), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n569), .A2(KEYINPUT113), .A3(new_n965), .A4(new_n573), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n528), .A2(G48), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n513), .A2(G86), .A3(new_n517), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n967), .A2(new_n573), .A3(new_n965), .A4(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(G305), .A2(G1981), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT49), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(G8), .B1(new_n943), .B2(new_n902), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT111), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n979), .B(G8), .C1(new_n943), .C2(new_n902), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n972), .A2(KEYINPUT49), .A3(new_n973), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n976), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G288), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n978), .A2(new_n980), .B1(G1976), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(KEYINPUT112), .ZN(new_n987));
  NOR2_X1   g562(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n985), .A2(new_n987), .B1(G288), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n984), .A2(G1976), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n981), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n987), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n983), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n902), .A2(KEYINPUT50), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n995), .A2(new_n899), .A3(new_n948), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n996), .A2(KEYINPUT110), .A3(new_n740), .A4(new_n947), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n944), .A2(new_n740), .A3(new_n947), .A4(new_n948), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n935), .A2(new_n785), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(G303), .A2(G8), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT55), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(G8), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n945), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n506), .A2(KEYINPUT115), .A3(new_n937), .A4(new_n901), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n944), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1001), .B1(new_n1010), .B2(G2090), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G8), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n1004), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n994), .A2(new_n1006), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n933), .A2(new_n694), .A3(new_n899), .A4(new_n934), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT53), .ZN(new_n1017));
  AND3_X1   g592(.A1(KEYINPUT72), .A2(KEYINPUT4), .A3(G138), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n466), .B2(new_n467), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n500), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n1020), .A2(new_n465), .B1(new_n504), .B2(new_n503), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n1021), .B2(new_n497), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n899), .B(new_n948), .C1(new_n937), .C2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT109), .B1(new_n1022), .B2(new_n937), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT120), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT120), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n944), .A2(new_n1026), .A3(new_n947), .A4(new_n948), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(new_n724), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(G301), .B1(new_n1017), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n954), .A2(new_n959), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT62), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n961), .A4(new_n962), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n964), .A2(new_n1015), .A3(new_n1029), .A4(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n976), .A2(new_n981), .A3(new_n982), .ZN(new_n1034));
  INV_X1    g609(.A(new_n980), .ZN(new_n1035));
  NAND4_X1  g610(.A1(G160), .A2(G40), .A3(new_n901), .A4(new_n506), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n979), .B1(new_n1036), .B2(G8), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n990), .B(new_n987), .C1(new_n1035), .C2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G288), .A2(new_n988), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n987), .B1(new_n981), .B2(new_n990), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1034), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(KEYINPUT114), .B(new_n1034), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1006), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OR3_X1    g621(.A1(new_n983), .A2(G1976), .A3(G288), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1047), .A2(new_n972), .B1(new_n980), .B2(new_n978), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1033), .A2(new_n1049), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n956), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1025), .A2(new_n743), .A3(new_n1027), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1036), .A2(G2067), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n587), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n1055));
  XNOR2_X1  g630(.A(G299), .B(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1956), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n995), .A2(new_n899), .A3(new_n1009), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1008), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT56), .B(G2072), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n933), .A2(new_n899), .A3(new_n934), .A4(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1056), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n933), .A2(new_n899), .A3(new_n934), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1057), .A2(new_n1010), .B1(new_n1065), .B2(new_n1061), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1066), .B2(new_n1056), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1060), .A2(new_n1056), .A3(new_n1064), .A4(new_n1062), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n1054), .A2(new_n1063), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1052), .A2(new_n587), .A3(new_n1053), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(new_n1054), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT60), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT58), .B(G1341), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1075), .B(KEYINPUT121), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n943), .B2(new_n902), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1036), .A2(KEYINPUT122), .A3(new_n1076), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n933), .A2(new_n915), .A3(new_n899), .A4(new_n934), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1079), .A2(new_n1081), .A3(new_n1080), .A4(KEYINPUT123), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1074), .B1(new_n1086), .B2(new_n547), .ZN(new_n1087));
  AOI211_X1 g662(.A(KEYINPUT59), .B(new_n813), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1072), .A2(new_n1073), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT61), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1063), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1060), .A2(new_n1056), .A3(new_n1062), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n587), .A2(KEYINPUT60), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1092), .A2(KEYINPUT119), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1063), .B1(new_n1097), .B2(new_n1068), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1093), .B(new_n1096), .C1(new_n1098), .C2(KEYINPUT61), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1070), .B1(new_n1089), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1030), .A2(new_n961), .A3(new_n962), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1029), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1017), .A2(new_n1028), .A3(G301), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(KEYINPUT54), .A3(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT125), .B(KEYINPUT54), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1103), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(new_n1029), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1101), .A2(new_n1104), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1051), .B1(new_n1100), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1050), .B1(new_n1110), .B2(new_n1014), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT63), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1002), .A2(new_n1114), .A3(G8), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1114), .B1(new_n1002), .B2(G8), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1004), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1113), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  AND4_X1   g697(.A1(G8), .A2(new_n1006), .A3(G168), .A4(new_n955), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1112), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n929), .B(new_n931), .C1(new_n1111), .C2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n813), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(new_n1074), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1063), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1090), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1092), .A2(new_n1091), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT60), .B1(new_n1071), .B2(new_n1054), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1128), .A2(new_n1131), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1108), .B1(new_n1134), .B2(new_n1070), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1015), .B1(new_n1135), .B2(new_n1051), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1113), .A2(new_n1120), .A3(new_n1117), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1120), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1123), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT63), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1136), .A2(new_n1140), .A3(new_n1050), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n929), .B1(new_n1141), .B2(new_n931), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n928), .B1(new_n1126), .B2(new_n1142), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g718(.A1(G229), .A2(new_n463), .A3(G227), .ZN(new_n1145));
  AND3_X1   g719(.A1(new_n642), .A2(new_n845), .A3(new_n1145), .ZN(new_n1146));
  AND2_X1   g720(.A1(new_n888), .A2(new_n889), .ZN(new_n1147));
  AND2_X1   g721(.A1(new_n1146), .A2(new_n1147), .ZN(G308));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(G225));
endmodule


