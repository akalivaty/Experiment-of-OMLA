//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1212, new_n1213,
    new_n1214, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT64), .B(G77), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  XOR2_X1   g0014(.A(KEYINPUT65), .B(G244), .Z(new_n215));
  AND2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G107), .A2(G264), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G20), .ZN(new_n225));
  INV_X1    g0025(.A(new_n201), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n212), .B1(KEYINPUT1), .B2(new_n222), .C1(new_n225), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G13), .ZN(new_n245));
  NOR3_X1   g0045(.A1(new_n245), .A2(new_n207), .A3(G1), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n223), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT66), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(new_n207), .B2(G1), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n206), .A2(KEYINPUT66), .A3(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(new_n202), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n250), .B1(new_n256), .B2(KEYINPUT67), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(KEYINPUT67), .B2(new_n256), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n203), .A2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(G150), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT8), .B(G58), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n259), .B1(new_n260), .B2(new_n262), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n267), .A2(new_n248), .B1(new_n202), .B2(new_n246), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n258), .A2(KEYINPUT9), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n273), .B1(G226), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G222), .A2(G1698), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G223), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n279), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n283), .B(new_n270), .C1(new_n214), .C2(new_n279), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G190), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(KEYINPUT9), .B1(new_n258), .B2(new_n268), .ZN(new_n289));
  NOR3_X1   g0089(.A1(new_n269), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT70), .ZN(new_n291));
  AOI21_X1  g0091(.A(KEYINPUT10), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n290), .B1(new_n293), .B2(new_n285), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(new_n294), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n286), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n258), .A2(new_n268), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n285), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n298), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n295), .A2(new_n296), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G58), .ZN(new_n304));
  INV_X1    g0104(.A(G68), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(G20), .B1(new_n306), .B2(new_n201), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n261), .A2(G159), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT7), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n263), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(new_n279), .B2(KEYINPUT71), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n311), .B1(new_n313), .B2(new_n207), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT71), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT71), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(new_n315), .A3(G33), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n318), .A2(new_n311), .A3(new_n207), .A4(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G68), .ZN(new_n322));
  OAI211_X1 g0122(.A(KEYINPUT16), .B(new_n310), .C1(new_n314), .C2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT16), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n311), .B1(new_n279), .B2(G20), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n316), .A2(new_n317), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n305), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n324), .B1(new_n328), .B2(new_n309), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n323), .A2(new_n248), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n273), .B1(G232), .B2(new_n277), .ZN(new_n331));
  INV_X1    g0131(.A(new_n270), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n318), .A2(new_n320), .ZN(new_n333));
  NOR2_X1   g0133(.A1(G223), .A2(G1698), .ZN(new_n334));
  INV_X1    g0134(.A(G226), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n334), .B1(new_n335), .B2(G1698), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n333), .A2(new_n336), .B1(G33), .B2(G87), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n331), .B1(new_n332), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G200), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n250), .A2(new_n255), .A3(new_n266), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n246), .B2(new_n266), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n331), .B(G190), .C1(new_n332), .C2(new_n337), .ZN(new_n342));
  AND4_X1   g0142(.A1(new_n330), .A2(new_n339), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT72), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT17), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n330), .A2(new_n341), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n338), .A2(G169), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n331), .B(G179), .C1(new_n332), .C2(new_n337), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT18), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n330), .A2(new_n341), .B1(new_n347), .B2(new_n348), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT18), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n330), .A2(new_n339), .A3(new_n341), .A4(new_n342), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n344), .A2(KEYINPUT17), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n344), .A2(KEYINPUT17), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n345), .A2(new_n351), .A3(new_n354), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n246), .A2(new_n305), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT12), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n261), .A2(G50), .B1(G20), .B2(new_n305), .ZN(new_n362));
  INV_X1    g0162(.A(G77), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n362), .B1(new_n265), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(KEYINPUT11), .A3(new_n248), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n249), .A2(G68), .A3(new_n254), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n361), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT11), .B1(new_n364), .B2(new_n248), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n277), .A2(G238), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n270), .A2(new_n271), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n370), .B1(new_n372), .B2(new_n272), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n335), .A2(new_n281), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n279), .B(new_n374), .C1(G232), .C2(new_n281), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G97), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n332), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT13), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(new_n376), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n270), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n273), .B1(G238), .B2(new_n277), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT13), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n369), .B1(new_n384), .B2(new_n287), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n293), .B1(new_n378), .B2(new_n383), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(G169), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT14), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT14), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n384), .A2(new_n390), .A3(G169), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n389), .B(new_n391), .C1(new_n300), .C2(new_n384), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n367), .A2(new_n368), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n387), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n250), .A2(new_n255), .A3(new_n363), .ZN(new_n395));
  INV_X1    g0195(.A(new_n266), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(new_n261), .B1(new_n214), .B2(G20), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT15), .B(G87), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n398), .B(KEYINPUT69), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n397), .B1(new_n399), .B2(new_n265), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n400), .A2(new_n248), .ZN(new_n401));
  AOI211_X1 g0201(.A(new_n395), .B(new_n401), .C1(new_n213), .C2(new_n246), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n273), .B1(new_n215), .B2(new_n277), .ZN(new_n403));
  NOR2_X1   g0203(.A1(G232), .A2(G1698), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n281), .A2(G238), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n279), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n406), .B(new_n270), .C1(G107), .C2(new_n279), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(G169), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n408), .A2(new_n300), .ZN(new_n410));
  NOR3_X1   g0210(.A1(new_n402), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n408), .A2(G190), .ZN(new_n413));
  XOR2_X1   g0213(.A(new_n413), .B(KEYINPUT68), .Z(new_n414));
  OAI211_X1 g0214(.A(new_n414), .B(new_n402), .C1(new_n293), .C2(new_n408), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n394), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n303), .A2(new_n359), .A3(new_n416), .ZN(new_n417));
  OR2_X1    g0217(.A1(G250), .A2(G1698), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G257), .B2(new_n281), .ZN(new_n419));
  INV_X1    g0219(.A(G294), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n313), .A2(new_n419), .B1(new_n263), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n270), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT5), .B(G41), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n275), .A2(G1), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n371), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n270), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G264), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n422), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n293), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n422), .A2(new_n287), .A3(new_n428), .A4(new_n426), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT81), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT23), .ZN(new_n435));
  INV_X1    g0235(.A(G107), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n433), .A2(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(G20), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n438), .A2(KEYINPUT81), .B1(new_n439), .B2(G20), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT82), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G116), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n435), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n433), .A2(new_n434), .B1(new_n443), .B2(new_n207), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT82), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n438), .A2(KEYINPUT81), .B1(KEYINPUT23), .B2(G107), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT24), .ZN(new_n449));
  AOI21_X1  g0249(.A(G20), .B1(new_n318), .B2(new_n320), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT22), .ZN(new_n451));
  INV_X1    g0251(.A(G87), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n279), .A2(new_n207), .A3(G87), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n450), .A2(new_n453), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n448), .A2(new_n449), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n449), .B1(new_n448), .B2(new_n455), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n248), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n249), .B1(G1), .B2(new_n263), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT25), .B1(new_n246), .B2(new_n436), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n246), .A2(KEYINPUT25), .A3(new_n436), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n460), .A2(G107), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n432), .A2(new_n458), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT84), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT84), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n432), .A2(new_n458), .A3(new_n467), .A4(new_n464), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n458), .A2(new_n464), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n429), .A2(KEYINPUT83), .A3(G169), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n300), .B2(new_n429), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT83), .B1(new_n429), .B2(G169), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  INV_X1    g0276(.A(G97), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n476), .B(new_n207), .C1(G33), .C2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n478), .B(new_n248), .C1(new_n207), .C2(G116), .ZN(new_n479));
  XOR2_X1   g0279(.A(new_n479), .B(KEYINPUT20), .Z(new_n480));
  INV_X1    g0280(.A(G116), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n246), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n480), .B(new_n482), .C1(new_n481), .C2(new_n459), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT21), .ZN(new_n484));
  OR2_X1    g0284(.A1(G257), .A2(G1698), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(G264), .B2(new_n281), .ZN(new_n486));
  INV_X1    g0286(.A(G303), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n313), .A2(new_n486), .B1(new_n487), .B2(new_n279), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT79), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT79), .ZN(new_n490));
  OAI221_X1 g0290(.A(new_n490), .B1(new_n487), .B2(new_n279), .C1(new_n313), .C2(new_n486), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n270), .A3(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n427), .A2(G270), .B1(new_n371), .B2(new_n425), .ZN(new_n493));
  AOI211_X1 g0293(.A(new_n484), .B(new_n297), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n492), .A2(G179), .A3(new_n493), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n483), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT80), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(KEYINPUT80), .B(new_n483), .C1(new_n494), .C2(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n492), .A2(new_n493), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n483), .A2(new_n500), .A3(G169), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n484), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n483), .B1(new_n500), .B2(G200), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n287), .B2(new_n500), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n498), .A2(new_n499), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n417), .A2(new_n475), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT6), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n508), .A2(new_n477), .A3(G107), .ZN(new_n509));
  XNOR2_X1  g0309(.A(G97), .B(G107), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n509), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  OAI22_X1  g0311(.A1(new_n511), .A2(new_n207), .B1(new_n363), .B2(new_n262), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n436), .B1(new_n325), .B2(new_n327), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n248), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n246), .A2(new_n477), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n460), .A2(G97), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n515), .B1(new_n459), .B2(new_n477), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n262), .A2(new_n363), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n510), .A2(new_n508), .ZN(new_n521));
  INV_X1    g0321(.A(new_n509), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n520), .B1(new_n523), .B2(G20), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n279), .A2(new_n311), .A3(G20), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT7), .B1(new_n326), .B2(new_n207), .ZN(new_n526));
  OAI21_X1  g0326(.A(G107), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n519), .B1(new_n528), .B2(new_n248), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT73), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n423), .A2(new_n424), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(new_n332), .A3(G257), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n426), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G250), .A2(G1698), .ZN(new_n535));
  NAND2_X1  g0335(.A1(KEYINPUT4), .A2(G244), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n535), .B1(new_n536), .B2(G1698), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n476), .B1(new_n538), .B2(new_n326), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G244), .ZN(new_n541));
  AOI211_X1 g0341(.A(new_n541), .B(G1698), .C1(new_n318), .C2(new_n320), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n540), .B1(new_n542), .B2(KEYINPUT4), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n534), .B1(new_n543), .B2(new_n270), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G190), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n426), .A2(new_n533), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n333), .A2(G244), .A3(new_n281), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT4), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n539), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n546), .B1(new_n549), .B2(new_n332), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G200), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n518), .A2(new_n531), .A3(new_n545), .A4(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT74), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(G169), .ZN(new_n554));
  OAI211_X1 g0354(.A(G179), .B(new_n546), .C1(new_n549), .C2(new_n332), .ZN(new_n555));
  AOI211_X1 g0355(.A(new_n553), .B(new_n529), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n555), .B1(new_n544), .B2(new_n297), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT74), .B1(new_n557), .B2(new_n517), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n552), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT75), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT75), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n561), .B(new_n552), .C1(new_n556), .C2(new_n558), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT78), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n332), .A2(G250), .ZN(new_n565));
  XOR2_X1   g0365(.A(new_n424), .B(KEYINPUT76), .Z(new_n566));
  AOI22_X1  g0366(.A1(new_n565), .A2(new_n566), .B1(new_n371), .B2(new_n424), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n333), .A2(G244), .A3(G1698), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n333), .A2(G238), .A3(new_n281), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n442), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT77), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n332), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT77), .A4(new_n442), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n568), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G190), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n313), .A2(new_n541), .A3(new_n281), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n281), .A2(G238), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n442), .B1(new_n313), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n572), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(new_n574), .A3(new_n270), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n567), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G200), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n399), .A2(new_n246), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT19), .B1(new_n264), .B2(G97), .ZN(new_n585));
  NAND3_X1  g0385(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n586));
  NOR2_X1   g0386(.A1(G97), .A2(G107), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n207), .A2(new_n586), .B1(new_n587), .B2(new_n452), .ZN(new_n588));
  AOI211_X1 g0388(.A(new_n585), .B(new_n588), .C1(new_n450), .C2(G68), .ZN(new_n589));
  INV_X1    g0389(.A(new_n248), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n584), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n459), .A2(new_n452), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n576), .A2(new_n583), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n581), .A2(new_n300), .A3(new_n567), .ZN(new_n595));
  OAI221_X1 g0395(.A(new_n584), .B1(new_n459), .B2(new_n399), .C1(new_n589), .C2(new_n590), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n595), .B(new_n596), .C1(new_n575), .C2(G169), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n563), .A2(new_n564), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n557), .A2(new_n517), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n553), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n557), .A2(KEYINPUT74), .A3(new_n517), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n561), .B1(new_n604), .B2(new_n552), .ZN(new_n605));
  INV_X1    g0405(.A(new_n562), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n599), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT78), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n507), .B1(new_n600), .B2(new_n608), .ZN(G372));
  INV_X1    g0409(.A(new_n552), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n602), .B2(new_n603), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT85), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n583), .A2(new_n612), .A3(new_n593), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n293), .B1(new_n581), .B2(new_n567), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n591), .A2(new_n592), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT85), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n613), .A2(new_n616), .A3(new_n576), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n611), .A2(new_n597), .A3(new_n469), .A4(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n474), .A2(new_n496), .A3(new_n502), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n597), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n594), .A2(new_n602), .A3(new_n597), .A4(new_n603), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT26), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n518), .A2(new_n531), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n557), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT86), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT86), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n627), .A3(new_n557), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n617), .A2(new_n597), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n623), .B1(new_n622), .B2(new_n629), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n620), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n417), .ZN(new_n632));
  INV_X1    g0432(.A(new_n302), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n295), .A2(new_n296), .ZN(new_n634));
  INV_X1    g0434(.A(new_n387), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n411), .A2(new_n635), .B1(new_n392), .B2(new_n393), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n345), .A2(new_n358), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n351), .B(new_n354), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n633), .B1(new_n634), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n632), .A2(new_n639), .ZN(G369));
  NAND3_X1  g0440(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G213), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT87), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n645), .A2(G343), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(G343), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n474), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n498), .A2(new_n499), .A3(new_n502), .ZN(new_n650));
  INV_X1    g0450(.A(new_n648), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n469), .A2(new_n474), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT88), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n475), .A2(new_n650), .A3(new_n651), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT88), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(new_n649), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n496), .A2(new_n502), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n483), .A2(new_n648), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n505), .B2(new_n661), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G330), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n470), .A2(new_n648), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n475), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n474), .A2(new_n651), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n659), .A2(new_n670), .ZN(G399));
  INV_X1    g0471(.A(new_n210), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n587), .A2(new_n452), .A3(new_n481), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT89), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n673), .A2(new_n206), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n227), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(new_n673), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT28), .Z(new_n679));
  INV_X1    g0479(.A(new_n597), .ZN(new_n680));
  INV_X1    g0480(.A(new_n621), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n622), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n629), .A2(KEYINPUT26), .ZN(new_n683));
  AND4_X1   g0483(.A1(new_n474), .A2(new_n498), .A3(new_n499), .A4(new_n502), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n682), .B(new_n683), .C1(new_n618), .C2(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n685), .A2(KEYINPUT29), .A3(new_n651), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n631), .A2(new_n651), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT29), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G330), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n505), .A2(new_n653), .A3(new_n648), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n564), .B1(new_n563), .B2(new_n599), .ZN(new_n692));
  AOI211_X1 g0492(.A(KEYINPUT78), .B(new_n598), .C1(new_n560), .C2(new_n562), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n429), .A2(new_n300), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n582), .A2(new_n695), .A3(new_n550), .A4(new_n500), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n495), .A2(new_n544), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT90), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n422), .A2(new_n428), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n575), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n581), .A2(new_n567), .A3(new_n699), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT90), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n697), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n696), .B1(new_n703), .B2(KEYINPUT30), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  AOI211_X1 g0505(.A(new_n705), .B(new_n697), .C1(new_n700), .C2(new_n702), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n648), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT31), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OAI211_X1 g0509(.A(KEYINPUT31), .B(new_n648), .C1(new_n704), .C2(new_n706), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n690), .B1(new_n694), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n689), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n679), .B1(new_n713), .B2(G1), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT91), .ZN(G364));
  NOR2_X1   g0515(.A1(new_n245), .A2(G20), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n206), .B1(new_n716), .B2(G45), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n673), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n665), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(G330), .B2(new_n663), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n672), .A2(new_n326), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G355), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(G116), .B2(new_n210), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n672), .A2(new_n333), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n275), .B2(new_n677), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n240), .A2(new_n275), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G13), .A2(G33), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n223), .B1(G20), .B2(new_n297), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n719), .B1(new_n729), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n207), .A2(G179), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G190), .A2(G200), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n739), .A2(KEYINPUT93), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(KEYINPUT93), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G159), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT32), .Z(new_n745));
  NAND2_X1  g0545(.A1(G20), .A2(G179), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT92), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G200), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n287), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G50), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n737), .A2(G190), .A3(G200), .ZN(new_n751));
  OAI211_X1 g0551(.A(KEYINPUT94), .B(new_n279), .C1(new_n751), .C2(new_n452), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n751), .A2(new_n452), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n326), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n748), .A2(G190), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n753), .B1(KEYINPUT94), .B2(new_n755), .C1(new_n305), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n287), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n747), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n304), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n207), .B1(new_n759), .B2(new_n300), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n737), .A2(new_n287), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n763), .A2(G97), .B1(new_n765), .B2(G107), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n747), .A2(new_n738), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n213), .B2(new_n767), .ZN(new_n768));
  NOR4_X1   g0568(.A1(new_n745), .A2(new_n758), .A3(new_n761), .A4(new_n768), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n769), .A2(KEYINPUT95), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(KEYINPUT95), .ZN(new_n771));
  INV_X1    g0571(.A(G329), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n742), .A2(new_n772), .B1(new_n773), .B2(new_n767), .ZN(new_n774));
  INV_X1    g0574(.A(new_n760), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n774), .B1(G322), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G283), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n326), .B1(new_n764), .B2(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n762), .A2(new_n420), .B1(new_n751), .B2(new_n487), .ZN(new_n779));
  XNOR2_X1  g0579(.A(KEYINPUT33), .B(G317), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n778), .B(new_n779), .C1(new_n756), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G326), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n749), .B(KEYINPUT96), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n776), .B(new_n781), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n770), .A2(new_n771), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n736), .B1(new_n785), .B2(new_n733), .ZN(new_n786));
  INV_X1    g0586(.A(new_n732), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n663), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n721), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(G396));
  INV_X1    g0590(.A(new_n719), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n733), .A2(new_n730), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n791), .B1(new_n363), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n733), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n481), .A2(new_n767), .B1(new_n760), .B2(new_n420), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n764), .A2(new_n452), .B1(new_n751), .B2(new_n436), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n279), .B(new_n796), .C1(G97), .C2(new_n763), .ZN(new_n797));
  INV_X1    g0597(.A(new_n749), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n797), .B1(new_n777), .B2(new_n757), .C1(new_n487), .C2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n742), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n795), .B(new_n799), .C1(G311), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n767), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G143), .A2(new_n775), .B1(new_n802), .B2(G159), .ZN(new_n803));
  INV_X1    g0603(.A(G137), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n757), .B2(new_n260), .C1(new_n804), .C2(new_n798), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT34), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n764), .A2(new_n305), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(G58), .B2(new_n763), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n808), .B(new_n333), .C1(new_n202), .C2(new_n751), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(G132), .B2(new_n800), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n801), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n411), .A2(new_n651), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n402), .A2(new_n651), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n415), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n813), .B1(new_n815), .B2(new_n412), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n793), .B1(new_n794), .B2(new_n811), .C1(new_n816), .C2(new_n731), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n412), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n812), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n687), .A2(new_n819), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n651), .B(new_n816), .C1(new_n620), .C2(new_n630), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n712), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n719), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n822), .A2(new_n823), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n817), .B1(new_n825), .B2(new_n826), .ZN(G384));
  AOI211_X1 g0627(.A(new_n481), .B(new_n225), .C1(new_n523), .C2(KEYINPUT35), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(KEYINPUT35), .B2(new_n523), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT36), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n227), .A2(new_n306), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n831), .A2(new_n213), .B1(G50), .B2(new_n305), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n832), .A2(G1), .A3(new_n245), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT97), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT104), .ZN(new_n836));
  XNOR2_X1  g0636(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT101), .ZN(new_n838));
  INV_X1    g0638(.A(new_n644), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(new_n346), .B2(new_n839), .ZN(new_n840));
  AOI211_X1 g0640(.A(KEYINPUT101), .B(new_n644), .C1(new_n330), .C2(new_n341), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n350), .A2(new_n355), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT37), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n343), .A2(new_n352), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n845), .B(new_n846), .C1(new_n841), .C2(new_n840), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n359), .A2(new_n842), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n837), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n323), .A2(new_n248), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT7), .B1(new_n333), .B2(G20), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(G68), .A3(new_n321), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT16), .B1(new_n853), .B2(new_n310), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n341), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n349), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n839), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(new_n857), .A3(new_n355), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT37), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n847), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n857), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n359), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n862), .A3(KEYINPUT38), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n836), .B1(new_n850), .B2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n844), .A2(new_n847), .B1(new_n359), .B2(new_n842), .ZN(new_n865));
  INV_X1    g0665(.A(new_n837), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n863), .B(new_n836), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n393), .B(new_n648), .C1(new_n392), .C2(new_n387), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT100), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n393), .A2(new_n648), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT99), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n872), .B(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n871), .B1(new_n394), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n391), .B1(new_n300), .B2(new_n384), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n390), .B1(new_n384), .B2(G169), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n393), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND4_X1   g0678(.A1(new_n871), .A2(new_n878), .A3(new_n874), .A4(new_n635), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n870), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n816), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n694), .B2(new_n711), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n869), .A2(new_n882), .A3(KEYINPUT40), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n860), .A2(new_n862), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n863), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n878), .A2(new_n874), .A3(new_n635), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT100), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n819), .B1(new_n889), .B2(new_n870), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n506), .A2(new_n475), .A3(new_n651), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n608), .B2(new_n600), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n709), .A2(new_n710), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n887), .B(new_n890), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n883), .A2(new_n896), .A3(G330), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n712), .A2(new_n417), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n899), .B(KEYINPUT105), .Z(new_n900));
  NAND2_X1  g0700(.A1(new_n694), .A2(new_n711), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n883), .A2(new_n896), .A3(new_n417), .A4(new_n901), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n392), .A2(new_n393), .A3(new_n651), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  INV_X1    g0706(.A(new_n887), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n850), .A2(KEYINPUT103), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n850), .A2(new_n863), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n905), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n880), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n812), .B(KEYINPUT98), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n914), .B1(new_n821), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n887), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n351), .A2(new_n354), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n644), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n913), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n689), .A2(new_n417), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n639), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n920), .B(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n903), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n903), .A2(new_n923), .B1(new_n206), .B2(new_n716), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n835), .B1(new_n925), .B2(new_n926), .ZN(G367));
  OAI221_X1 g0727(.A(new_n734), .B1(new_n210), .B2(new_n399), .C1(new_n726), .C2(new_n236), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n928), .A2(new_n719), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n742), .A2(new_n804), .B1(new_n202), .B2(new_n767), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(G150), .B2(new_n775), .ZN(new_n931));
  INV_X1    g0731(.A(new_n751), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n932), .A2(G58), .B1(new_n765), .B2(new_n214), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n763), .A2(G68), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n933), .A2(new_n279), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(G159), .B2(new_n756), .ZN(new_n936));
  INV_X1    g0736(.A(G143), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n931), .B(new_n936), .C1(new_n937), .C2(new_n783), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n783), .A2(new_n773), .ZN(new_n939));
  XOR2_X1   g0739(.A(KEYINPUT109), .B(G317), .Z(new_n940));
  OAI22_X1  g0740(.A1(new_n742), .A2(new_n940), .B1(new_n487), .B2(new_n760), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(G283), .B2(new_n802), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n313), .B1(new_n477), .B2(new_n764), .C1(new_n436), .C2(new_n762), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n756), .B2(G294), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT108), .B1(new_n751), .B2(new_n481), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT46), .Z(new_n946));
  NAND3_X1  g0746(.A1(new_n942), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n938), .B1(new_n939), .B2(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT47), .Z(new_n949));
  NAND2_X1  g0749(.A1(new_n615), .A2(new_n648), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n617), .A2(new_n597), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n597), .B2(new_n950), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n929), .B1(new_n949), .B2(new_n794), .C1(new_n952), .C2(new_n787), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n673), .B(KEYINPUT41), .Z(new_n954));
  INV_X1    g0754(.A(new_n670), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n624), .A2(new_n648), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n611), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n624), .A2(new_n557), .A3(new_n648), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n655), .A2(new_n658), .A3(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT44), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n654), .A2(KEYINPUT88), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n657), .B1(new_n656), .B2(new_n649), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n659), .A2(new_n959), .A3(new_n966), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n955), .B1(new_n962), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT44), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n961), .B(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n973), .A2(new_n670), .A3(new_n969), .A4(new_n968), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n667), .A2(new_n668), .A3(new_n652), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n656), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(new_n664), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n689), .A2(new_n977), .A3(new_n712), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n971), .A2(new_n974), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n954), .B1(new_n979), .B2(new_n713), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n980), .A2(new_n718), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT42), .ZN(new_n982));
  OR3_X1    g0782(.A1(new_n960), .A2(new_n656), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n982), .B1(new_n960), .B2(new_n656), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n604), .B1(new_n960), .B2(new_n474), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n983), .A2(new_n984), .B1(new_n651), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT106), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n952), .B(KEYINPUT43), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n987), .B1(new_n986), .B2(new_n988), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n670), .A2(new_n960), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n993), .B(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n953), .B1(new_n981), .B2(new_n996), .ZN(G387));
  INV_X1    g0797(.A(new_n978), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n977), .B1(new_n689), .B2(new_n712), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n998), .A2(new_n673), .A3(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n722), .A2(new_n675), .B1(new_n436), .B2(new_n672), .ZN(new_n1001));
  AOI211_X1 g0801(.A(G45), .B(new_n675), .C1(G68), .C2(G77), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT110), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n396), .A2(new_n202), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT50), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n725), .B1(new_n233), .B2(new_n275), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1001), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n791), .B1(new_n1010), .B2(new_n734), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n333), .B1(new_n477), .B2(new_n764), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n214), .B2(new_n932), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n757), .B2(new_n266), .C1(new_n743), .C2(new_n798), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n399), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n763), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n305), .B2(new_n767), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n742), .A2(new_n260), .B1(new_n202), .B2(new_n760), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1014), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n802), .A2(G303), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n760), .B2(new_n940), .C1(new_n757), .C2(new_n773), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n783), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1021), .B1(new_n1022), .B2(G322), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1023), .A2(KEYINPUT48), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(KEYINPUT48), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n763), .A2(G283), .B1(new_n932), .B2(G294), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT49), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n313), .B1(new_n481), .B2(new_n764), .C1(new_n742), .C2(new_n782), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT111), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1019), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1011), .B1(new_n669), .B2(new_n787), .C1(new_n1034), .C2(new_n794), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1000), .B(new_n1035), .C1(new_n717), .C2(new_n977), .ZN(G393));
  NAND2_X1  g0836(.A1(new_n971), .A2(new_n974), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n998), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1038), .A2(new_n673), .A3(new_n979), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n971), .A2(new_n974), .A3(new_n718), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n734), .B1(new_n477), .B2(new_n210), .C1(new_n726), .C2(new_n243), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n719), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n762), .A2(new_n363), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n333), .B1(new_n452), .B2(new_n764), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1043), .B(new_n1044), .C1(G68), .C2(new_n932), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n800), .A2(G143), .B1(new_n396), .B2(new_n802), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(new_n202), .C2(new_n757), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n749), .A2(G150), .B1(new_n775), .B2(G159), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT51), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n749), .A2(G317), .B1(new_n775), .B2(G311), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT52), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n800), .A2(G322), .B1(G294), .B2(new_n802), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n762), .A2(new_n481), .B1(new_n751), .B2(new_n777), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n279), .B(new_n1053), .C1(G107), .C2(new_n765), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1052), .B(new_n1054), .C1(new_n487), .C2(new_n757), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1047), .A2(new_n1049), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1042), .B1(new_n1056), .B2(new_n733), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n959), .B2(new_n787), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1040), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1039), .A2(new_n1059), .ZN(G390));
  INV_X1    g0860(.A(new_n792), .ZN(new_n1061));
  INV_X1    g0861(.A(G132), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n760), .A2(new_n1062), .B1(new_n743), .B2(new_n762), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n751), .A2(new_n260), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1064), .B(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(G128), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1066), .B1(new_n757), .B2(new_n804), .C1(new_n1067), .C2(new_n798), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT54), .B(G143), .Z(new_n1069));
  AOI211_X1 g0869(.A(new_n1063), .B(new_n1068), .C1(new_n802), .C2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n279), .B1(new_n764), .B2(new_n202), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n800), .B2(G125), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT113), .Z(new_n1073));
  OAI22_X1  g0873(.A1(new_n477), .A2(new_n767), .B1(new_n760), .B2(new_n481), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G294), .B2(new_n800), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n757), .A2(new_n436), .ZN(new_n1076));
  OR4_X1    g0876(.A1(new_n279), .A2(new_n1043), .A3(new_n754), .A4(new_n807), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(G283), .C2(new_n749), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1070), .A2(new_n1073), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n719), .B1(new_n396), .B2(new_n1061), .C1(new_n1079), .C2(new_n794), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n865), .A2(new_n866), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT103), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n886), .B(new_n863), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n863), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1083), .A2(KEYINPUT39), .B1(new_n1085), .B2(new_n910), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1080), .B1(new_n1086), .B2(new_n730), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n821), .A2(new_n915), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n905), .B1(new_n1089), .B2(new_n880), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1083), .A2(KEYINPUT39), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n911), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n685), .A2(new_n651), .A3(new_n816), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n914), .B1(new_n1093), .B2(new_n915), .ZN(new_n1094));
  OAI21_X1  g0894(.A(KEYINPUT104), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(new_n904), .A3(new_n867), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1090), .A2(new_n1092), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(G330), .B(new_n816), .C1(new_n892), .C2(new_n893), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1098), .A2(new_n914), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1093), .A2(new_n915), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n880), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1096), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1086), .B1(new_n916), .B2(new_n905), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n712), .A2(new_n816), .A3(new_n880), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1100), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1088), .B1(new_n1108), .B2(new_n717), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n921), .A2(new_n898), .A3(new_n639), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1098), .A2(new_n914), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(KEYINPUT112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1101), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT112), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1098), .A2(new_n1115), .A3(new_n914), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1113), .A2(new_n1114), .A3(new_n1106), .A4(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1112), .A2(new_n1106), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n1089), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1111), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1106), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n673), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1110), .B1(new_n1125), .B2(new_n1126), .ZN(G378));
  OAI21_X1  g0927(.A(new_n719), .B1(new_n1061), .B2(G50), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n934), .B1(new_n304), .B2(new_n764), .C1(new_n399), .C2(new_n767), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n313), .A2(new_n274), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n214), .B2(new_n932), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT115), .Z(new_n1132));
  OAI22_X1  g0932(.A1(new_n742), .A2(new_n777), .B1(new_n436), .B2(new_n760), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n477), .A2(new_n757), .B1(new_n798), .B2(new_n481), .ZN(new_n1134));
  OR4_X1    g0934(.A1(new_n1129), .A2(new_n1132), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT58), .ZN(new_n1136));
  AOI21_X1  g0936(.A(G50), .B1(new_n263), .B2(new_n274), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1135), .A2(new_n1136), .B1(new_n1130), .B2(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n802), .A2(G137), .B1(new_n932), .B2(new_n1069), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n1067), .B2(new_n760), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(G132), .B2(new_n756), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n749), .A2(G125), .B1(G150), .B2(new_n763), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1142), .A2(KEYINPUT116), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1142), .A2(KEYINPUT116), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1141), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(KEYINPUT59), .ZN(new_n1146));
  AOI211_X1 g0946(.A(G33), .B(G41), .C1(new_n765), .C2(G159), .ZN(new_n1147));
  INV_X1    g0947(.A(G124), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(new_n1148), .B2(new_n742), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT117), .Z(new_n1150));
  NAND2_X1  g0950(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1145), .A2(KEYINPUT59), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1138), .B1(new_n1136), .B2(new_n1135), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1128), .B1(new_n1153), .B2(new_n733), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n299), .A2(new_n839), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n634), .A2(new_n302), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n303), .A2(new_n299), .A3(new_n839), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1158), .B(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1154), .B1(new_n1161), .B2(new_n731), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT118), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1161), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n897), .A2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1161), .A2(new_n883), .A3(new_n896), .A4(G330), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n920), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1165), .A2(new_n920), .A3(new_n1166), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1163), .B1(new_n1171), .B2(new_n718), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1165), .A2(new_n920), .A3(new_n1166), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n920), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1174));
  OAI21_X1  g0974(.A(KEYINPUT57), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1111), .B1(new_n1123), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n673), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1111), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1116), .A2(new_n1114), .A3(new_n1106), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1180), .A2(new_n1113), .B1(new_n1089), .B2(new_n1118), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1179), .B1(new_n1181), .B2(new_n1108), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT57), .B1(new_n1171), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1172), .B1(new_n1178), .B2(new_n1183), .ZN(G375));
  AOI21_X1  g0984(.A(new_n791), .B1(new_n305), .B2(new_n792), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n279), .B1(new_n932), .B2(G97), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1186), .B1(new_n363), .B2(new_n764), .C1(new_n742), .C2(new_n487), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1016), .B1(new_n777), .B2(new_n760), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT120), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1187), .B(new_n1189), .C1(G294), .C2(new_n749), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n756), .A2(G116), .B1(new_n802), .B2(G107), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT119), .Z(new_n1192));
  AOI22_X1  g0992(.A1(new_n756), .A2(new_n1069), .B1(new_n775), .B2(G137), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n1062), .B2(new_n798), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT121), .Z(new_n1195));
  OAI22_X1  g0995(.A1(new_n742), .A2(new_n1067), .B1(new_n260), .B2(new_n767), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n333), .B1(new_n304), .B2(new_n764), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n762), .A2(new_n202), .B1(new_n751), .B2(new_n743), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1190), .A2(new_n1192), .B1(new_n1195), .B2(new_n1199), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1185), .B1(new_n794), .B2(new_n1200), .C1(new_n880), .C2(new_n731), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n1181), .B2(new_n717), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1120), .A2(new_n954), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1203), .B1(new_n1204), .B2(new_n1205), .ZN(G381));
  NOR4_X1   g1006(.A1(G390), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n993), .B(new_n994), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n718), .B2(new_n980), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1209), .A3(new_n953), .ZN(new_n1210));
  OR4_X1    g1010(.A1(G378), .A2(new_n1210), .A3(G375), .A4(G381), .ZN(G407));
  NAND3_X1  g1011(.A1(new_n646), .A2(new_n647), .A3(G213), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(G375), .A2(G378), .A3(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT122), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(G213), .A3(G407), .ZN(G409));
  OAI211_X1 g1015(.A(G378), .B(new_n1172), .C1(new_n1178), .C2(new_n1183), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n673), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1217), .B1(new_n1218), .B2(new_n1108), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1109), .B1(new_n1219), .B2(new_n1124), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1221), .A2(new_n1177), .A3(new_n954), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1163), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1221), .B2(new_n717), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1220), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1216), .A2(new_n1225), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1117), .A2(new_n1111), .A3(KEYINPUT60), .A4(new_n1119), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n673), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1218), .A2(KEYINPUT60), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1181), .A2(new_n1111), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1228), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(G384), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n1202), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1227), .A2(new_n673), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT60), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1120), .A2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1234), .B1(new_n1236), .B2(new_n1205), .ZN(new_n1237));
  AOI21_X1  g1037(.A(G384), .B1(new_n1237), .B2(new_n1203), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1233), .A2(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1226), .A2(new_n1239), .A3(KEYINPUT63), .A4(new_n1212), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1209), .A2(new_n953), .A3(G390), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT125), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT124), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G390), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1039), .A2(KEYINPUT124), .A3(new_n1059), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(G387), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(G393), .B(new_n789), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT125), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1209), .A2(new_n1249), .A3(G390), .A4(new_n953), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1242), .A2(new_n1246), .A3(new_n1248), .A4(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1241), .ZN(new_n1252));
  AOI21_X1  g1052(.A(G390), .B1(new_n1209), .B2(new_n953), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1247), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1251), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT61), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1240), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1226), .A2(KEYINPUT123), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT123), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1216), .A2(new_n1225), .A3(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1212), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1212), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(G2897), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1233), .A2(new_n1238), .A3(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1232), .B1(new_n1231), .B2(new_n1202), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1237), .A2(G384), .A3(new_n1203), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1265), .A2(new_n1266), .B1(G2897), .B2(new_n1262), .ZN(new_n1267));
  OR2_X1    g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1261), .A2(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1258), .A2(new_n1212), .A3(new_n1239), .A4(new_n1260), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1257), .B(new_n1269), .C1(new_n1271), .C2(KEYINPUT63), .ZN(new_n1272));
  XOR2_X1   g1072(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1273));
  NOR2_X1   g1073(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1262), .B1(new_n1216), .B2(new_n1225), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  XOR2_X1   g1076(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1277));
  NAND2_X1  g1077(.A1(new_n1270), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1275), .A2(KEYINPUT62), .A3(new_n1239), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1276), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1272), .B1(new_n1280), .B2(new_n1255), .ZN(G405));
  NAND2_X1  g1081(.A1(G375), .A2(new_n1220), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1255), .A2(new_n1216), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1216), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1284), .A2(new_n1254), .A3(new_n1251), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1286), .B(new_n1239), .ZN(G402));
endmodule


