

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U321 ( .A(n304), .B(n303), .ZN(n306) );
  XNOR2_X1 U322 ( .A(n302), .B(n301), .ZN(n303) );
  OR2_X1 U323 ( .A1(n549), .A2(n567), .ZN(n366) );
  NOR2_X1 U324 ( .A1(n542), .A2(n368), .ZN(n369) );
  XNOR2_X1 U325 ( .A(n359), .B(KEYINPUT45), .ZN(n360) );
  XNOR2_X1 U326 ( .A(G120GAT), .B(G148GAT), .ZN(n309) );
  XNOR2_X1 U327 ( .A(n361), .B(n360), .ZN(n362) );
  INV_X1 U328 ( .A(KEYINPUT90), .ZN(n379) );
  XNOR2_X1 U329 ( .A(n309), .B(G57GAT), .ZN(n394) );
  XNOR2_X1 U330 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U331 ( .A(n313), .B(n312), .ZN(n314) );
  INV_X1 U332 ( .A(KEYINPUT97), .ZN(n469) );
  XNOR2_X1 U333 ( .A(n315), .B(n314), .ZN(n319) );
  XNOR2_X1 U334 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n430) );
  XNOR2_X1 U335 ( .A(n333), .B(KEYINPUT71), .ZN(n334) );
  XNOR2_X1 U336 ( .A(n431), .B(n430), .ZN(n446) );
  XNOR2_X1 U337 ( .A(n335), .B(n334), .ZN(n337) );
  NOR2_X1 U338 ( .A1(n446), .A2(n531), .ZN(n562) );
  XOR2_X1 U339 ( .A(n308), .B(n307), .Z(n555) );
  INV_X1 U340 ( .A(G43GAT), .ZN(n475) );
  XOR2_X1 U341 ( .A(n392), .B(n391), .Z(n518) );
  XNOR2_X1 U342 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n447) );
  XNOR2_X1 U343 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U344 ( .A(n448), .B(n447), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(n478), .B(n477), .ZN(G1330GAT) );
  XOR2_X1 U346 ( .A(G92GAT), .B(KEYINPUT11), .Z(n290) );
  XNOR2_X1 U347 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n289) );
  XNOR2_X1 U348 ( .A(n290), .B(n289), .ZN(n308) );
  XNOR2_X1 U349 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n291) );
  XNOR2_X1 U350 ( .A(n291), .B(G29GAT), .ZN(n292) );
  XOR2_X1 U351 ( .A(n292), .B(KEYINPUT8), .Z(n294) );
  XNOR2_X1 U352 ( .A(G43GAT), .B(G50GAT), .ZN(n293) );
  XOR2_X1 U353 ( .A(n294), .B(n293), .Z(n336) );
  INV_X1 U354 ( .A(G134GAT), .ZN(n295) );
  XNOR2_X1 U355 ( .A(n336), .B(n295), .ZN(n304) );
  XNOR2_X1 U356 ( .A(G99GAT), .B(G85GAT), .ZN(n296) );
  XNOR2_X1 U357 ( .A(n296), .B(KEYINPUT76), .ZN(n317) );
  XOR2_X1 U358 ( .A(n317), .B(G162GAT), .Z(n302) );
  XOR2_X1 U359 ( .A(KEYINPUT68), .B(KEYINPUT66), .Z(n298) );
  XNOR2_X1 U360 ( .A(G190GAT), .B(KEYINPUT9), .ZN(n297) );
  XNOR2_X1 U361 ( .A(n298), .B(n297), .ZN(n300) );
  XOR2_X1 U362 ( .A(G218GAT), .B(KEYINPUT67), .Z(n299) );
  XNOR2_X1 U363 ( .A(n300), .B(n299), .ZN(n301) );
  NAND2_X1 U364 ( .A1(G232GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U365 ( .A(n306), .B(n305), .ZN(n307) );
  INV_X1 U366 ( .A(n555), .ZN(n542) );
  XOR2_X1 U367 ( .A(G71GAT), .B(KEYINPUT13), .Z(n345) );
  XOR2_X1 U368 ( .A(n394), .B(n345), .Z(n315) );
  XOR2_X1 U369 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n311) );
  XNOR2_X1 U370 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n313) );
  NAND2_X1 U372 ( .A1(G230GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U373 ( .A(G106GAT), .B(G78GAT), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n316), .B(KEYINPUT75), .ZN(n422) );
  XOR2_X1 U375 ( .A(n422), .B(n317), .Z(n318) );
  XNOR2_X1 U376 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U377 ( .A(G64GAT), .B(KEYINPUT77), .Z(n321) );
  XNOR2_X1 U378 ( .A(G204GAT), .B(G92GAT), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U380 ( .A(G176GAT), .B(n322), .Z(n384) );
  XNOR2_X1 U381 ( .A(n323), .B(n384), .ZN(n364) );
  INV_X1 U382 ( .A(n364), .ZN(n572) );
  XOR2_X1 U383 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n325) );
  XNOR2_X1 U384 ( .A(KEYINPUT70), .B(KEYINPUT73), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U386 ( .A(G169GAT), .B(G8GAT), .Z(n382) );
  XOR2_X1 U387 ( .A(G22GAT), .B(G15GAT), .Z(n346) );
  XNOR2_X1 U388 ( .A(n382), .B(n346), .ZN(n327) );
  XOR2_X1 U389 ( .A(KEYINPUT69), .B(G197GAT), .Z(n326) );
  XNOR2_X1 U390 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U391 ( .A(n329), .B(n328), .Z(n331) );
  NAND2_X1 U392 ( .A1(G229GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n331), .B(n330), .ZN(n335) );
  XNOR2_X1 U394 ( .A(G141GAT), .B(G113GAT), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n332), .B(G1GAT), .ZN(n408) );
  XNOR2_X1 U396 ( .A(n408), .B(KEYINPUT72), .ZN(n333) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n567) );
  XOR2_X1 U398 ( .A(KEYINPUT74), .B(n567), .Z(n532) );
  INV_X1 U399 ( .A(n532), .ZN(n338) );
  NAND2_X1 U400 ( .A1(n572), .A2(n338), .ZN(n363) );
  XOR2_X1 U401 ( .A(G78GAT), .B(G155GAT), .Z(n340) );
  XNOR2_X1 U402 ( .A(G183GAT), .B(G211GAT), .ZN(n339) );
  XNOR2_X1 U403 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U404 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n342) );
  XNOR2_X1 U405 ( .A(G8GAT), .B(KEYINPUT12), .ZN(n341) );
  XNOR2_X1 U406 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U407 ( .A(n344), .B(n343), .Z(n348) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U410 ( .A(KEYINPUT79), .B(KEYINPUT81), .Z(n350) );
  NAND2_X1 U411 ( .A1(G231GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U413 ( .A(n352), .B(n351), .Z(n357) );
  XOR2_X1 U414 ( .A(G64GAT), .B(G57GAT), .Z(n354) );
  XNOR2_X1 U415 ( .A(G1GAT), .B(G127GAT), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n355), .B(KEYINPUT80), .ZN(n356) );
  XOR2_X1 U418 ( .A(n357), .B(n356), .Z(n563) );
  INV_X1 U419 ( .A(n563), .ZN(n577) );
  XOR2_X1 U420 ( .A(KEYINPUT36), .B(KEYINPUT101), .Z(n358) );
  XNOR2_X1 U421 ( .A(n555), .B(n358), .ZN(n580) );
  NOR2_X1 U422 ( .A1(n577), .A2(n580), .ZN(n361) );
  INV_X1 U423 ( .A(KEYINPUT114), .ZN(n359) );
  OR2_X1 U424 ( .A1(n363), .A2(n362), .ZN(n373) );
  XOR2_X1 U425 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n367) );
  XNOR2_X1 U426 ( .A(n364), .B(KEYINPUT64), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n365), .B(KEYINPUT41), .ZN(n549) );
  XNOR2_X1 U428 ( .A(n367), .B(n366), .ZN(n368) );
  NAND2_X1 U429 ( .A1(n577), .A2(n369), .ZN(n370) );
  XNOR2_X1 U430 ( .A(KEYINPUT113), .B(n370), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n371), .B(KEYINPUT47), .ZN(n372) );
  NAND2_X1 U432 ( .A1(n373), .A2(n372), .ZN(n375) );
  INV_X1 U433 ( .A(KEYINPUT48), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n527) );
  XOR2_X1 U435 ( .A(KEYINPUT17), .B(G190GAT), .Z(n377) );
  XNOR2_X1 U436 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U438 ( .A(KEYINPUT19), .B(n378), .Z(n445) );
  NAND2_X1 U439 ( .A1(G226GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U441 ( .A(n383), .B(KEYINPUT91), .Z(n386) );
  XNOR2_X1 U442 ( .A(G36GAT), .B(n384), .ZN(n385) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n445), .B(n387), .ZN(n392) );
  XOR2_X1 U445 ( .A(KEYINPUT83), .B(G218GAT), .Z(n389) );
  XNOR2_X1 U446 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U448 ( .A(G197GAT), .B(n390), .ZN(n427) );
  INV_X1 U449 ( .A(n427), .ZN(n391) );
  NOR2_X1 U450 ( .A1(n527), .A2(n518), .ZN(n393) );
  XNOR2_X1 U451 ( .A(KEYINPUT54), .B(n393), .ZN(n411) );
  XOR2_X1 U452 ( .A(G85GAT), .B(n394), .Z(n396) );
  XNOR2_X1 U453 ( .A(G29GAT), .B(KEYINPUT4), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U455 ( .A(n397), .B(KEYINPUT1), .Z(n402) );
  XOR2_X1 U456 ( .A(KEYINPUT88), .B(KEYINPUT5), .Z(n399) );
  NAND2_X1 U457 ( .A1(G225GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U459 ( .A(KEYINPUT6), .B(n400), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U461 ( .A(KEYINPUT84), .B(G162GAT), .Z(n404) );
  XNOR2_X1 U462 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U464 ( .A(KEYINPUT2), .B(n405), .Z(n419) );
  XOR2_X1 U465 ( .A(n406), .B(n419), .Z(n410) );
  XNOR2_X1 U466 ( .A(G134GAT), .B(G127GAT), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n407), .B(KEYINPUT0), .ZN(n432) );
  XNOR2_X1 U468 ( .A(n408), .B(n432), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n410), .B(n409), .ZN(n466) );
  XNOR2_X1 U470 ( .A(KEYINPUT89), .B(n466), .ZN(n515) );
  NAND2_X1 U471 ( .A1(n411), .A2(n515), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n412), .B(KEYINPUT65), .ZN(n565) );
  XOR2_X1 U473 ( .A(G148GAT), .B(G204GAT), .Z(n414) );
  XNOR2_X1 U474 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U476 ( .A(G22GAT), .B(n415), .Z(n417) );
  NAND2_X1 U477 ( .A1(G228GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U479 ( .A(n418), .B(KEYINPUT24), .Z(n421) );
  XNOR2_X1 U480 ( .A(G141GAT), .B(n419), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n426) );
  XOR2_X1 U482 ( .A(KEYINPUT23), .B(n422), .Z(n424) );
  XNOR2_X1 U483 ( .A(G50GAT), .B(KEYINPUT87), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U485 ( .A(n426), .B(n425), .Z(n429) );
  XOR2_X1 U486 ( .A(n427), .B(KEYINPUT22), .Z(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n457) );
  NAND2_X1 U488 ( .A1(n565), .A2(n457), .ZN(n431) );
  XOR2_X1 U489 ( .A(n432), .B(G99GAT), .Z(n434) );
  NAND2_X1 U490 ( .A1(G227GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U492 ( .A(G120GAT), .B(G71GAT), .Z(n436) );
  XNOR2_X1 U493 ( .A(G113GAT), .B(G15GAT), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U495 ( .A(n438), .B(n437), .Z(n443) );
  XOR2_X1 U496 ( .A(G176GAT), .B(KEYINPUT82), .Z(n440) );
  XNOR2_X1 U497 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n439) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U499 ( .A(G43GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U501 ( .A(n445), .B(n444), .Z(n458) );
  INV_X1 U502 ( .A(n458), .ZN(n531) );
  NAND2_X1 U503 ( .A1(n542), .A2(n562), .ZN(n448) );
  XOR2_X1 U504 ( .A(KEYINPUT102), .B(KEYINPUT37), .Z(n473) );
  XNOR2_X1 U505 ( .A(n457), .B(KEYINPUT28), .ZN(n529) );
  INV_X1 U506 ( .A(n529), .ZN(n451) );
  XNOR2_X1 U507 ( .A(KEYINPUT27), .B(KEYINPUT92), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n449), .B(n518), .ZN(n460) );
  NOR2_X1 U509 ( .A1(n460), .A2(n515), .ZN(n450) );
  XNOR2_X1 U510 ( .A(n450), .B(KEYINPUT93), .ZN(n526) );
  NOR2_X1 U511 ( .A1(n451), .A2(n526), .ZN(n452) );
  XOR2_X1 U512 ( .A(KEYINPUT94), .B(n452), .Z(n453) );
  NOR2_X1 U513 ( .A1(n458), .A2(n453), .ZN(n468) );
  NOR2_X1 U514 ( .A1(n531), .A2(n518), .ZN(n454) );
  XOR2_X1 U515 ( .A(KEYINPUT96), .B(n454), .Z(n455) );
  NAND2_X1 U516 ( .A1(n457), .A2(n455), .ZN(n456) );
  XNOR2_X1 U517 ( .A(KEYINPUT25), .B(n456), .ZN(n464) );
  NOR2_X1 U518 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U519 ( .A(KEYINPUT26), .B(n459), .ZN(n566) );
  INV_X1 U520 ( .A(n566), .ZN(n461) );
  NOR2_X1 U521 ( .A1(n461), .A2(n460), .ZN(n462) );
  XOR2_X1 U522 ( .A(KEYINPUT95), .B(n462), .Z(n463) );
  NOR2_X1 U523 ( .A1(n464), .A2(n463), .ZN(n465) );
  NOR2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n468), .A2(n467), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n470), .B(n469), .ZN(n483) );
  NOR2_X1 U527 ( .A1(n483), .A2(n580), .ZN(n471) );
  NAND2_X1 U528 ( .A1(n471), .A2(n577), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n473), .B(n472), .ZN(n514) );
  NAND2_X1 U530 ( .A1(n572), .A2(n532), .ZN(n485) );
  NOR2_X1 U531 ( .A1(n514), .A2(n485), .ZN(n474) );
  XOR2_X1 U532 ( .A(KEYINPUT38), .B(n474), .Z(n499) );
  NOR2_X1 U533 ( .A1(n499), .A2(n531), .ZN(n478) );
  XNOR2_X1 U534 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n476) );
  NAND2_X1 U535 ( .A1(n532), .A2(n562), .ZN(n480) );
  XNOR2_X1 U536 ( .A(KEYINPUT122), .B(G169GAT), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n480), .B(n479), .ZN(G1348GAT) );
  NOR2_X1 U538 ( .A1(n577), .A2(n542), .ZN(n481) );
  XOR2_X1 U539 ( .A(KEYINPUT16), .B(n481), .Z(n482) );
  NOR2_X1 U540 ( .A1(n483), .A2(n482), .ZN(n484) );
  XOR2_X1 U541 ( .A(KEYINPUT98), .B(n484), .Z(n502) );
  OR2_X1 U542 ( .A1(n502), .A2(n485), .ZN(n493) );
  NOR2_X1 U543 ( .A1(n515), .A2(n493), .ZN(n486) );
  XOR2_X1 U544 ( .A(n486), .B(KEYINPUT34), .Z(n487) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  NOR2_X1 U546 ( .A1(n518), .A2(n493), .ZN(n488) );
  XOR2_X1 U547 ( .A(G8GAT), .B(n488), .Z(G1325GAT) );
  NOR2_X1 U548 ( .A1(n493), .A2(n531), .ZN(n492) );
  XOR2_X1 U549 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n490) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1326GAT) );
  NOR2_X1 U553 ( .A1(n529), .A2(n493), .ZN(n494) );
  XOR2_X1 U554 ( .A(G22GAT), .B(n494), .Z(G1327GAT) );
  NOR2_X1 U555 ( .A1(n499), .A2(n515), .ZN(n496) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  NOR2_X1 U558 ( .A1(n499), .A2(n518), .ZN(n498) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1329GAT) );
  NOR2_X1 U561 ( .A1(n499), .A2(n529), .ZN(n500) );
  XOR2_X1 U562 ( .A(G50GAT), .B(n500), .Z(G1331GAT) );
  INV_X1 U563 ( .A(n549), .ZN(n557) );
  NAND2_X1 U564 ( .A1(n567), .A2(n557), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n501), .B(KEYINPUT106), .ZN(n513) );
  OR2_X1 U566 ( .A1(n502), .A2(n513), .ZN(n509) );
  NOR2_X1 U567 ( .A1(n515), .A2(n509), .ZN(n504) );
  XNOR2_X1 U568 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  NOR2_X1 U571 ( .A1(n518), .A2(n509), .ZN(n506) );
  XOR2_X1 U572 ( .A(G64GAT), .B(n506), .Z(G1333GAT) );
  NOR2_X1 U573 ( .A1(n531), .A2(n509), .ZN(n508) );
  XNOR2_X1 U574 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(G1334GAT) );
  NOR2_X1 U576 ( .A1(n529), .A2(n509), .ZN(n511) );
  XNOR2_X1 U577 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(n512), .ZN(G1335GAT) );
  OR2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n522) );
  NOR2_X1 U581 ( .A1(n515), .A2(n522), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(G1336GAT) );
  NOR2_X1 U584 ( .A1(n518), .A2(n522), .ZN(n519) );
  XOR2_X1 U585 ( .A(KEYINPUT110), .B(n519), .Z(n520) );
  XNOR2_X1 U586 ( .A(G92GAT), .B(n520), .ZN(G1337GAT) );
  NOR2_X1 U587 ( .A1(n531), .A2(n522), .ZN(n521) );
  XOR2_X1 U588 ( .A(G99GAT), .B(n521), .Z(G1338GAT) );
  NOR2_X1 U589 ( .A1(n529), .A2(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(KEYINPUT111), .B(KEYINPUT44), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  NOR2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U594 ( .A(n528), .B(KEYINPUT115), .Z(n547) );
  NAND2_X1 U595 ( .A1(n547), .A2(n529), .ZN(n530) );
  NOR2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n543), .A2(n532), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U600 ( .A1(n543), .A2(n557), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(G120GAT), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n538) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(KEYINPUT118), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U606 ( .A(KEYINPUT117), .B(n539), .Z(n541) );
  NAND2_X1 U607 ( .A1(n543), .A2(n563), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(G134GAT), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U613 ( .A1(n547), .A2(n566), .ZN(n554) );
  NOR2_X1 U614 ( .A1(n567), .A2(n554), .ZN(n548) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n548), .Z(G1344GAT) );
  NOR2_X1 U616 ( .A1(n549), .A2(n554), .ZN(n551) );
  XNOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(n552), .ZN(G1345GAT) );
  NOR2_X1 U620 ( .A1(n577), .A2(n554), .ZN(n553) );
  XOR2_X1 U621 ( .A(G155GAT), .B(n553), .Z(G1346GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U623 ( .A(G162GAT), .B(n556), .Z(G1347GAT) );
  NAND2_X1 U624 ( .A1(n562), .A2(n557), .ZN(n559) );
  XOR2_X1 U625 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n561) );
  XOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT56), .Z(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n566), .ZN(n579) );
  NOR2_X1 U632 ( .A1(n567), .A2(n579), .ZN(n571) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(KEYINPUT60), .ZN(n569) );
  XNOR2_X1 U635 ( .A(KEYINPUT124), .B(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  NOR2_X1 U637 ( .A1(n579), .A2(n572), .ZN(n576) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n574) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n579), .ZN(n578) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n578), .Z(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

