

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U556 ( .A(n682), .B(n681), .ZN(n711) );
  AND2_X2 U557 ( .A1(n680), .A2(n679), .ZN(n682) );
  NOR2_X1 U558 ( .A1(n724), .A2(n723), .ZN(n725) );
  OR2_X1 U559 ( .A1(n666), .A2(n665), .ZN(n712) );
  OR2_X2 U560 ( .A1(n702), .A2(n703), .ZN(n672) );
  AND2_X1 U561 ( .A1(n545), .A2(n544), .ZN(n546) );
  OR2_X2 U562 ( .A1(n623), .A2(n973), .ZN(n624) );
  XNOR2_X2 U563 ( .A(n546), .B(KEYINPUT84), .ZN(G164) );
  AND2_X1 U564 ( .A1(n708), .A2(n522), .ZN(n709) );
  XNOR2_X1 U565 ( .A(n525), .B(KEYINPUT17), .ZN(n537) );
  NOR2_X1 U566 ( .A1(n619), .A2(n618), .ZN(n620) );
  INV_X1 U567 ( .A(G2105), .ZN(n524) );
  OR2_X1 U568 ( .A1(n707), .A2(n720), .ZN(n522) );
  INV_X1 U569 ( .A(n672), .ZN(n642) );
  NAND2_X1 U570 ( .A1(G8), .A2(n672), .ZN(n720) );
  NOR2_X1 U571 ( .A1(G1384), .A2(G164), .ZN(n597) );
  XNOR2_X1 U572 ( .A(n597), .B(KEYINPUT65), .ZN(n702) );
  INV_X1 U573 ( .A(G2104), .ZN(n523) );
  INV_X1 U574 ( .A(n702), .ZN(n704) );
  NAND2_X1 U575 ( .A1(n524), .A2(n523), .ZN(n525) );
  AND2_X2 U576 ( .A1(n524), .A2(G2104), .ZN(n891) );
  INV_X1 U577 ( .A(KEYINPUT23), .ZN(n529) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n800) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n895) );
  INV_X1 U580 ( .A(KEYINPUT67), .ZN(n533) );
  NOR2_X1 U581 ( .A1(n536), .A2(n535), .ZN(G160) );
  INV_X1 U582 ( .A(n537), .ZN(n526) );
  INV_X1 U583 ( .A(n526), .ZN(n890) );
  NAND2_X1 U584 ( .A1(G137), .A2(n890), .ZN(n528) );
  NAND2_X1 U585 ( .A1(G113), .A2(n895), .ZN(n527) );
  NAND2_X1 U586 ( .A1(n528), .A2(n527), .ZN(n536) );
  AND2_X1 U587 ( .A1(G2105), .A2(n523), .ZN(n894) );
  NAND2_X1 U588 ( .A1(n894), .A2(G125), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n891), .A2(G101), .ZN(n530) );
  XNOR2_X1 U590 ( .A(n530), .B(n529), .ZN(n531) );
  NAND2_X1 U591 ( .A1(n532), .A2(n531), .ZN(n534) );
  XNOR2_X1 U592 ( .A(n534), .B(n533), .ZN(n535) );
  NAND2_X1 U593 ( .A1(G138), .A2(n537), .ZN(n539) );
  NAND2_X1 U594 ( .A1(G102), .A2(n891), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U596 ( .A(n540), .B(KEYINPUT83), .ZN(n545) );
  AND2_X1 U597 ( .A1(G2105), .A2(G126), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n523), .A2(n541), .ZN(n543) );
  NAND2_X1 U599 ( .A1(G114), .A2(n895), .ZN(n542) );
  AND2_X1 U600 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U601 ( .A1(n800), .A2(G89), .ZN(n547) );
  XNOR2_X1 U602 ( .A(n547), .B(KEYINPUT4), .ZN(n549) );
  XOR2_X1 U603 ( .A(G543), .B(KEYINPUT0), .Z(n572) );
  INV_X1 U604 ( .A(G651), .ZN(n551) );
  NOR2_X1 U605 ( .A1(n572), .A2(n551), .ZN(n801) );
  NAND2_X1 U606 ( .A1(G76), .A2(n801), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U608 ( .A(KEYINPUT5), .B(n550), .ZN(n559) );
  NOR2_X1 U609 ( .A1(G543), .A2(n551), .ZN(n552) );
  XOR2_X2 U610 ( .A(KEYINPUT1), .B(n552), .Z(n796) );
  NAND2_X1 U611 ( .A1(n796), .A2(G63), .ZN(n553) );
  XOR2_X1 U612 ( .A(KEYINPUT71), .B(n553), .Z(n556) );
  NOR2_X1 U613 ( .A1(G651), .A2(n572), .ZN(n554) );
  XNOR2_X1 U614 ( .A(KEYINPUT66), .B(n554), .ZN(n797) );
  NAND2_X1 U615 ( .A1(G51), .A2(n797), .ZN(n555) );
  NAND2_X1 U616 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U617 ( .A(KEYINPUT6), .B(n557), .Z(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U619 ( .A(KEYINPUT7), .B(n560), .ZN(G168) );
  NAND2_X1 U620 ( .A1(n800), .A2(G90), .ZN(n561) );
  XNOR2_X1 U621 ( .A(n561), .B(KEYINPUT68), .ZN(n563) );
  NAND2_X1 U622 ( .A1(G77), .A2(n801), .ZN(n562) );
  NAND2_X1 U623 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U624 ( .A(KEYINPUT9), .B(n564), .ZN(n568) );
  NAND2_X1 U625 ( .A1(n797), .A2(G52), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G64), .A2(n796), .ZN(n565) );
  AND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n568), .A2(n567), .ZN(G301) );
  INV_X1 U629 ( .A(G301), .ZN(G171) );
  NAND2_X1 U630 ( .A1(G651), .A2(G74), .ZN(n570) );
  NAND2_X1 U631 ( .A1(G49), .A2(n797), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U633 ( .A1(n796), .A2(n571), .ZN(n574) );
  NAND2_X1 U634 ( .A1(n572), .A2(G87), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(G288) );
  XOR2_X1 U636 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U637 ( .A1(G88), .A2(n800), .ZN(n576) );
  NAND2_X1 U638 ( .A1(G75), .A2(n801), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U640 ( .A1(G62), .A2(n796), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G50), .A2(n797), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U643 ( .A1(n580), .A2(n579), .ZN(G166) );
  INV_X1 U644 ( .A(G166), .ZN(G303) );
  NAND2_X1 U645 ( .A1(n797), .A2(G48), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT78), .ZN(n590) );
  NAND2_X1 U647 ( .A1(G73), .A2(n801), .ZN(n582) );
  XOR2_X1 U648 ( .A(KEYINPUT2), .B(n582), .Z(n583) );
  XNOR2_X1 U649 ( .A(n583), .B(KEYINPUT77), .ZN(n585) );
  NAND2_X1 U650 ( .A1(G61), .A2(n796), .ZN(n584) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U652 ( .A1(n800), .A2(G86), .ZN(n586) );
  XOR2_X1 U653 ( .A(KEYINPUT76), .B(n586), .Z(n587) );
  NOR2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U655 ( .A1(n590), .A2(n589), .ZN(G305) );
  AND2_X1 U656 ( .A1(n796), .A2(G60), .ZN(n594) );
  NAND2_X1 U657 ( .A1(G85), .A2(n800), .ZN(n592) );
  NAND2_X1 U658 ( .A1(G72), .A2(n801), .ZN(n591) );
  NAND2_X1 U659 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U660 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U661 ( .A1(G47), .A2(n797), .ZN(n595) );
  NAND2_X1 U662 ( .A1(n596), .A2(n595), .ZN(G290) );
  NAND2_X1 U663 ( .A1(G160), .A2(G40), .ZN(n703) );
  NOR2_X1 U664 ( .A1(n720), .A2(G1966), .ZN(n663) );
  NOR2_X1 U665 ( .A1(G2084), .A2(n672), .ZN(n662) );
  NOR2_X1 U666 ( .A1(n663), .A2(n662), .ZN(n598) );
  XNOR2_X1 U667 ( .A(KEYINPUT94), .B(n598), .ZN(n599) );
  NAND2_X1 U668 ( .A1(n599), .A2(G8), .ZN(n600) );
  XNOR2_X1 U669 ( .A(n600), .B(KEYINPUT30), .ZN(n601) );
  NOR2_X1 U670 ( .A1(n601), .A2(G168), .ZN(n606) );
  XNOR2_X1 U671 ( .A(KEYINPUT91), .B(G1961), .ZN(n1025) );
  NAND2_X1 U672 ( .A1(n672), .A2(n1025), .ZN(n603) );
  XNOR2_X1 U673 ( .A(G2078), .B(KEYINPUT25), .ZN(n991) );
  NAND2_X1 U674 ( .A1(n642), .A2(n991), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(n610) );
  OR2_X1 U676 ( .A1(n610), .A2(G171), .ZN(n604) );
  XNOR2_X1 U677 ( .A(n604), .B(KEYINPUT95), .ZN(n605) );
  NOR2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n609) );
  XNOR2_X1 U679 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n607) );
  XNOR2_X1 U680 ( .A(n607), .B(KEYINPUT31), .ZN(n608) );
  XNOR2_X1 U681 ( .A(n609), .B(n608), .ZN(n670) );
  NAND2_X1 U682 ( .A1(n610), .A2(G171), .ZN(n661) );
  INV_X1 U683 ( .A(G1996), .ZN(n984) );
  NOR2_X1 U684 ( .A1(n672), .A2(n984), .ZN(n611) );
  XNOR2_X1 U685 ( .A(n611), .B(KEYINPUT26), .ZN(n625) );
  AND2_X1 U686 ( .A1(n672), .A2(G1341), .ZN(n623) );
  NAND2_X1 U687 ( .A1(n800), .A2(G81), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n612), .B(KEYINPUT12), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G68), .A2(n801), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U691 ( .A(KEYINPUT13), .B(n615), .Z(n619) );
  NAND2_X1 U692 ( .A1(G56), .A2(n796), .ZN(n616) );
  XNOR2_X1 U693 ( .A(n616), .B(KEYINPUT14), .ZN(n617) );
  XNOR2_X1 U694 ( .A(n617), .B(KEYINPUT69), .ZN(n618) );
  XNOR2_X1 U695 ( .A(n620), .B(KEYINPUT70), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G43), .A2(n797), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n973) );
  NOR2_X2 U698 ( .A1(n625), .A2(n624), .ZN(n638) );
  NAND2_X1 U699 ( .A1(G92), .A2(n800), .ZN(n627) );
  NAND2_X1 U700 ( .A1(G79), .A2(n801), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U702 ( .A1(G66), .A2(n796), .ZN(n629) );
  NAND2_X1 U703 ( .A1(G54), .A2(n797), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U706 ( .A(KEYINPUT15), .B(n632), .Z(n918) );
  NAND2_X1 U707 ( .A1(n638), .A2(n918), .ZN(n637) );
  NAND2_X1 U708 ( .A1(G1348), .A2(n672), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G2067), .A2(n642), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U711 ( .A(KEYINPUT93), .B(n635), .Z(n636) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n640) );
  OR2_X1 U713 ( .A1(n918), .A2(n638), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n652) );
  NAND2_X1 U715 ( .A1(n642), .A2(G2072), .ZN(n641) );
  XNOR2_X1 U716 ( .A(n641), .B(KEYINPUT27), .ZN(n644) );
  INV_X1 U717 ( .A(G1956), .ZN(n1016) );
  NOR2_X1 U718 ( .A1(n1016), .A2(n642), .ZN(n643) );
  NOR2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n653) );
  NAND2_X1 U720 ( .A1(G65), .A2(n796), .ZN(n646) );
  NAND2_X1 U721 ( .A1(G53), .A2(n797), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n646), .A2(n645), .ZN(n650) );
  NAND2_X1 U723 ( .A1(G91), .A2(n800), .ZN(n648) );
  NAND2_X1 U724 ( .A1(G78), .A2(n801), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n956) );
  NAND2_X1 U727 ( .A1(n653), .A2(n956), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n652), .A2(n651), .ZN(n657) );
  NOR2_X1 U729 ( .A1(n653), .A2(n956), .ZN(n655) );
  XOR2_X1 U730 ( .A(KEYINPUT28), .B(KEYINPUT92), .Z(n654) );
  XNOR2_X1 U731 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U733 ( .A(KEYINPUT29), .B(n658), .ZN(n659) );
  INV_X1 U734 ( .A(n659), .ZN(n660) );
  NAND2_X1 U735 ( .A1(n661), .A2(n660), .ZN(n669) );
  AND2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n666) );
  AND2_X1 U737 ( .A1(G8), .A2(n662), .ZN(n664) );
  OR2_X1 U738 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U739 ( .A1(G1976), .A2(G288), .ZN(n967) );
  INV_X1 U740 ( .A(n967), .ZN(n667) );
  OR2_X1 U741 ( .A1(n720), .A2(n667), .ZN(n687) );
  INV_X1 U742 ( .A(n687), .ZN(n668) );
  AND2_X1 U743 ( .A1(n712), .A2(n668), .ZN(n683) );
  NAND2_X1 U744 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U745 ( .A1(n671), .A2(G286), .ZN(n680) );
  INV_X1 U746 ( .A(G8), .ZN(n678) );
  NOR2_X1 U747 ( .A1(G1971), .A2(n720), .ZN(n674) );
  NOR2_X1 U748 ( .A1(G2090), .A2(n672), .ZN(n673) );
  NOR2_X1 U749 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U750 ( .A(n675), .B(KEYINPUT98), .ZN(n676) );
  NAND2_X1 U751 ( .A1(n676), .A2(G303), .ZN(n677) );
  OR2_X1 U752 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U753 ( .A(KEYINPUT99), .B(KEYINPUT32), .Z(n681) );
  NAND2_X1 U754 ( .A1(n683), .A2(n711), .ZN(n689) );
  NOR2_X1 U755 ( .A1(G1976), .A2(G288), .ZN(n965) );
  NOR2_X1 U756 ( .A1(G1971), .A2(G303), .ZN(n684) );
  NOR2_X1 U757 ( .A1(n965), .A2(n684), .ZN(n685) );
  XNOR2_X1 U758 ( .A(n685), .B(KEYINPUT100), .ZN(n686) );
  OR2_X1 U759 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U760 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U761 ( .A(n690), .B(KEYINPUT64), .ZN(n691) );
  NOR2_X1 U762 ( .A1(KEYINPUT33), .A2(n691), .ZN(n692) );
  INV_X1 U763 ( .A(n692), .ZN(n710) );
  XOR2_X1 U764 ( .A(G1981), .B(G305), .Z(n962) );
  XOR2_X1 U765 ( .A(KEYINPUT37), .B(G2067), .Z(n762) );
  NAND2_X1 U766 ( .A1(G128), .A2(n894), .ZN(n694) );
  NAND2_X1 U767 ( .A1(G116), .A2(n895), .ZN(n693) );
  NAND2_X1 U768 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U769 ( .A(n695), .B(KEYINPUT35), .ZN(n700) );
  NAND2_X1 U770 ( .A1(G140), .A2(n890), .ZN(n697) );
  NAND2_X1 U771 ( .A1(G104), .A2(n891), .ZN(n696) );
  NAND2_X1 U772 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U773 ( .A(KEYINPUT34), .B(n698), .Z(n699) );
  NAND2_X1 U774 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U775 ( .A(n701), .B(KEYINPUT36), .ZN(n903) );
  NAND2_X1 U776 ( .A1(n762), .A2(n903), .ZN(n933) );
  NOR2_X1 U777 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U778 ( .A(KEYINPUT85), .B(n705), .ZN(n728) );
  NOR2_X1 U779 ( .A1(n933), .A2(n728), .ZN(n724) );
  INV_X1 U780 ( .A(n724), .ZN(n706) );
  AND2_X1 U781 ( .A1(n962), .A2(n706), .ZN(n708) );
  NAND2_X1 U782 ( .A1(n965), .A2(KEYINPUT33), .ZN(n707) );
  NAND2_X1 U783 ( .A1(n710), .A2(n709), .ZN(n727) );
  NAND2_X1 U784 ( .A1(n712), .A2(n711), .ZN(n715) );
  NOR2_X1 U785 ( .A1(G2090), .A2(G303), .ZN(n713) );
  NAND2_X1 U786 ( .A1(G8), .A2(n713), .ZN(n714) );
  NAND2_X1 U787 ( .A1(n715), .A2(n714), .ZN(n716) );
  AND2_X1 U788 ( .A1(n716), .A2(n720), .ZN(n722) );
  NOR2_X1 U789 ( .A1(G1981), .A2(G305), .ZN(n717) );
  XOR2_X1 U790 ( .A(n717), .B(KEYINPUT90), .Z(n718) );
  XNOR2_X1 U791 ( .A(KEYINPUT24), .B(n718), .ZN(n719) );
  NOR2_X1 U792 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U793 ( .A1(n722), .A2(n721), .ZN(n723) );
  INV_X1 U794 ( .A(n725), .ZN(n726) );
  NAND2_X1 U795 ( .A1(n727), .A2(n726), .ZN(n748) );
  INV_X1 U796 ( .A(n728), .ZN(n766) );
  XNOR2_X1 U797 ( .A(KEYINPUT88), .B(n766), .ZN(n746) );
  NAND2_X1 U798 ( .A1(G131), .A2(n890), .ZN(n730) );
  NAND2_X1 U799 ( .A1(G119), .A2(n894), .ZN(n729) );
  NAND2_X1 U800 ( .A1(n730), .A2(n729), .ZN(n734) );
  NAND2_X1 U801 ( .A1(G95), .A2(n891), .ZN(n732) );
  NAND2_X1 U802 ( .A1(G107), .A2(n895), .ZN(n731) );
  NAND2_X1 U803 ( .A1(n732), .A2(n731), .ZN(n733) );
  OR2_X1 U804 ( .A1(n734), .A2(n733), .ZN(n902) );
  NAND2_X1 U805 ( .A1(G1991), .A2(n902), .ZN(n745) );
  XOR2_X1 U806 ( .A(KEYINPUT86), .B(KEYINPUT38), .Z(n736) );
  NAND2_X1 U807 ( .A1(G105), .A2(n891), .ZN(n735) );
  XNOR2_X1 U808 ( .A(n736), .B(n735), .ZN(n740) );
  NAND2_X1 U809 ( .A1(G129), .A2(n894), .ZN(n738) );
  NAND2_X1 U810 ( .A1(G117), .A2(n895), .ZN(n737) );
  NAND2_X1 U811 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U812 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U813 ( .A(KEYINPUT87), .B(n741), .Z(n743) );
  NAND2_X1 U814 ( .A1(n890), .A2(G141), .ZN(n742) );
  NAND2_X1 U815 ( .A1(n743), .A2(n742), .ZN(n908) );
  NAND2_X1 U816 ( .A1(G1996), .A2(n908), .ZN(n744) );
  NAND2_X1 U817 ( .A1(n745), .A2(n744), .ZN(n936) );
  NAND2_X1 U818 ( .A1(n746), .A2(n936), .ZN(n747) );
  XOR2_X1 U819 ( .A(KEYINPUT89), .B(n747), .Z(n753) );
  NAND2_X1 U820 ( .A1(n748), .A2(n753), .ZN(n749) );
  XNOR2_X1 U821 ( .A(n749), .B(KEYINPUT101), .ZN(n751) );
  XNOR2_X1 U822 ( .A(G1986), .B(G290), .ZN(n959) );
  NAND2_X1 U823 ( .A1(n766), .A2(n959), .ZN(n750) );
  NAND2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U825 ( .A(n752), .B(KEYINPUT102), .ZN(n768) );
  NOR2_X1 U826 ( .A1(G1996), .A2(n908), .ZN(n945) );
  INV_X1 U827 ( .A(n753), .ZN(n757) );
  NOR2_X1 U828 ( .A1(G1991), .A2(n902), .ZN(n938) );
  NOR2_X1 U829 ( .A1(G1986), .A2(G290), .ZN(n754) );
  NOR2_X1 U830 ( .A1(n938), .A2(n754), .ZN(n755) );
  XOR2_X1 U831 ( .A(KEYINPUT103), .B(n755), .Z(n756) );
  NOR2_X1 U832 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U833 ( .A1(n945), .A2(n758), .ZN(n759) );
  XNOR2_X1 U834 ( .A(n759), .B(KEYINPUT39), .ZN(n760) );
  NAND2_X1 U835 ( .A1(n760), .A2(n933), .ZN(n761) );
  XNOR2_X1 U836 ( .A(n761), .B(KEYINPUT104), .ZN(n764) );
  NOR2_X1 U837 ( .A1(n903), .A2(n762), .ZN(n763) );
  XNOR2_X1 U838 ( .A(n763), .B(KEYINPUT105), .ZN(n950) );
  NAND2_X1 U839 ( .A1(n764), .A2(n950), .ZN(n765) );
  NAND2_X1 U840 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U841 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U842 ( .A(n769), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U843 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U844 ( .A(G57), .ZN(G237) );
  INV_X1 U845 ( .A(G132), .ZN(G219) );
  INV_X1 U846 ( .A(G82), .ZN(G220) );
  NAND2_X1 U847 ( .A1(G7), .A2(G661), .ZN(n770) );
  XNOR2_X1 U848 ( .A(n770), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U849 ( .A(G223), .ZN(n847) );
  NAND2_X1 U850 ( .A1(n847), .A2(G567), .ZN(n771) );
  XOR2_X1 U851 ( .A(KEYINPUT11), .B(n771), .Z(G234) );
  INV_X1 U852 ( .A(n973), .ZN(n772) );
  NAND2_X1 U853 ( .A1(n772), .A2(G860), .ZN(G153) );
  NAND2_X1 U854 ( .A1(G868), .A2(G301), .ZN(n774) );
  INV_X1 U855 ( .A(n918), .ZN(n957) );
  INV_X1 U856 ( .A(G868), .ZN(n818) );
  NAND2_X1 U857 ( .A1(n957), .A2(n818), .ZN(n773) );
  NAND2_X1 U858 ( .A1(n774), .A2(n773), .ZN(G284) );
  INV_X1 U859 ( .A(n956), .ZN(G299) );
  XNOR2_X1 U860 ( .A(KEYINPUT72), .B(n818), .ZN(n775) );
  NOR2_X1 U861 ( .A1(G286), .A2(n775), .ZN(n777) );
  NOR2_X1 U862 ( .A1(G868), .A2(G299), .ZN(n776) );
  NOR2_X1 U863 ( .A1(n777), .A2(n776), .ZN(G297) );
  INV_X1 U864 ( .A(G559), .ZN(n778) );
  NOR2_X1 U865 ( .A1(G860), .A2(n778), .ZN(n779) );
  XNOR2_X1 U866 ( .A(KEYINPUT73), .B(n779), .ZN(n780) );
  NAND2_X1 U867 ( .A1(n780), .A2(n918), .ZN(n781) );
  XNOR2_X1 U868 ( .A(n781), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U869 ( .A1(G868), .A2(n973), .ZN(n784) );
  NAND2_X1 U870 ( .A1(G868), .A2(n918), .ZN(n782) );
  NOR2_X1 U871 ( .A1(G559), .A2(n782), .ZN(n783) );
  NOR2_X1 U872 ( .A1(n784), .A2(n783), .ZN(G282) );
  NAND2_X1 U873 ( .A1(G123), .A2(n894), .ZN(n785) );
  XNOR2_X1 U874 ( .A(n785), .B(KEYINPUT18), .ZN(n786) );
  XNOR2_X1 U875 ( .A(n786), .B(KEYINPUT74), .ZN(n788) );
  NAND2_X1 U876 ( .A1(G99), .A2(n891), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n792) );
  NAND2_X1 U878 ( .A1(G135), .A2(n890), .ZN(n790) );
  NAND2_X1 U879 ( .A1(G111), .A2(n895), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n937) );
  XOR2_X1 U882 ( .A(n937), .B(G2096), .Z(n793) );
  NOR2_X1 U883 ( .A1(G2100), .A2(n793), .ZN(n794) );
  XNOR2_X1 U884 ( .A(KEYINPUT75), .B(n794), .ZN(G156) );
  NAND2_X1 U885 ( .A1(n918), .A2(G559), .ZN(n815) );
  XNOR2_X1 U886 ( .A(n973), .B(n815), .ZN(n795) );
  NOR2_X1 U887 ( .A1(n795), .A2(G860), .ZN(n806) );
  NAND2_X1 U888 ( .A1(G67), .A2(n796), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G55), .A2(n797), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n805) );
  NAND2_X1 U891 ( .A1(G93), .A2(n800), .ZN(n803) );
  NAND2_X1 U892 ( .A1(G80), .A2(n801), .ZN(n802) );
  NAND2_X1 U893 ( .A1(n803), .A2(n802), .ZN(n804) );
  OR2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n817) );
  XOR2_X1 U895 ( .A(n806), .B(n817), .Z(G145) );
  XNOR2_X1 U896 ( .A(KEYINPUT79), .B(KEYINPUT80), .ZN(n808) );
  XNOR2_X1 U897 ( .A(G288), .B(KEYINPUT19), .ZN(n807) );
  XNOR2_X1 U898 ( .A(n808), .B(n807), .ZN(n809) );
  XNOR2_X1 U899 ( .A(G305), .B(n809), .ZN(n811) );
  XNOR2_X1 U900 ( .A(n956), .B(G166), .ZN(n810) );
  XNOR2_X1 U901 ( .A(n811), .B(n810), .ZN(n812) );
  XNOR2_X1 U902 ( .A(n817), .B(n812), .ZN(n813) );
  XNOR2_X1 U903 ( .A(G290), .B(n813), .ZN(n814) );
  XNOR2_X1 U904 ( .A(n814), .B(n973), .ZN(n915) );
  XNOR2_X1 U905 ( .A(n815), .B(n915), .ZN(n816) );
  NAND2_X1 U906 ( .A1(n816), .A2(G868), .ZN(n820) );
  NAND2_X1 U907 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U908 ( .A1(n820), .A2(n819), .ZN(G295) );
  NAND2_X1 U909 ( .A1(G2084), .A2(G2078), .ZN(n821) );
  XOR2_X1 U910 ( .A(KEYINPUT20), .B(n821), .Z(n822) );
  NAND2_X1 U911 ( .A1(G2090), .A2(n822), .ZN(n823) );
  XNOR2_X1 U912 ( .A(KEYINPUT21), .B(n823), .ZN(n824) );
  NAND2_X1 U913 ( .A1(n824), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U914 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U915 ( .A1(G220), .A2(G219), .ZN(n825) );
  XOR2_X1 U916 ( .A(KEYINPUT22), .B(n825), .Z(n826) );
  NOR2_X1 U917 ( .A1(G218), .A2(n826), .ZN(n827) );
  NAND2_X1 U918 ( .A1(G96), .A2(n827), .ZN(n851) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n851), .ZN(n831) );
  NAND2_X1 U920 ( .A1(G69), .A2(G120), .ZN(n828) );
  NOR2_X1 U921 ( .A1(G237), .A2(n828), .ZN(n829) );
  NAND2_X1 U922 ( .A1(G108), .A2(n829), .ZN(n852) );
  NAND2_X1 U923 ( .A1(G567), .A2(n852), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U925 ( .A(KEYINPUT81), .B(n832), .ZN(G319) );
  INV_X1 U926 ( .A(G319), .ZN(n834) );
  NAND2_X1 U927 ( .A1(G661), .A2(G483), .ZN(n833) );
  NOR2_X1 U928 ( .A1(n834), .A2(n833), .ZN(n850) );
  NAND2_X1 U929 ( .A1(n850), .A2(G36), .ZN(n835) );
  XNOR2_X1 U930 ( .A(KEYINPUT82), .B(n835), .ZN(G176) );
  XNOR2_X1 U931 ( .A(G2427), .B(G2443), .ZN(n845) );
  XOR2_X1 U932 ( .A(G2430), .B(KEYINPUT107), .Z(n837) );
  XNOR2_X1 U933 ( .A(G2454), .B(G2435), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U935 ( .A(G2438), .B(KEYINPUT106), .Z(n839) );
  XNOR2_X1 U936 ( .A(G1341), .B(G1348), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U938 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U939 ( .A(G2446), .B(G2451), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n845), .B(n844), .ZN(n846) );
  NAND2_X1 U942 ( .A1(n846), .A2(G14), .ZN(n921) );
  XOR2_X1 U943 ( .A(KEYINPUT108), .B(n921), .Z(G401) );
  NAND2_X1 U944 ( .A1(G2106), .A2(n847), .ZN(G217) );
  AND2_X1 U945 ( .A1(G15), .A2(G2), .ZN(n848) );
  NAND2_X1 U946 ( .A1(G661), .A2(n848), .ZN(G259) );
  NAND2_X1 U947 ( .A1(G3), .A2(G1), .ZN(n849) );
  NAND2_X1 U948 ( .A1(n850), .A2(n849), .ZN(G188) );
  NOR2_X1 U949 ( .A1(n852), .A2(n851), .ZN(G325) );
  XNOR2_X1 U950 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U952 ( .A(G120), .ZN(G236) );
  INV_X1 U953 ( .A(G96), .ZN(G221) );
  INV_X1 U954 ( .A(G69), .ZN(G235) );
  XOR2_X1 U955 ( .A(G2096), .B(KEYINPUT43), .Z(n854) );
  XNOR2_X1 U956 ( .A(G2090), .B(KEYINPUT110), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U958 ( .A(n855), .B(G2678), .Z(n857) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n856) );
  XNOR2_X1 U960 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U961 ( .A(KEYINPUT42), .B(G2100), .Z(n859) );
  XNOR2_X1 U962 ( .A(G2084), .B(G2078), .ZN(n858) );
  XNOR2_X1 U963 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U964 ( .A(n861), .B(n860), .ZN(G227) );
  XOR2_X1 U965 ( .A(G1976), .B(G1981), .Z(n863) );
  XNOR2_X1 U966 ( .A(G1966), .B(G1956), .ZN(n862) );
  XNOR2_X1 U967 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U968 ( .A(G1971), .B(G1986), .Z(n865) );
  XNOR2_X1 U969 ( .A(G1996), .B(G1991), .ZN(n864) );
  XNOR2_X1 U970 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U971 ( .A(n867), .B(n866), .Z(n869) );
  XNOR2_X1 U972 ( .A(KEYINPUT111), .B(G2474), .ZN(n868) );
  XNOR2_X1 U973 ( .A(n869), .B(n868), .ZN(n871) );
  XOR2_X1 U974 ( .A(G1961), .B(KEYINPUT41), .Z(n870) );
  XNOR2_X1 U975 ( .A(n871), .B(n870), .ZN(G229) );
  NAND2_X1 U976 ( .A1(n894), .A2(G124), .ZN(n873) );
  XNOR2_X1 U977 ( .A(KEYINPUT44), .B(KEYINPUT112), .ZN(n872) );
  XNOR2_X1 U978 ( .A(n873), .B(n872), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G136), .A2(n890), .ZN(n875) );
  NAND2_X1 U980 ( .A1(G100), .A2(n891), .ZN(n874) );
  NAND2_X1 U981 ( .A1(n875), .A2(n874), .ZN(n878) );
  NAND2_X1 U982 ( .A1(G112), .A2(n895), .ZN(n876) );
  XNOR2_X1 U983 ( .A(KEYINPUT113), .B(n876), .ZN(n877) );
  NOR2_X1 U984 ( .A1(n878), .A2(n877), .ZN(n879) );
  NAND2_X1 U985 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U986 ( .A(KEYINPUT114), .B(n881), .Z(G162) );
  NAND2_X1 U987 ( .A1(G130), .A2(n894), .ZN(n883) );
  NAND2_X1 U988 ( .A1(G118), .A2(n895), .ZN(n882) );
  NAND2_X1 U989 ( .A1(n883), .A2(n882), .ZN(n888) );
  NAND2_X1 U990 ( .A1(G142), .A2(n890), .ZN(n885) );
  NAND2_X1 U991 ( .A1(G106), .A2(n891), .ZN(n884) );
  NAND2_X1 U992 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U993 ( .A(KEYINPUT45), .B(n886), .Z(n887) );
  NOR2_X1 U994 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U995 ( .A(G160), .B(n889), .ZN(n912) );
  NAND2_X1 U996 ( .A1(G139), .A2(n890), .ZN(n893) );
  NAND2_X1 U997 ( .A1(G103), .A2(n891), .ZN(n892) );
  NAND2_X1 U998 ( .A1(n893), .A2(n892), .ZN(n901) );
  NAND2_X1 U999 ( .A1(G127), .A2(n894), .ZN(n897) );
  NAND2_X1 U1000 ( .A1(G115), .A2(n895), .ZN(n896) );
  NAND2_X1 U1001 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U1002 ( .A(KEYINPUT47), .B(n898), .ZN(n899) );
  XNOR2_X1 U1003 ( .A(KEYINPUT115), .B(n899), .ZN(n900) );
  NOR2_X1 U1004 ( .A1(n901), .A2(n900), .ZN(n927) );
  XNOR2_X1 U1005 ( .A(n903), .B(n902), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n904) );
  XNOR2_X1 U1007 ( .A(n904), .B(G162), .ZN(n905) );
  XNOR2_X1 U1008 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1009 ( .A(n927), .B(n907), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(n908), .B(n937), .ZN(n909) );
  XNOR2_X1 U1011 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1013 ( .A(n913), .B(G164), .Z(n914) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n914), .ZN(G395) );
  XOR2_X1 U1015 ( .A(KEYINPUT116), .B(n915), .Z(n917) );
  XNOR2_X1 U1016 ( .A(G171), .B(G286), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n917), .B(n916), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n920), .ZN(G397) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n921), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1024 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1026 ( .A(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1028 ( .A(n927), .B(KEYINPUT119), .Z(n928) );
  XOR2_X1 U1029 ( .A(G2072), .B(n928), .Z(n930) );
  XOR2_X1 U1030 ( .A(G164), .B(G2078), .Z(n929) );
  NOR2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1032 ( .A(n931), .B(KEYINPUT120), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(n932), .B(KEYINPUT50), .ZN(n943) );
  XNOR2_X1 U1034 ( .A(G2084), .B(G160), .ZN(n934) );
  NAND2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n940) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(KEYINPUT117), .B(n941), .ZN(n942) );
  NAND2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n949) );
  XOR2_X1 U1041 ( .A(G2090), .B(G162), .Z(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(KEYINPUT118), .B(n946), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(KEYINPUT51), .B(n947), .ZN(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1047 ( .A(KEYINPUT52), .B(n952), .Z(n954) );
  INV_X1 U1048 ( .A(KEYINPUT55), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n955), .A2(G29), .ZN(n1010) );
  XOR2_X1 U1051 ( .A(G16), .B(KEYINPUT56), .Z(n982) );
  XNOR2_X1 U1052 ( .A(n956), .B(G1956), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(G1348), .B(n957), .ZN(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n979) );
  XNOR2_X1 U1056 ( .A(G1966), .B(G168), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(n964), .B(KEYINPUT57), .ZN(n977) );
  INV_X1 U1059 ( .A(n965), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(n968), .B(KEYINPUT125), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(G301), .B(G1961), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(G303), .B(G1971), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(G1341), .B(n973), .ZN(n974) );
  NOR2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(n980), .B(KEYINPUT126), .ZN(n981) );
  NOR2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n1008) );
  XOR2_X1 U1072 ( .A(G29), .B(KEYINPUT124), .Z(n1005) );
  XNOR2_X1 U1073 ( .A(KEYINPUT121), .B(G2090), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(n983), .B(G35), .ZN(n999) );
  XOR2_X1 U1075 ( .A(KEYINPUT123), .B(KEYINPUT53), .Z(n997) );
  XOR2_X1 U1076 ( .A(G2067), .B(G26), .Z(n986) );
  XNOR2_X1 U1077 ( .A(n984), .B(G32), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n990) );
  XOR2_X1 U1079 ( .A(G1991), .B(G25), .Z(n987) );
  NAND2_X1 U1080 ( .A1(n987), .A2(G28), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(KEYINPUT122), .B(n988), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n995) );
  XOR2_X1 U1083 ( .A(n991), .B(G27), .Z(n993) );
  XNOR2_X1 U1084 ( .A(G2072), .B(G33), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(n997), .B(n996), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(G34), .B(G2084), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(KEYINPUT54), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1003), .B(KEYINPUT55), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(G11), .A2(n1006), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1036) );
  XOR2_X1 U1097 ( .A(G1976), .B(G23), .Z(n1012) );
  XOR2_X1 U1098 ( .A(G1971), .B(G22), .Z(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G24), .B(G1986), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT58), .B(n1015), .Z(n1032) );
  XNOR2_X1 U1103 ( .A(G20), .B(n1016), .ZN(n1020) );
  XNOR2_X1 U1104 ( .A(G1341), .B(G19), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(G6), .B(G1981), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1023) );
  XOR2_X1 U1108 ( .A(KEYINPUT59), .B(G1348), .Z(n1021) );
  XNOR2_X1 U1109 ( .A(G4), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1111 ( .A(KEYINPUT60), .B(n1024), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(n1025), .B(G5), .ZN(n1026) );
  NAND2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(G21), .B(G1966), .ZN(n1028) );
  NOR2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1116 ( .A(KEYINPUT127), .B(n1030), .ZN(n1031) );
  NOR2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1118 ( .A(KEYINPUT61), .B(n1033), .Z(n1034) );
  NOR2_X1 U1119 ( .A1(G16), .A2(n1034), .ZN(n1035) );
  NOR2_X1 U1120 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XNOR2_X1 U1121 ( .A(n1037), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1122 ( .A(G311), .ZN(G150) );
endmodule

