

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U551 ( .A1(n750), .A2(n749), .ZN(n752) );
  XNOR2_X1 U552 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n523) );
  AND2_X2 U553 ( .A1(n537), .A2(n536), .ZN(n683) );
  AND2_X1 U554 ( .A1(n830), .A2(n521), .ZN(n831) );
  NOR2_X1 U555 ( .A1(G164), .A2(G1384), .ZN(n684) );
  BUF_X1 U556 ( .A(n588), .Z(n540) );
  BUF_X1 U557 ( .A(n615), .Z(n616) );
  NOR2_X2 U558 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X2 U559 ( .A1(n683), .A2(G40), .ZN(n797) );
  NOR2_X2 U560 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U561 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U562 ( .A1(G1966), .A2(n778), .ZN(n729) );
  OR2_X1 U563 ( .A1(n767), .A2(n519), .ZN(n757) );
  INV_X2 U564 ( .A(G2105), .ZN(n526) );
  XOR2_X1 U565 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  NOR2_X1 U566 ( .A1(n591), .A2(n590), .ZN(n593) );
  NOR2_X1 U567 ( .A1(n778), .A2(n763), .ZN(n517) );
  NAND2_X1 U568 ( .A1(n764), .A2(KEYINPUT33), .ZN(n518) );
  XOR2_X1 U569 ( .A(KEYINPUT100), .B(n955), .Z(n519) );
  AND2_X1 U570 ( .A1(n615), .A2(G137), .ZN(n520) );
  NAND2_X1 U571 ( .A1(n829), .A2(n828), .ZN(n521) );
  INV_X1 U572 ( .A(KEYINPUT27), .ZN(n702) );
  XNOR2_X1 U573 ( .A(n703), .B(n702), .ZN(n705) );
  XNOR2_X1 U574 ( .A(KEYINPUT96), .B(KEYINPUT30), .ZN(n722) );
  INV_X1 U575 ( .A(KEYINPUT95), .ZN(n709) );
  INV_X1 U576 ( .A(KEYINPUT32), .ZN(n751) );
  XNOR2_X1 U577 ( .A(n752), .B(n751), .ZN(n753) );
  BUF_X1 U578 ( .A(n695), .Z(n736) );
  XNOR2_X1 U579 ( .A(KEYINPUT76), .B(KEYINPUT12), .ZN(n582) );
  XNOR2_X1 U580 ( .A(n583), .B(n582), .ZN(n585) );
  NOR2_X2 U581 ( .A1(n634), .A2(n544), .ZN(n645) );
  NAND2_X1 U582 ( .A1(n593), .A2(n592), .ZN(n959) );
  NOR2_X1 U583 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XNOR2_X1 U584 ( .A(n523), .B(n522), .ZN(n615) );
  NAND2_X1 U585 ( .A1(n615), .A2(G138), .ZN(n525) );
  AND2_X4 U586 ( .A1(n526), .A2(G2104), .ZN(n534) );
  NAND2_X1 U587 ( .A1(G102), .A2(n534), .ZN(n524) );
  NAND2_X1 U588 ( .A1(n525), .A2(n524), .ZN(n530) );
  NOR2_X4 U589 ( .A1(G2104), .A2(n526), .ZN(n888) );
  NAND2_X1 U590 ( .A1(G126), .A2(n888), .ZN(n528) );
  AND2_X1 U591 ( .A1(G2105), .A2(G2104), .ZN(n886) );
  NAND2_X1 U592 ( .A1(G114), .A2(n886), .ZN(n527) );
  NAND2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X2 U594 ( .A1(n530), .A2(n529), .ZN(G164) );
  NAND2_X1 U595 ( .A1(G125), .A2(n888), .ZN(n532) );
  NAND2_X1 U596 ( .A1(G113), .A2(n886), .ZN(n531) );
  NAND2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U598 ( .A1(n533), .A2(n520), .ZN(n537) );
  NAND2_X1 U599 ( .A1(G101), .A2(n534), .ZN(n535) );
  XOR2_X1 U600 ( .A(KEYINPUT23), .B(n535), .Z(n536) );
  BUF_X1 U601 ( .A(n683), .Z(G160) );
  INV_X1 U602 ( .A(G651), .ZN(n544) );
  NOR2_X1 U603 ( .A1(G543), .A2(n544), .ZN(n539) );
  XOR2_X1 U604 ( .A(KEYINPUT1), .B(n539), .Z(n588) );
  NAND2_X1 U605 ( .A1(G64), .A2(n540), .ZN(n543) );
  NOR2_X1 U606 ( .A1(G651), .A2(n634), .ZN(n541) );
  XNOR2_X2 U607 ( .A(KEYINPUT66), .B(n541), .ZN(n646) );
  NAND2_X1 U608 ( .A1(G52), .A2(n646), .ZN(n542) );
  NAND2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n551) );
  XNOR2_X1 U610 ( .A(KEYINPUT9), .B(KEYINPUT70), .ZN(n549) );
  NAND2_X1 U611 ( .A1(n649), .A2(G90), .ZN(n547) );
  NAND2_X1 U612 ( .A1(n645), .A2(G77), .ZN(n545) );
  XOR2_X1 U613 ( .A(KEYINPUT69), .B(n545), .Z(n546) );
  NAND2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U615 ( .A(n549), .B(n548), .Z(n550) );
  NOR2_X1 U616 ( .A1(n551), .A2(n550), .ZN(G171) );
  INV_X1 U617 ( .A(G57), .ZN(G237) );
  INV_X1 U618 ( .A(G82), .ZN(G220) );
  NAND2_X1 U619 ( .A1(G88), .A2(n649), .ZN(n553) );
  NAND2_X1 U620 ( .A1(G75), .A2(n645), .ZN(n552) );
  NAND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n540), .A2(G62), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n554), .B(KEYINPUT82), .ZN(n556) );
  NAND2_X1 U624 ( .A1(G50), .A2(n646), .ZN(n555) );
  NAND2_X1 U625 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U626 ( .A1(n558), .A2(n557), .ZN(G166) );
  NAND2_X1 U627 ( .A1(G53), .A2(n646), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n559), .B(KEYINPUT72), .ZN(n561) );
  NAND2_X1 U629 ( .A1(G65), .A2(n540), .ZN(n560) );
  NAND2_X1 U630 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U631 ( .A(KEYINPUT73), .B(n562), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G91), .A2(n649), .ZN(n564) );
  NAND2_X1 U633 ( .A1(G78), .A2(n645), .ZN(n563) );
  AND2_X1 U634 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U635 ( .A1(n566), .A2(n565), .ZN(G299) );
  NAND2_X1 U636 ( .A1(G63), .A2(n540), .ZN(n568) );
  NAND2_X1 U637 ( .A1(G51), .A2(n646), .ZN(n567) );
  NAND2_X1 U638 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U639 ( .A(KEYINPUT6), .B(n569), .Z(n577) );
  NAND2_X1 U640 ( .A1(n645), .A2(G76), .ZN(n570) );
  XNOR2_X1 U641 ( .A(KEYINPUT79), .B(n570), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n649), .A2(G89), .ZN(n571) );
  XOR2_X1 U643 ( .A(n571), .B(KEYINPUT4), .Z(n572) );
  NOR2_X1 U644 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U645 ( .A(KEYINPUT5), .B(n574), .Z(n575) );
  XNOR2_X1 U646 ( .A(KEYINPUT80), .B(n575), .ZN(n576) );
  NAND2_X1 U647 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U648 ( .A(KEYINPUT7), .B(n578), .ZN(G168) );
  XOR2_X1 U649 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U650 ( .A1(G94), .A2(G452), .ZN(n579) );
  XNOR2_X1 U651 ( .A(n579), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U652 ( .A1(G7), .A2(G661), .ZN(n580) );
  XNOR2_X1 U653 ( .A(n580), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U654 ( .A(G223), .B(KEYINPUT75), .ZN(n832) );
  NAND2_X1 U655 ( .A1(n832), .A2(G567), .ZN(n581) );
  XOR2_X1 U656 ( .A(KEYINPUT11), .B(n581), .Z(G234) );
  XNOR2_X1 U657 ( .A(KEYINPUT13), .B(KEYINPUT77), .ZN(n587) );
  NAND2_X1 U658 ( .A1(G81), .A2(n649), .ZN(n583) );
  NAND2_X1 U659 ( .A1(G68), .A2(n645), .ZN(n584) );
  NAND2_X1 U660 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U661 ( .A(n587), .B(n586), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n588), .A2(G56), .ZN(n589) );
  XOR2_X1 U663 ( .A(KEYINPUT14), .B(n589), .Z(n590) );
  NAND2_X1 U664 ( .A1(G43), .A2(n646), .ZN(n592) );
  INV_X1 U665 ( .A(G860), .ZN(n606) );
  OR2_X1 U666 ( .A1(n959), .A2(n606), .ZN(G153) );
  INV_X1 U667 ( .A(G171), .ZN(G301) );
  NAND2_X1 U668 ( .A1(G868), .A2(G301), .ZN(n603) );
  NAND2_X1 U669 ( .A1(n646), .A2(G54), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G92), .A2(n649), .ZN(n595) );
  NAND2_X1 U671 ( .A1(G66), .A2(n540), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n645), .A2(G79), .ZN(n596) );
  XOR2_X1 U674 ( .A(KEYINPUT78), .B(n596), .Z(n597) );
  NOR2_X1 U675 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X2 U677 ( .A(n601), .B(KEYINPUT15), .ZN(n958) );
  OR2_X1 U678 ( .A1(n958), .A2(G868), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n603), .A2(n602), .ZN(G284) );
  INV_X1 U680 ( .A(G868), .ZN(n665) );
  NOR2_X1 U681 ( .A1(G286), .A2(n665), .ZN(n605) );
  NOR2_X1 U682 ( .A1(G868), .A2(G299), .ZN(n604) );
  NOR2_X1 U683 ( .A1(n605), .A2(n604), .ZN(G297) );
  NAND2_X1 U684 ( .A1(n606), .A2(G559), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n607), .A2(n958), .ZN(n608) );
  XNOR2_X1 U686 ( .A(n608), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U687 ( .A1(G868), .A2(n959), .ZN(n611) );
  NAND2_X1 U688 ( .A1(G868), .A2(n958), .ZN(n609) );
  NOR2_X1 U689 ( .A1(G559), .A2(n609), .ZN(n610) );
  NOR2_X1 U690 ( .A1(n611), .A2(n610), .ZN(G282) );
  NAND2_X1 U691 ( .A1(G123), .A2(n888), .ZN(n612) );
  XNOR2_X1 U692 ( .A(n612), .B(KEYINPUT18), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n534), .A2(G99), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n620) );
  NAND2_X1 U695 ( .A1(G135), .A2(n616), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G111), .A2(n886), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n928) );
  XNOR2_X1 U699 ( .A(G2096), .B(n928), .ZN(n622) );
  INV_X1 U700 ( .A(G2100), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(G156) );
  NAND2_X1 U702 ( .A1(n958), .A2(G559), .ZN(n662) );
  XNOR2_X1 U703 ( .A(n959), .B(n662), .ZN(n623) );
  NOR2_X1 U704 ( .A1(n623), .A2(G860), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G93), .A2(n649), .ZN(n625) );
  NAND2_X1 U706 ( .A1(G80), .A2(n645), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G67), .A2(n540), .ZN(n627) );
  NAND2_X1 U709 ( .A1(G55), .A2(n646), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n628) );
  OR2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n664) );
  XOR2_X1 U712 ( .A(n630), .B(n664), .Z(G145) );
  NAND2_X1 U713 ( .A1(G651), .A2(G74), .ZN(n632) );
  NAND2_X1 U714 ( .A1(G49), .A2(n646), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U716 ( .A1(n540), .A2(n633), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n634), .A2(G87), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U719 ( .A1(G73), .A2(n645), .ZN(n637) );
  XOR2_X1 U720 ( .A(KEYINPUT2), .B(n637), .Z(n642) );
  NAND2_X1 U721 ( .A1(G86), .A2(n649), .ZN(n639) );
  NAND2_X1 U722 ( .A1(G61), .A2(n540), .ZN(n638) );
  NAND2_X1 U723 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U724 ( .A(KEYINPUT81), .B(n640), .Z(n641) );
  NOR2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U726 ( .A1(G48), .A2(n646), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n644), .A2(n643), .ZN(G305) );
  NAND2_X1 U728 ( .A1(G72), .A2(n645), .ZN(n648) );
  NAND2_X1 U729 ( .A1(G47), .A2(n646), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U731 ( .A1(G85), .A2(n649), .ZN(n650) );
  XOR2_X1 U732 ( .A(KEYINPUT68), .B(n650), .Z(n651) );
  NOR2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U734 ( .A1(n540), .A2(G60), .ZN(n653) );
  NAND2_X1 U735 ( .A1(n654), .A2(n653), .ZN(G290) );
  XNOR2_X1 U736 ( .A(KEYINPUT83), .B(n959), .ZN(n655) );
  XNOR2_X1 U737 ( .A(n655), .B(G288), .ZN(n656) );
  XNOR2_X1 U738 ( .A(KEYINPUT19), .B(n656), .ZN(n658) );
  XNOR2_X1 U739 ( .A(G305), .B(G166), .ZN(n657) );
  XNOR2_X1 U740 ( .A(n658), .B(n657), .ZN(n659) );
  XOR2_X1 U741 ( .A(n664), .B(n659), .Z(n660) );
  XNOR2_X1 U742 ( .A(n660), .B(G290), .ZN(n661) );
  XNOR2_X1 U743 ( .A(G299), .B(n661), .ZN(n904) );
  XNOR2_X1 U744 ( .A(n662), .B(n904), .ZN(n663) );
  NAND2_X1 U745 ( .A1(n663), .A2(G868), .ZN(n667) );
  NAND2_X1 U746 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U747 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U752 ( .A1(n671), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U754 ( .A(KEYINPUT74), .B(G132), .Z(G219) );
  NOR2_X1 U755 ( .A1(G219), .A2(G220), .ZN(n672) );
  XOR2_X1 U756 ( .A(KEYINPUT84), .B(n672), .Z(n673) );
  XNOR2_X1 U757 ( .A(n673), .B(KEYINPUT22), .ZN(n674) );
  NOR2_X1 U758 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U759 ( .A1(G96), .A2(n675), .ZN(n838) );
  NAND2_X1 U760 ( .A1(G2106), .A2(n838), .ZN(n679) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n676) );
  NOR2_X1 U762 ( .A1(G237), .A2(n676), .ZN(n677) );
  NAND2_X1 U763 ( .A1(G108), .A2(n677), .ZN(n837) );
  NAND2_X1 U764 ( .A1(G567), .A2(n837), .ZN(n678) );
  NAND2_X1 U765 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U766 ( .A(KEYINPUT85), .B(n680), .ZN(G319) );
  INV_X1 U767 ( .A(G319), .ZN(n682) );
  NAND2_X1 U768 ( .A1(G661), .A2(G483), .ZN(n681) );
  NOR2_X1 U769 ( .A1(n682), .A2(n681), .ZN(n834) );
  NAND2_X1 U770 ( .A1(n834), .A2(G36), .ZN(G176) );
  INV_X1 U771 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U772 ( .A(KEYINPUT91), .B(n797), .ZN(n685) );
  XNOR2_X1 U773 ( .A(n684), .B(KEYINPUT64), .ZN(n798) );
  NAND2_X1 U774 ( .A1(n685), .A2(n798), .ZN(n695) );
  INV_X1 U775 ( .A(G1996), .ZN(n1009) );
  NOR2_X2 U776 ( .A1(n695), .A2(n1009), .ZN(n686) );
  XNOR2_X1 U777 ( .A(n686), .B(KEYINPUT26), .ZN(n690) );
  NAND2_X1 U778 ( .A1(n695), .A2(G1341), .ZN(n688) );
  INV_X1 U779 ( .A(n959), .ZN(n687) );
  NAND2_X1 U780 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U781 ( .A1(n690), .A2(n689), .ZN(n692) );
  INV_X1 U782 ( .A(KEYINPUT65), .ZN(n691) );
  XNOR2_X1 U783 ( .A(n692), .B(n691), .ZN(n694) );
  NOR2_X2 U784 ( .A1(n694), .A2(n958), .ZN(n693) );
  XNOR2_X1 U785 ( .A(n693), .B(KEYINPUT93), .ZN(n701) );
  NAND2_X1 U786 ( .A1(n694), .A2(n958), .ZN(n699) );
  INV_X1 U787 ( .A(n695), .ZN(n716) );
  NOR2_X1 U788 ( .A1(n716), .A2(G1348), .ZN(n697) );
  NOR2_X1 U789 ( .A1(G2067), .A2(n736), .ZN(n696) );
  NOR2_X1 U790 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U792 ( .A1(n701), .A2(n700), .ZN(n708) );
  NAND2_X1 U793 ( .A1(n716), .A2(G2072), .ZN(n703) );
  NAND2_X1 U794 ( .A1(G1956), .A2(n736), .ZN(n704) );
  NAND2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n711) );
  NOR2_X1 U796 ( .A1(G299), .A2(n711), .ZN(n706) );
  XOR2_X1 U797 ( .A(KEYINPUT94), .B(n706), .Z(n707) );
  NAND2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n710) );
  XNOR2_X1 U799 ( .A(n710), .B(n709), .ZN(n714) );
  NAND2_X1 U800 ( .A1(G299), .A2(n711), .ZN(n712) );
  XNOR2_X1 U801 ( .A(KEYINPUT28), .B(n712), .ZN(n713) );
  NAND2_X1 U802 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U803 ( .A(n715), .B(KEYINPUT29), .ZN(n720) );
  NOR2_X1 U804 ( .A1(n716), .A2(G1961), .ZN(n718) );
  XOR2_X1 U805 ( .A(G2078), .B(KEYINPUT25), .Z(n1015) );
  NOR2_X1 U806 ( .A1(n736), .A2(n1015), .ZN(n717) );
  NOR2_X1 U807 ( .A1(n718), .A2(n717), .ZN(n725) );
  NOR2_X1 U808 ( .A1(G301), .A2(n725), .ZN(n719) );
  NOR2_X2 U809 ( .A1(n720), .A2(n719), .ZN(n746) );
  NAND2_X1 U810 ( .A1(G8), .A2(n736), .ZN(n778) );
  NOR2_X1 U811 ( .A1(G2084), .A2(n736), .ZN(n732) );
  NOR2_X1 U812 ( .A1(n729), .A2(n732), .ZN(n721) );
  NAND2_X1 U813 ( .A1(G8), .A2(n721), .ZN(n723) );
  NOR2_X1 U814 ( .A1(G168), .A2(n724), .ZN(n727) );
  AND2_X1 U815 ( .A1(G301), .A2(n725), .ZN(n726) );
  NOR2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U817 ( .A(n728), .B(KEYINPUT31), .ZN(n744) );
  NOR2_X1 U818 ( .A1(n746), .A2(n744), .ZN(n730) );
  NOR2_X1 U819 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U820 ( .A(n731), .B(KEYINPUT97), .ZN(n735) );
  NAND2_X1 U821 ( .A1(G8), .A2(n732), .ZN(n733) );
  XOR2_X1 U822 ( .A(KEYINPUT92), .B(n733), .Z(n734) );
  NOR2_X1 U823 ( .A1(n735), .A2(n734), .ZN(n754) );
  INV_X1 U824 ( .A(G8), .ZN(n742) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n736), .ZN(n737) );
  XNOR2_X1 U826 ( .A(n737), .B(KEYINPUT98), .ZN(n739) );
  NOR2_X1 U827 ( .A1(n778), .A2(G1971), .ZN(n738) );
  NOR2_X1 U828 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U829 ( .A1(n740), .A2(G303), .ZN(n741) );
  OR2_X1 U830 ( .A1(n742), .A2(n741), .ZN(n748) );
  INV_X1 U831 ( .A(n748), .ZN(n743) );
  OR2_X1 U832 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n750) );
  NAND2_X1 U834 ( .A1(G286), .A2(G8), .ZN(n747) );
  AND2_X1 U835 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U836 ( .A1(n754), .A2(n753), .ZN(n767) );
  NOR2_X1 U837 ( .A1(G288), .A2(G1976), .ZN(n755) );
  XOR2_X1 U838 ( .A(n755), .B(KEYINPUT99), .Z(n759) );
  NOR2_X1 U839 ( .A1(G1971), .A2(G303), .ZN(n756) );
  NOR2_X1 U840 ( .A1(n759), .A2(n756), .ZN(n955) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n954) );
  NAND2_X1 U842 ( .A1(n757), .A2(n954), .ZN(n758) );
  XNOR2_X1 U843 ( .A(n758), .B(KEYINPUT101), .ZN(n762) );
  XOR2_X1 U844 ( .A(G1981), .B(G305), .Z(n968) );
  INV_X1 U845 ( .A(n778), .ZN(n771) );
  AND2_X1 U846 ( .A1(n771), .A2(n759), .ZN(n760) );
  NAND2_X1 U847 ( .A1(KEYINPUT33), .A2(n760), .ZN(n761) );
  NAND2_X1 U848 ( .A1(n968), .A2(n761), .ZN(n763) );
  NAND2_X1 U849 ( .A1(n762), .A2(n517), .ZN(n765) );
  INV_X1 U850 ( .A(n763), .ZN(n764) );
  NAND2_X1 U851 ( .A1(n765), .A2(n518), .ZN(n766) );
  XNOR2_X1 U852 ( .A(n766), .B(KEYINPUT102), .ZN(n774) );
  NAND2_X1 U853 ( .A1(G8), .A2(G166), .ZN(n768) );
  NOR2_X1 U854 ( .A1(G2090), .A2(n768), .ZN(n769) );
  NOR2_X1 U855 ( .A1(n767), .A2(n769), .ZN(n770) );
  NOR2_X1 U856 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U857 ( .A(KEYINPUT103), .B(n772), .Z(n773) );
  XNOR2_X1 U858 ( .A(n775), .B(KEYINPUT104), .ZN(n821) );
  NOR2_X1 U859 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U860 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  NOR2_X1 U861 ( .A1(n778), .A2(n777), .ZN(n819) );
  NAND2_X1 U862 ( .A1(G129), .A2(n888), .ZN(n780) );
  NAND2_X1 U863 ( .A1(G141), .A2(n616), .ZN(n779) );
  NAND2_X1 U864 ( .A1(n780), .A2(n779), .ZN(n785) );
  XOR2_X1 U865 ( .A(KEYINPUT38), .B(KEYINPUT89), .Z(n782) );
  NAND2_X1 U866 ( .A1(G105), .A2(n534), .ZN(n781) );
  XNOR2_X1 U867 ( .A(n782), .B(n781), .ZN(n783) );
  XOR2_X1 U868 ( .A(KEYINPUT88), .B(n783), .Z(n784) );
  NOR2_X1 U869 ( .A1(n785), .A2(n784), .ZN(n787) );
  NAND2_X1 U870 ( .A1(n886), .A2(G117), .ZN(n786) );
  NAND2_X1 U871 ( .A1(n787), .A2(n786), .ZN(n868) );
  NOR2_X1 U872 ( .A1(G1996), .A2(n868), .ZN(n938) );
  NAND2_X1 U873 ( .A1(G119), .A2(n888), .ZN(n789) );
  NAND2_X1 U874 ( .A1(G107), .A2(n886), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U876 ( .A(KEYINPUT87), .B(n790), .ZN(n794) );
  NAND2_X1 U877 ( .A1(n534), .A2(G95), .ZN(n792) );
  NAND2_X1 U878 ( .A1(G131), .A2(n616), .ZN(n791) );
  AND2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U880 ( .A1(n794), .A2(n793), .ZN(n869) );
  NAND2_X1 U881 ( .A1(G1991), .A2(n869), .ZN(n796) );
  NAND2_X1 U882 ( .A1(G1996), .A2(n868), .ZN(n795) );
  NAND2_X1 U883 ( .A1(n796), .A2(n795), .ZN(n931) );
  NOR2_X1 U884 ( .A1(n797), .A2(n798), .ZN(n822) );
  NAND2_X1 U885 ( .A1(n931), .A2(n822), .ZN(n799) );
  XOR2_X1 U886 ( .A(KEYINPUT90), .B(n799), .Z(n823) );
  NOR2_X1 U887 ( .A1(G1991), .A2(n869), .ZN(n929) );
  NOR2_X1 U888 ( .A1(G1986), .A2(G290), .ZN(n800) );
  NOR2_X1 U889 ( .A1(n929), .A2(n800), .ZN(n801) );
  NOR2_X1 U890 ( .A1(n823), .A2(n801), .ZN(n802) );
  NOR2_X1 U891 ( .A1(n938), .A2(n802), .ZN(n803) );
  XNOR2_X1 U892 ( .A(n803), .B(KEYINPUT39), .ZN(n814) );
  XNOR2_X1 U893 ( .A(G2067), .B(KEYINPUT37), .ZN(n815) );
  NAND2_X1 U894 ( .A1(G104), .A2(n534), .ZN(n805) );
  NAND2_X1 U895 ( .A1(G140), .A2(n616), .ZN(n804) );
  NAND2_X1 U896 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U897 ( .A(KEYINPUT34), .B(n806), .ZN(n811) );
  NAND2_X1 U898 ( .A1(G128), .A2(n888), .ZN(n808) );
  NAND2_X1 U899 ( .A1(G116), .A2(n886), .ZN(n807) );
  NAND2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U901 ( .A(KEYINPUT35), .B(n809), .Z(n810) );
  NOR2_X1 U902 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U903 ( .A(KEYINPUT36), .B(n812), .ZN(n899) );
  NOR2_X1 U904 ( .A1(n815), .A2(n899), .ZN(n935) );
  NAND2_X1 U905 ( .A1(n935), .A2(n822), .ZN(n813) );
  XNOR2_X1 U906 ( .A(n813), .B(KEYINPUT86), .ZN(n825) );
  NAND2_X1 U907 ( .A1(n814), .A2(n825), .ZN(n816) );
  NAND2_X1 U908 ( .A1(n815), .A2(n899), .ZN(n946) );
  NAND2_X1 U909 ( .A1(n816), .A2(n946), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n817), .A2(n822), .ZN(n829) );
  INV_X1 U911 ( .A(n829), .ZN(n818) );
  NOR2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U913 ( .A1(n821), .A2(n820), .ZN(n830) );
  XNOR2_X1 U914 ( .A(G1986), .B(G290), .ZN(n961) );
  AND2_X1 U915 ( .A1(n961), .A2(n822), .ZN(n827) );
  INV_X1 U916 ( .A(n823), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n825), .A2(n824), .ZN(n826) );
  OR2_X1 U918 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U919 ( .A(n831), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U922 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G1), .A2(G3), .ZN(n835) );
  NAND2_X1 U924 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U925 ( .A(n836), .B(KEYINPUT106), .ZN(G188) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G69), .ZN(G235) );
  NOR2_X1 U929 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U930 ( .A(n839), .B(KEYINPUT107), .ZN(G261) );
  INV_X1 U931 ( .A(G261), .ZN(G325) );
  XOR2_X1 U932 ( .A(G2096), .B(KEYINPUT43), .Z(n841) );
  XNOR2_X1 U933 ( .A(G2072), .B(KEYINPUT108), .ZN(n840) );
  XNOR2_X1 U934 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U935 ( .A(n842), .B(G2678), .Z(n844) );
  XNOR2_X1 U936 ( .A(G2067), .B(G2090), .ZN(n843) );
  XNOR2_X1 U937 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U938 ( .A(KEYINPUT42), .B(G2100), .Z(n846) );
  XNOR2_X1 U939 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U940 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U941 ( .A(n848), .B(n847), .ZN(G227) );
  XOR2_X1 U942 ( .A(G1976), .B(G1971), .Z(n850) );
  XNOR2_X1 U943 ( .A(G1986), .B(G1961), .ZN(n849) );
  XNOR2_X1 U944 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U945 ( .A(G1966), .B(G1981), .Z(n852) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U947 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U948 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U949 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n855) );
  XNOR2_X1 U950 ( .A(n856), .B(n855), .ZN(n858) );
  XOR2_X1 U951 ( .A(G1956), .B(G2474), .Z(n857) );
  XNOR2_X1 U952 ( .A(n858), .B(n857), .ZN(G229) );
  NAND2_X1 U953 ( .A1(G124), .A2(n888), .ZN(n859) );
  XNOR2_X1 U954 ( .A(n859), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U955 ( .A1(G112), .A2(n886), .ZN(n860) );
  XOR2_X1 U956 ( .A(KEYINPUT111), .B(n860), .Z(n861) );
  NAND2_X1 U957 ( .A1(n862), .A2(n861), .ZN(n867) );
  NAND2_X1 U958 ( .A1(G136), .A2(n616), .ZN(n863) );
  XNOR2_X1 U959 ( .A(n863), .B(KEYINPUT110), .ZN(n865) );
  NAND2_X1 U960 ( .A1(n534), .A2(G100), .ZN(n864) );
  NAND2_X1 U961 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U962 ( .A1(n867), .A2(n866), .ZN(G162) );
  XNOR2_X1 U963 ( .A(G160), .B(n868), .ZN(n870) );
  XNOR2_X1 U964 ( .A(n870), .B(n869), .ZN(n898) );
  NAND2_X1 U965 ( .A1(G106), .A2(n534), .ZN(n872) );
  NAND2_X1 U966 ( .A1(G142), .A2(n616), .ZN(n871) );
  NAND2_X1 U967 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U968 ( .A(n873), .B(KEYINPUT45), .ZN(n875) );
  NAND2_X1 U969 ( .A1(G130), .A2(n888), .ZN(n874) );
  NAND2_X1 U970 ( .A1(n875), .A2(n874), .ZN(n878) );
  NAND2_X1 U971 ( .A1(n886), .A2(G118), .ZN(n876) );
  XOR2_X1 U972 ( .A(KEYINPUT112), .B(n876), .Z(n877) );
  NOR2_X1 U973 ( .A1(n878), .A2(n877), .ZN(n882) );
  XOR2_X1 U974 ( .A(KEYINPUT116), .B(KEYINPUT46), .Z(n880) );
  XNOR2_X1 U975 ( .A(G164), .B(KEYINPUT48), .ZN(n879) );
  XNOR2_X1 U976 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U977 ( .A(n882), .B(n881), .ZN(n896) );
  NAND2_X1 U978 ( .A1(G103), .A2(n534), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G139), .A2(n616), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U981 ( .A(KEYINPUT113), .B(n885), .ZN(n894) );
  NAND2_X1 U982 ( .A1(n886), .A2(G115), .ZN(n887) );
  XNOR2_X1 U983 ( .A(n887), .B(KEYINPUT114), .ZN(n890) );
  NAND2_X1 U984 ( .A1(G127), .A2(n888), .ZN(n889) );
  NAND2_X1 U985 ( .A1(n890), .A2(n889), .ZN(n892) );
  XOR2_X1 U986 ( .A(KEYINPUT115), .B(KEYINPUT47), .Z(n891) );
  XNOR2_X1 U987 ( .A(n892), .B(n891), .ZN(n893) );
  NAND2_X1 U988 ( .A1(n894), .A2(n893), .ZN(n923) );
  XNOR2_X1 U989 ( .A(n923), .B(G162), .ZN(n895) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U991 ( .A(n898), .B(n897), .ZN(n901) );
  XNOR2_X1 U992 ( .A(n899), .B(n928), .ZN(n900) );
  XNOR2_X1 U993 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U994 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U995 ( .A(n958), .B(G286), .Z(n903) );
  XNOR2_X1 U996 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U997 ( .A(n905), .B(G171), .ZN(n906) );
  NOR2_X1 U998 ( .A1(G37), .A2(n906), .ZN(G397) );
  XOR2_X1 U999 ( .A(KEYINPUT105), .B(G2427), .Z(n908) );
  XNOR2_X1 U1000 ( .A(G2435), .B(G2438), .ZN(n907) );
  XNOR2_X1 U1001 ( .A(n908), .B(n907), .ZN(n915) );
  XOR2_X1 U1002 ( .A(G2443), .B(G2430), .Z(n910) );
  XNOR2_X1 U1003 ( .A(G2454), .B(G2446), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1005 ( .A(n911), .B(G2451), .Z(n913) );
  XNOR2_X1 U1006 ( .A(G1348), .B(G1341), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1008 ( .A(n915), .B(n914), .ZN(n916) );
  NAND2_X1 U1009 ( .A1(n916), .A2(G14), .ZN(n922) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n922), .ZN(n919) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1015 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G96), .ZN(G221) );
  INV_X1 U1018 ( .A(G108), .ZN(G238) );
  INV_X1 U1019 ( .A(n922), .ZN(G401) );
  XNOR2_X1 U1020 ( .A(G164), .B(G2078), .ZN(n926) );
  XNOR2_X1 U1021 ( .A(G2072), .B(KEYINPUT119), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(n924), .B(n923), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(n927), .B(KEYINPUT50), .ZN(n944) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n933) );
  XOR2_X1 U1026 ( .A(G160), .B(G2084), .Z(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1030 ( .A(KEYINPUT117), .B(n936), .ZN(n941) );
  XOR2_X1 U1031 ( .A(G2090), .B(G162), .Z(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(KEYINPUT51), .B(n939), .ZN(n940) );
  NOR2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1035 ( .A(KEYINPUT118), .B(n942), .Z(n943) );
  NOR2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1037 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1038 ( .A(n947), .B(KEYINPUT52), .ZN(n948) );
  XNOR2_X1 U1039 ( .A(n948), .B(KEYINPUT120), .ZN(n949) );
  NOR2_X1 U1040 ( .A1(KEYINPUT55), .A2(n949), .ZN(n950) );
  XNOR2_X1 U1041 ( .A(KEYINPUT121), .B(n950), .ZN(n951) );
  NAND2_X1 U1042 ( .A1(n951), .A2(G29), .ZN(n1004) );
  XNOR2_X1 U1043 ( .A(G1961), .B(G171), .ZN(n953) );
  NAND2_X1 U1044 ( .A1(G1971), .A2(G303), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n957) );
  NAND2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1047 ( .A1(n957), .A2(n956), .ZN(n967) );
  XNOR2_X1 U1048 ( .A(G1348), .B(n958), .ZN(n963) );
  XNOR2_X1 U1049 ( .A(G1341), .B(n959), .ZN(n960) );
  NOR2_X1 U1050 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1051 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1052 ( .A(G1956), .B(G299), .ZN(n964) );
  NOR2_X1 U1053 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1054 ( .A1(n967), .A2(n966), .ZN(n972) );
  XNOR2_X1 U1055 ( .A(G1966), .B(G168), .ZN(n969) );
  NAND2_X1 U1056 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1057 ( .A(KEYINPUT57), .B(n970), .Z(n971) );
  NOR2_X1 U1058 ( .A1(n972), .A2(n971), .ZN(n974) );
  XOR2_X1 U1059 ( .A(KEYINPUT56), .B(G16), .Z(n973) );
  NOR2_X1 U1060 ( .A1(n974), .A2(n973), .ZN(n1002) );
  XNOR2_X1 U1061 ( .A(KEYINPUT125), .B(G1961), .ZN(n975) );
  XNOR2_X1 U1062 ( .A(n975), .B(G5), .ZN(n985) );
  XOR2_X1 U1063 ( .A(G1966), .B(KEYINPUT127), .Z(n976) );
  XNOR2_X1 U1064 ( .A(G21), .B(n976), .ZN(n983) );
  XNOR2_X1 U1065 ( .A(G1971), .B(G22), .ZN(n978) );
  XNOR2_X1 U1066 ( .A(G23), .B(G1976), .ZN(n977) );
  NOR2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n980) );
  XOR2_X1 U1068 ( .A(G1986), .B(G24), .Z(n979) );
  NAND2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(KEYINPUT58), .B(n981), .ZN(n982) );
  NOR2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1072 ( .A1(n985), .A2(n984), .ZN(n996) );
  XOR2_X1 U1073 ( .A(G1341), .B(G19), .Z(n989) );
  XNOR2_X1 U1074 ( .A(G1981), .B(G6), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(G20), .B(G1956), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(KEYINPUT126), .B(n990), .ZN(n993) );
  XOR2_X1 U1079 ( .A(KEYINPUT59), .B(G1348), .Z(n991) );
  XNOR2_X1 U1080 ( .A(G4), .B(n991), .ZN(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1082 ( .A(KEYINPUT60), .B(n994), .Z(n995) );
  NOR2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(KEYINPUT61), .B(n997), .ZN(n999) );
  INV_X1 U1085 ( .A(G16), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(G11), .ZN(n1001) );
  NOR2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1089 ( .A1(n1004), .A2(n1003), .ZN(n1028) );
  XNOR2_X1 U1090 ( .A(G2084), .B(G34), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(n1005), .B(KEYINPUT54), .ZN(n1023) );
  XNOR2_X1 U1092 ( .A(G2090), .B(G35), .ZN(n1020) );
  XNOR2_X1 U1093 ( .A(G1991), .B(G25), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G33), .B(G2072), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1014) );
  XOR2_X1 U1096 ( .A(G2067), .B(G26), .Z(n1008) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(G28), .ZN(n1012) );
  XOR2_X1 U1098 ( .A(KEYINPUT122), .B(n1009), .Z(n1010) );
  XNOR2_X1 U1099 ( .A(G32), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(G27), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT53), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(n1021), .B(KEYINPUT123), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1108 ( .A(KEYINPUT55), .B(n1024), .Z(n1025) );
  XNOR2_X1 U1109 ( .A(KEYINPUT124), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1110 ( .A1(G29), .A2(n1026), .ZN(n1027) );
  NOR2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1112 ( .A(n1029), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

