

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n369, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819;

  INV_X1 U392 ( .A(n622), .ZN(n374) );
  XNOR2_X1 U393 ( .A(G143), .B(G131), .ZN(n467) );
  XNOR2_X1 U394 ( .A(G107), .B(G110), .ZN(n538) );
  XNOR2_X1 U395 ( .A(G116), .B(G107), .ZN(n480) );
  XNOR2_X1 U396 ( .A(KEYINPUT78), .B(KEYINPUT4), .ZN(n485) );
  XNOR2_X1 U397 ( .A(KEYINPUT16), .B(G110), .ZN(n479) );
  INV_X1 U398 ( .A(G104), .ZN(n463) );
  XNOR2_X2 U399 ( .A(n369), .B(KEYINPUT32), .ZN(n739) );
  NAND2_X1 U400 ( .A1(n431), .A2(n627), .ZN(n369) );
  NAND2_X4 U401 ( .A1(n675), .A2(n409), .ZN(n736) );
  NAND2_X4 U402 ( .A1(n488), .A2(G214), .ZN(n748) );
  XOR2_X2 U403 ( .A(KEYINPUT62), .B(n705), .Z(n706) );
  XNOR2_X2 U404 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X2 U405 ( .A(n723), .B(KEYINPUT59), .ZN(n724) );
  XOR2_X2 U406 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n658) );
  XNOR2_X2 U407 ( .A(n809), .B(n399), .ZN(n669) );
  AND2_X2 U408 ( .A1(n382), .A2(n387), .ZN(n386) );
  XNOR2_X1 U409 ( .A(n590), .B(n447), .ZN(n446) );
  XNOR2_X1 U410 ( .A(G101), .B(G104), .ZN(n537) );
  INV_X1 U411 ( .A(G237), .ZN(n487) );
  INV_X1 U412 ( .A(G902), .ZN(n500) );
  INV_X1 U413 ( .A(n759), .ZN(n649) );
  BUF_X1 U414 ( .A(G113), .Z(n694) );
  XNOR2_X2 U415 ( .A(n570), .B(KEYINPUT41), .ZN(n781) );
  NOR2_X2 U416 ( .A1(n753), .A2(n750), .ZN(n570) );
  NAND2_X2 U417 ( .A1(n440), .A2(n667), .ZN(n668) );
  NOR2_X1 U418 ( .A1(n649), .A2(n764), .ZN(n621) );
  NAND2_X1 U419 ( .A1(n391), .A2(n439), .ZN(n385) );
  NAND2_X1 U420 ( .A1(n383), .A2(n384), .ZN(n391) );
  AND2_X1 U421 ( .A1(n558), .A2(n375), .ZN(n377) );
  INV_X1 U422 ( .A(n645), .ZN(n754) );
  INV_X1 U423 ( .A(n595), .ZN(n375) );
  NOR2_X1 U424 ( .A1(n557), .A2(n376), .ZN(n379) );
  AND2_X1 U425 ( .A1(n419), .A2(n390), .ZN(n439) );
  XNOR2_X1 U426 ( .A(n484), .B(n456), .ZN(n492) );
  INV_X1 U427 ( .A(KEYINPUT31), .ZN(n394) );
  INV_X1 U428 ( .A(KEYINPUT80), .ZN(n432) );
  INV_X1 U429 ( .A(KEYINPUT66), .ZN(n390) );
  NAND2_X1 U430 ( .A1(n386), .A2(n385), .ZN(n440) );
  AND2_X1 U431 ( .A1(n388), .A2(n437), .ZN(n387) );
  NOR2_X1 U432 ( .A1(n554), .A2(n553), .ZN(n566) );
  XNOR2_X1 U433 ( .A(n395), .B(n394), .ZN(n692) );
  AND2_X1 U434 ( .A1(n417), .A2(n414), .ZN(n403) );
  XNOR2_X1 U435 ( .A(n536), .B(n381), .ZN(n380) );
  AND2_X1 U436 ( .A1(n417), .A2(KEYINPUT67), .ZN(n405) );
  XNOR2_X1 U437 ( .A(n626), .B(n432), .ZN(n627) );
  NOR2_X1 U438 ( .A1(n575), .A2(n574), .ZN(n576) );
  OR2_X1 U439 ( .A1(n621), .A2(KEYINPUT67), .ZN(n427) );
  BUF_X2 U440 ( .A(n555), .Z(n764) );
  XNOR2_X1 U441 ( .A(n504), .B(n503), .ZN(n555) );
  OR2_X1 U442 ( .A1(n712), .A2(G902), .ZN(n436) );
  XNOR2_X1 U443 ( .A(n545), .B(n424), .ZN(n501) );
  XNOR2_X1 U444 ( .A(n545), .B(n544), .ZN(n712) );
  XNOR2_X1 U445 ( .A(n426), .B(n425), .ZN(n424) );
  INV_X1 U446 ( .A(n762), .ZN(n376) );
  XNOR2_X1 U447 ( .A(n495), .B(n499), .ZN(n426) );
  XNOR2_X1 U448 ( .A(n696), .B(G146), .ZN(n545) );
  XNOR2_X1 U449 ( .A(n492), .B(n491), .ZN(n696) );
  XNOR2_X1 U450 ( .A(n615), .B(KEYINPUT69), .ZN(n616) );
  INV_X1 U451 ( .A(n535), .ZN(n381) );
  XNOR2_X2 U452 ( .A(G122), .B(KEYINPUT9), .ZN(n454) );
  XNOR2_X2 U453 ( .A(G902), .B(KEYINPUT15), .ZN(n660) );
  NOR2_X2 U454 ( .A1(G953), .A2(G237), .ZN(n496) );
  XNOR2_X1 U455 ( .A(n430), .B(n619), .ZN(n431) );
  NOR2_X1 U456 ( .A1(n818), .A2(n819), .ZN(n580) );
  XNOR2_X1 U457 ( .A(n577), .B(n578), .ZN(n818) );
  NAND2_X1 U458 ( .A1(n378), .A2(n377), .ZN(n575) );
  INV_X1 U459 ( .A(n559), .ZN(n378) );
  NAND2_X1 U460 ( .A1(n374), .A2(n379), .ZN(n588) );
  NAND2_X1 U461 ( .A1(n380), .A2(n375), .ZN(n571) );
  NAND2_X1 U462 ( .A1(n407), .A2(n389), .ZN(n382) );
  INV_X1 U463 ( .A(n444), .ZN(n383) );
  INV_X1 U464 ( .A(n441), .ZN(n384) );
  NAND2_X1 U465 ( .A1(n695), .A2(n439), .ZN(n388) );
  NOR2_X1 U466 ( .A1(n695), .A2(n390), .ZN(n389) );
  XNOR2_X2 U467 ( .A(n659), .B(n658), .ZN(n664) );
  AND2_X1 U468 ( .A1(n404), .A2(n402), .ZN(n730) );
  XNOR2_X1 U469 ( .A(n620), .B(n619), .ZN(n421) );
  XNOR2_X1 U470 ( .A(n400), .B(n486), .ZN(n399) );
  XNOR2_X1 U471 ( .A(n392), .B(n482), .ZN(n398) );
  XNOR2_X1 U472 ( .A(n392), .B(KEYINPUT10), .ZN(n519) );
  XNOR2_X2 U473 ( .A(G146), .B(G125), .ZN(n392) );
  XNOR2_X2 U474 ( .A(n393), .B(n493), .ZN(n401) );
  XNOR2_X2 U475 ( .A(n464), .B(n463), .ZN(n393) );
  XNOR2_X1 U476 ( .A(n393), .B(n519), .ZN(n471) );
  NAND2_X1 U477 ( .A1(n692), .A2(n686), .ZN(n646) );
  NAND2_X1 U478 ( .A1(n644), .A2(n396), .ZN(n395) );
  INV_X1 U479 ( .A(n770), .ZN(n396) );
  XNOR2_X2 U480 ( .A(n397), .B(n489), .ZN(n590) );
  NAND2_X2 U481 ( .A1(n562), .A2(n748), .ZN(n397) );
  XNOR2_X2 U482 ( .A(n410), .B(n411), .ZN(n562) );
  XNOR2_X1 U483 ( .A(n398), .B(n483), .ZN(n400) );
  XNOR2_X2 U484 ( .A(n401), .B(n481), .ZN(n809) );
  XNOR2_X2 U485 ( .A(n478), .B(n477), .ZN(n493) );
  NAND2_X1 U486 ( .A1(n421), .A2(n403), .ZN(n402) );
  NAND2_X1 U487 ( .A1(n420), .A2(n405), .ZN(n404) );
  NAND2_X1 U488 ( .A1(n739), .A2(n730), .ZN(n638) );
  XNOR2_X1 U489 ( .A(n498), .B(n494), .ZN(n425) );
  NOR2_X1 U490 ( .A1(n441), .A2(n444), .ZN(n407) );
  BUF_X1 U491 ( .A(n729), .Z(n408) );
  XNOR2_X1 U492 ( .A(n433), .B(KEYINPUT35), .ZN(n729) );
  INV_X2 U493 ( .A(n811), .ZN(n409) );
  INV_X4 U494 ( .A(G953), .ZN(n811) );
  NOR2_X2 U495 ( .A1(n669), .A2(n662), .ZN(n410) );
  NAND2_X1 U496 ( .A1(n488), .A2(G210), .ZN(n411) );
  BUF_X1 U497 ( .A(n739), .Z(n412) );
  INV_X1 U498 ( .A(KEYINPUT6), .ZN(n423) );
  NAND2_X1 U499 ( .A1(n660), .A2(n661), .ZN(n442) );
  NAND2_X1 U500 ( .A1(n438), .A2(KEYINPUT66), .ZN(n437) );
  XOR2_X1 U501 ( .A(G116), .B(KEYINPUT98), .Z(n494) );
  INV_X1 U502 ( .A(G134), .ZN(n456) );
  OR2_X2 U503 ( .A1(n589), .A2(n422), .ZN(n603) );
  NAND2_X1 U504 ( .A1(n501), .A2(n500), .ZN(n504) );
  XNOR2_X1 U505 ( .A(G140), .B(KEYINPUT71), .ZN(n518) );
  INV_X1 U506 ( .A(n501), .ZN(n705) );
  NAND2_X1 U507 ( .A1(n650), .A2(n422), .ZN(n651) );
  NOR2_X1 U508 ( .A1(n759), .A2(n758), .ZN(n413) );
  NAND2_X1 U509 ( .A1(n621), .A2(KEYINPUT67), .ZN(n414) );
  AND2_X1 U510 ( .A1(n614), .A2(n613), .ZN(n415) );
  NOR2_X1 U511 ( .A1(n757), .A2(n435), .ZN(n416) );
  AND2_X1 U512 ( .A1(n427), .A2(n374), .ZN(n417) );
  XOR2_X1 U513 ( .A(n630), .B(KEYINPUT34), .Z(n418) );
  NAND2_X1 U514 ( .A1(n662), .A2(KEYINPUT2), .ZN(n419) );
  INV_X1 U515 ( .A(n421), .ZN(n420) );
  NAND2_X1 U516 ( .A1(n413), .A2(n623), .ZN(n628) );
  INV_X1 U517 ( .A(n623), .ZN(n422) );
  XNOR2_X2 U518 ( .A(n764), .B(n423), .ZN(n623) );
  BUF_X1 U519 ( .A(n446), .Z(n428) );
  XNOR2_X2 U520 ( .A(n668), .B(KEYINPUT65), .ZN(n429) );
  XNOR2_X1 U521 ( .A(n668), .B(KEYINPUT65), .ZN(n732) );
  BUF_X1 U522 ( .A(n493), .Z(n495) );
  NAND2_X1 U523 ( .A1(n629), .A2(n618), .ZN(n430) );
  NAND2_X1 U524 ( .A1(n629), .A2(n618), .ZN(n620) );
  NAND2_X1 U525 ( .A1(n508), .A2(G221), .ZN(n517) );
  XNOR2_X1 U526 ( .A(n452), .B(n451), .ZN(n508) );
  XNOR2_X2 U527 ( .A(KEYINPUT85), .B(KEYINPUT8), .ZN(n450) );
  NAND2_X1 U528 ( .A1(n664), .A2(n661), .ZN(n443) );
  XNOR2_X1 U529 ( .A(n580), .B(n579), .ZN(n581) );
  NAND2_X1 U530 ( .A1(n434), .A2(n633), .ZN(n433) );
  XNOR2_X1 U531 ( .A(n631), .B(n418), .ZN(n434) );
  INV_X1 U532 ( .A(n782), .ZN(n435) );
  XNOR2_X2 U533 ( .A(n628), .B(KEYINPUT33), .ZN(n782) );
  XNOR2_X2 U534 ( .A(n595), .B(KEYINPUT1), .ZN(n759) );
  XNOR2_X2 U535 ( .A(n436), .B(n546), .ZN(n595) );
  INV_X1 U536 ( .A(n419), .ZN(n438) );
  NAND2_X1 U537 ( .A1(n443), .A2(n442), .ZN(n441) );
  NOR2_X1 U538 ( .A1(n664), .A2(n445), .ZN(n444) );
  NAND2_X1 U539 ( .A1(n662), .A2(KEYINPUT87), .ZN(n445) );
  NAND2_X1 U540 ( .A1(n446), .A2(n415), .ZN(n617) );
  NAND2_X1 U541 ( .A1(n448), .A2(n428), .ZN(n547) );
  INV_X1 U542 ( .A(KEYINPUT19), .ZN(n447) );
  INV_X1 U543 ( .A(n571), .ZN(n448) );
  XNOR2_X2 U544 ( .A(G119), .B(G101), .ZN(n478) );
  NAND2_X1 U545 ( .A1(n429), .A2(G210), .ZN(n674) );
  XNOR2_X1 U546 ( .A(KEYINPUT74), .B(KEYINPUT39), .ZN(n449) );
  INV_X1 U547 ( .A(KEYINPUT46), .ZN(n579) );
  INV_X1 U548 ( .A(KEYINPUT87), .ZN(n661) );
  AND2_X1 U549 ( .A1(n598), .A2(n597), .ZN(n599) );
  AND2_X1 U550 ( .A1(n600), .A2(n599), .ZN(n601) );
  INV_X1 U551 ( .A(KEYINPUT22), .ZN(n619) );
  BUF_X1 U552 ( .A(n695), .Z(n741) );
  BUF_X1 U553 ( .A(n732), .Z(n716) );
  BUF_X1 U554 ( .A(n730), .Z(n731) );
  XNOR2_X1 U555 ( .A(n450), .B(KEYINPUT70), .ZN(n452) );
  NAND2_X1 U556 ( .A1(n811), .A2(G234), .ZN(n451) );
  NAND2_X1 U557 ( .A1(n508), .A2(G217), .ZN(n460) );
  XNOR2_X2 U558 ( .A(KEYINPUT100), .B(KEYINPUT7), .ZN(n453) );
  XNOR2_X1 U559 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U560 ( .A(n455), .B(n480), .ZN(n458) );
  XNOR2_X2 U561 ( .A(G128), .B(G143), .ZN(n484) );
  INV_X1 U562 ( .A(n492), .ZN(n457) );
  XNOR2_X1 U563 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U564 ( .A(n460), .B(n459), .ZN(n733) );
  OR2_X1 U565 ( .A1(n733), .A2(G902), .ZN(n462) );
  XNOR2_X1 U566 ( .A(G478), .B(KEYINPUT101), .ZN(n461) );
  XNOR2_X1 U567 ( .A(n462), .B(n461), .ZN(n569) );
  XNOR2_X2 U568 ( .A(G122), .B(G113), .ZN(n464) );
  NAND2_X1 U569 ( .A1(n496), .A2(G214), .ZN(n465) );
  XNOR2_X1 U570 ( .A(n465), .B(KEYINPUT11), .ZN(n469) );
  XNOR2_X1 U571 ( .A(G140), .B(KEYINPUT12), .ZN(n466) );
  XNOR2_X1 U572 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U573 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U574 ( .A(n471), .B(n470), .ZN(n723) );
  OR2_X1 U575 ( .A1(n723), .A2(G902), .ZN(n474) );
  INV_X1 U576 ( .A(KEYINPUT13), .ZN(n472) );
  XNOR2_X1 U577 ( .A(n472), .B(G475), .ZN(n473) );
  XNOR2_X1 U578 ( .A(n474), .B(n473), .ZN(n567) );
  NAND2_X1 U579 ( .A1(n569), .A2(n567), .ZN(n475) );
  XNOR2_X1 U580 ( .A(n475), .B(KEYINPUT102), .ZN(n795) );
  OR2_X1 U581 ( .A1(n569), .A2(n567), .ZN(n790) );
  NAND2_X1 U582 ( .A1(n795), .A2(n790), .ZN(n645) );
  AND2_X1 U583 ( .A1(n754), .A2(KEYINPUT84), .ZN(n476) );
  NOR2_X1 U584 ( .A1(KEYINPUT75), .A2(n476), .ZN(n548) );
  XNOR2_X2 U585 ( .A(KEYINPUT93), .B(KEYINPUT3), .ZN(n477) );
  XNOR2_X1 U586 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U587 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n483) );
  NAND2_X1 U588 ( .A1(n811), .A2(G224), .ZN(n482) );
  XNOR2_X1 U589 ( .A(n484), .B(n485), .ZN(n486) );
  INV_X1 U590 ( .A(n660), .ZN(n662) );
  NAND2_X1 U591 ( .A1(n487), .A2(n500), .ZN(n488) );
  INV_X1 U592 ( .A(KEYINPUT90), .ZN(n489) );
  XNOR2_X2 U593 ( .A(KEYINPUT4), .B(G131), .ZN(n490) );
  XNOR2_X1 U594 ( .A(n490), .B(KEYINPUT72), .ZN(n491) );
  NAND2_X1 U595 ( .A1(n496), .A2(G210), .ZN(n497) );
  XNOR2_X1 U596 ( .A(n497), .B(KEYINPUT5), .ZN(n499) );
  XNOR2_X1 U597 ( .A(G137), .B(n694), .ZN(n498) );
  INV_X1 U598 ( .A(KEYINPUT99), .ZN(n502) );
  XNOR2_X1 U599 ( .A(n502), .B(G472), .ZN(n503) );
  NAND2_X1 U600 ( .A1(n660), .A2(G234), .ZN(n505) );
  XNOR2_X1 U601 ( .A(n505), .B(KEYINPUT20), .ZN(n521) );
  NAND2_X1 U602 ( .A1(n521), .A2(G221), .ZN(n507) );
  INV_X1 U603 ( .A(KEYINPUT21), .ZN(n506) );
  XNOR2_X1 U604 ( .A(n507), .B(n506), .ZN(n762) );
  XOR2_X1 U605 ( .A(KEYINPUT95), .B(G110), .Z(n510) );
  XNOR2_X1 U606 ( .A(G128), .B(G119), .ZN(n509) );
  XNOR2_X1 U607 ( .A(n510), .B(n509), .ZN(n515) );
  XOR2_X1 U608 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n513) );
  XNOR2_X1 U609 ( .A(KEYINPUT94), .B(KEYINPUT96), .ZN(n511) );
  INV_X1 U610 ( .A(n511), .ZN(n512) );
  XNOR2_X1 U611 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U612 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U613 ( .A(n517), .B(n516), .ZN(n520) );
  XNOR2_X1 U614 ( .A(n518), .B(G137), .ZN(n542) );
  XNOR2_X1 U615 ( .A(n519), .B(n542), .ZN(n697) );
  XNOR2_X1 U616 ( .A(n520), .B(n697), .ZN(n717) );
  NAND2_X1 U617 ( .A1(n717), .A2(n500), .ZN(n527) );
  XOR2_X1 U618 ( .A(KEYINPUT97), .B(KEYINPUT76), .Z(n523) );
  NAND2_X1 U619 ( .A1(n521), .A2(G217), .ZN(n522) );
  XNOR2_X1 U620 ( .A(n523), .B(n522), .ZN(n525) );
  INV_X1 U621 ( .A(KEYINPUT25), .ZN(n524) );
  XNOR2_X1 U622 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X2 U623 ( .A(n527), .B(n526), .ZN(n622) );
  NAND2_X1 U624 ( .A1(G237), .A2(G234), .ZN(n528) );
  XNOR2_X1 U625 ( .A(n528), .B(KEYINPUT14), .ZN(n778) );
  NAND2_X1 U626 ( .A1(n811), .A2(G952), .ZN(n530) );
  NAND2_X1 U627 ( .A1(n409), .A2(G902), .ZN(n529) );
  NAND2_X1 U628 ( .A1(n530), .A2(n529), .ZN(n531) );
  AND2_X1 U629 ( .A1(n778), .A2(n531), .ZN(n614) );
  NAND2_X1 U630 ( .A1(n409), .A2(G900), .ZN(n532) );
  NAND2_X1 U631 ( .A1(n614), .A2(n532), .ZN(n533) );
  XOR2_X1 U632 ( .A(KEYINPUT83), .B(n533), .Z(n557) );
  INV_X1 U633 ( .A(n588), .ZN(n534) );
  NAND2_X1 U634 ( .A1(n764), .A2(n534), .ZN(n536) );
  XNOR2_X1 U635 ( .A(KEYINPUT106), .B(KEYINPUT28), .ZN(n535) );
  XNOR2_X1 U636 ( .A(n538), .B(n537), .ZN(n541) );
  NAND2_X1 U637 ( .A1(n811), .A2(G227), .ZN(n539) );
  XNOR2_X1 U638 ( .A(n539), .B(KEYINPUT77), .ZN(n540) );
  XNOR2_X1 U639 ( .A(n541), .B(n540), .ZN(n543) );
  XNOR2_X1 U640 ( .A(n543), .B(n542), .ZN(n544) );
  INV_X1 U641 ( .A(G469), .ZN(n546) );
  XNOR2_X1 U642 ( .A(n547), .B(KEYINPUT82), .ZN(n583) );
  INV_X2 U643 ( .A(n583), .ZN(n797) );
  NAND2_X1 U644 ( .A1(n548), .A2(n797), .ZN(n549) );
  NAND2_X1 U645 ( .A1(n549), .A2(KEYINPUT47), .ZN(n552) );
  AND2_X1 U646 ( .A1(n754), .A2(KEYINPUT75), .ZN(n550) );
  NAND2_X1 U647 ( .A1(n550), .A2(n797), .ZN(n551) );
  NAND2_X1 U648 ( .A1(n552), .A2(n551), .ZN(n554) );
  NOR2_X1 U649 ( .A1(KEYINPUT84), .A2(n754), .ZN(n553) );
  NAND2_X1 U650 ( .A1(n555), .A2(n748), .ZN(n556) );
  XNOR2_X1 U651 ( .A(n556), .B(KEYINPUT30), .ZN(n559) );
  NAND2_X1 U652 ( .A1(n622), .A2(n762), .ZN(n758) );
  NOR2_X1 U653 ( .A1(n758), .A2(n557), .ZN(n558) );
  INV_X1 U654 ( .A(n575), .ZN(n565) );
  INV_X1 U655 ( .A(n569), .ZN(n560) );
  NAND2_X1 U656 ( .A1(n560), .A2(n567), .ZN(n561) );
  XNOR2_X1 U657 ( .A(n561), .B(KEYINPUT104), .ZN(n632) );
  BUF_X1 U658 ( .A(n562), .Z(n563) );
  INV_X1 U659 ( .A(n563), .ZN(n608) );
  NOR2_X1 U660 ( .A1(n632), .A2(n608), .ZN(n564) );
  NAND2_X1 U661 ( .A1(n565), .A2(n564), .ZN(n679) );
  NAND2_X1 U662 ( .A1(n566), .A2(n679), .ZN(n582) );
  XNOR2_X1 U663 ( .A(n563), .B(KEYINPUT38), .ZN(n574) );
  INV_X1 U664 ( .A(n574), .ZN(n749) );
  NAND2_X1 U665 ( .A1(n749), .A2(n748), .ZN(n753) );
  INV_X1 U666 ( .A(n567), .ZN(n568) );
  NAND2_X1 U667 ( .A1(n569), .A2(n568), .ZN(n750) );
  NOR2_X1 U668 ( .A1(n781), .A2(n571), .ZN(n572) );
  XNOR2_X1 U669 ( .A(KEYINPUT42), .B(n572), .ZN(n819) );
  XNOR2_X1 U670 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n573) );
  XOR2_X1 U671 ( .A(n573), .B(KEYINPUT40), .Z(n578) );
  XNOR2_X1 U672 ( .A(n576), .B(n449), .ZN(n610) );
  NOR2_X1 U673 ( .A1(n795), .A2(n610), .ZN(n577) );
  NOR2_X1 U674 ( .A1(n582), .A2(n581), .ZN(n600) );
  NOR2_X1 U675 ( .A1(n583), .A2(KEYINPUT75), .ZN(n584) );
  NAND2_X1 U676 ( .A1(n645), .A2(n584), .ZN(n585) );
  NAND2_X1 U677 ( .A1(n585), .A2(KEYINPUT84), .ZN(n587) );
  INV_X1 U678 ( .A(KEYINPUT47), .ZN(n586) );
  NAND2_X1 U679 ( .A1(n587), .A2(n586), .ZN(n598) );
  OR2_X1 U680 ( .A1(n795), .A2(n588), .ZN(n589) );
  XNOR2_X1 U681 ( .A(n603), .B(KEYINPUT109), .ZN(n592) );
  BUF_X1 U682 ( .A(n590), .Z(n591) );
  NAND2_X1 U683 ( .A1(n592), .A2(n591), .ZN(n594) );
  INV_X1 U684 ( .A(KEYINPUT36), .ZN(n593) );
  XNOR2_X1 U685 ( .A(n594), .B(n593), .ZN(n596) );
  AND2_X1 U686 ( .A1(n596), .A2(n649), .ZN(n800) );
  INV_X1 U687 ( .A(n800), .ZN(n597) );
  XNOR2_X1 U688 ( .A(n601), .B(KEYINPUT48), .ZN(n612) );
  INV_X1 U689 ( .A(n748), .ZN(n602) );
  NOR2_X1 U690 ( .A1(n603), .A2(n602), .ZN(n605) );
  INV_X1 U691 ( .A(KEYINPUT105), .ZN(n604) );
  XNOR2_X1 U692 ( .A(n605), .B(n604), .ZN(n606) );
  NAND2_X1 U693 ( .A1(n606), .A2(n759), .ZN(n607) );
  XNOR2_X1 U694 ( .A(n607), .B(KEYINPUT43), .ZN(n609) );
  NAND2_X1 U695 ( .A1(n609), .A2(n608), .ZN(n689) );
  OR2_X1 U696 ( .A1(n610), .A2(n790), .ZN(n802) );
  AND2_X1 U697 ( .A1(n689), .A2(n802), .ZN(n611) );
  NAND2_X1 U698 ( .A1(n612), .A2(n611), .ZN(n663) );
  XNOR2_X2 U699 ( .A(n663), .B(KEYINPUT88), .ZN(n695) );
  NAND2_X1 U700 ( .A1(n409), .A2(G898), .ZN(n613) );
  XNOR2_X1 U701 ( .A(KEYINPUT92), .B(KEYINPUT0), .ZN(n615) );
  XNOR2_X2 U702 ( .A(n617), .B(n616), .ZN(n629) );
  NOR2_X1 U703 ( .A1(n750), .A2(n376), .ZN(n618) );
  XNOR2_X1 U704 ( .A(n623), .B(KEYINPUT81), .ZN(n625) );
  NOR2_X1 U705 ( .A1(n759), .A2(n622), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U707 ( .A(n638), .B(KEYINPUT89), .ZN(n635) );
  BUF_X2 U708 ( .A(n629), .Z(n644) );
  NAND2_X1 U709 ( .A1(n782), .A2(n644), .ZN(n631) );
  INV_X1 U710 ( .A(KEYINPUT79), .ZN(n630) );
  INV_X1 U711 ( .A(n632), .ZN(n633) );
  NOR2_X1 U712 ( .A1(n729), .A2(KEYINPUT44), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n637) );
  INV_X1 U714 ( .A(KEYINPUT73), .ZN(n636) );
  XNOR2_X1 U715 ( .A(n637), .B(n636), .ZN(n657) );
  OR2_X1 U716 ( .A1(n638), .A2(n729), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n639), .A2(KEYINPUT44), .ZN(n655) );
  INV_X1 U718 ( .A(n758), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n641), .A2(n764), .ZN(n640) );
  OR2_X1 U720 ( .A1(n759), .A2(n640), .ZN(n770) );
  NAND2_X1 U721 ( .A1(n641), .A2(n375), .ZN(n642) );
  NOR2_X1 U722 ( .A1(n642), .A2(n764), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n644), .A2(n643), .ZN(n686) );
  NAND2_X1 U724 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U725 ( .A(n647), .B(KEYINPUT103), .ZN(n653) );
  BUF_X1 U726 ( .A(n431), .Z(n648) );
  INV_X1 U727 ( .A(n648), .ZN(n652) );
  NOR2_X1 U728 ( .A1(n649), .A2(n374), .ZN(n650) );
  NOR2_X1 U729 ( .A1(n652), .A2(n651), .ZN(n690) );
  NOR2_X1 U730 ( .A1(n653), .A2(n690), .ZN(n654) );
  AND2_X1 U731 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n657), .A2(n656), .ZN(n659) );
  BUF_X1 U733 ( .A(n663), .Z(n666) );
  BUF_X1 U734 ( .A(n664), .Z(n665) );
  NOR2_X1 U735 ( .A1(n666), .A2(n665), .ZN(n743) );
  NAND2_X1 U736 ( .A1(n743), .A2(KEYINPUT2), .ZN(n667) );
  BUF_X1 U737 ( .A(n669), .Z(n672) );
  XNOR2_X1 U738 ( .A(KEYINPUT91), .B(KEYINPUT54), .ZN(n670) );
  XOR2_X1 U739 ( .A(n670), .B(KEYINPUT55), .Z(n671) );
  XNOR2_X1 U740 ( .A(n674), .B(n673), .ZN(n676) );
  INV_X1 U741 ( .A(G952), .ZN(n675) );
  NAND2_X1 U742 ( .A1(n676), .A2(n736), .ZN(n678) );
  INV_X1 U743 ( .A(KEYINPUT56), .ZN(n677) );
  XNOR2_X1 U744 ( .A(n678), .B(n677), .ZN(G51) );
  XNOR2_X1 U745 ( .A(n679), .B(G143), .ZN(G45) );
  XOR2_X1 U746 ( .A(G104), .B(KEYINPUT111), .Z(n681) );
  NOR2_X1 U747 ( .A1(n686), .A2(n795), .ZN(n680) );
  XOR2_X1 U748 ( .A(n681), .B(n680), .Z(G6) );
  XOR2_X1 U749 ( .A(KEYINPUT114), .B(KEYINPUT27), .Z(n683) );
  XNOR2_X1 U750 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n682) );
  XNOR2_X1 U751 ( .A(n683), .B(n682), .ZN(n685) );
  XOR2_X1 U752 ( .A(G107), .B(KEYINPUT26), .Z(n684) );
  XNOR2_X1 U753 ( .A(n685), .B(n684), .ZN(n688) );
  NOR2_X1 U754 ( .A1(n686), .A2(n790), .ZN(n687) );
  XOR2_X1 U755 ( .A(n688), .B(n687), .Z(G9) );
  XNOR2_X1 U756 ( .A(n689), .B(G140), .ZN(G42) );
  XOR2_X1 U757 ( .A(G101), .B(n690), .Z(G3) );
  NOR2_X1 U758 ( .A1(n692), .A2(n790), .ZN(n691) );
  XOR2_X1 U759 ( .A(G116), .B(n691), .Z(G18) );
  NOR2_X1 U760 ( .A1(n692), .A2(n795), .ZN(n693) );
  XOR2_X1 U761 ( .A(n694), .B(n693), .Z(G15) );
  XNOR2_X1 U762 ( .A(n696), .B(KEYINPUT127), .ZN(n698) );
  XNOR2_X1 U763 ( .A(n698), .B(n697), .ZN(n700) );
  XNOR2_X1 U764 ( .A(n741), .B(n700), .ZN(n699) );
  NAND2_X1 U765 ( .A1(n699), .A2(n811), .ZN(n704) );
  XNOR2_X1 U766 ( .A(n700), .B(G227), .ZN(n701) );
  NAND2_X1 U767 ( .A1(n701), .A2(G900), .ZN(n702) );
  NAND2_X1 U768 ( .A1(n409), .A2(n702), .ZN(n703) );
  NAND2_X1 U769 ( .A1(n704), .A2(n703), .ZN(G72) );
  NAND2_X1 U770 ( .A1(n429), .A2(G472), .ZN(n707) );
  XNOR2_X1 U771 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U772 ( .A1(n708), .A2(n736), .ZN(n710) );
  XNOR2_X1 U773 ( .A(KEYINPUT110), .B(KEYINPUT63), .ZN(n709) );
  XNOR2_X1 U774 ( .A(n710), .B(n709), .ZN(G57) );
  NAND2_X1 U775 ( .A1(n716), .A2(G469), .ZN(n714) );
  XOR2_X1 U776 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n711) );
  XNOR2_X1 U777 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U778 ( .A(n714), .B(n713), .ZN(n715) );
  INV_X1 U779 ( .A(n736), .ZN(n721) );
  NOR2_X1 U780 ( .A1(n715), .A2(n721), .ZN(G54) );
  NAND2_X1 U781 ( .A1(n716), .A2(G217), .ZN(n720) );
  BUF_X1 U782 ( .A(n717), .Z(n718) );
  XOR2_X1 U783 ( .A(KEYINPUT122), .B(n718), .Z(n719) );
  XNOR2_X1 U784 ( .A(n720), .B(n719), .ZN(n722) );
  NOR2_X1 U785 ( .A1(n722), .A2(n721), .ZN(G66) );
  NAND2_X1 U786 ( .A1(n429), .A2(G475), .ZN(n725) );
  XNOR2_X1 U787 ( .A(n725), .B(n724), .ZN(n726) );
  NAND2_X1 U788 ( .A1(n726), .A2(n736), .ZN(n728) );
  XOR2_X1 U789 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n727) );
  XNOR2_X1 U790 ( .A(n728), .B(n727), .ZN(G60) );
  XOR2_X1 U791 ( .A(G122), .B(n408), .Z(G24) );
  XNOR2_X1 U792 ( .A(n731), .B(G110), .ZN(G12) );
  NAND2_X1 U793 ( .A1(n732), .A2(G478), .ZN(n735) );
  INV_X1 U794 ( .A(n733), .ZN(n734) );
  XNOR2_X1 U795 ( .A(n735), .B(n734), .ZN(n737) );
  NAND2_X1 U796 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U797 ( .A(n738), .B(KEYINPUT121), .ZN(G63) );
  XNOR2_X1 U798 ( .A(n412), .B(G119), .ZN(G21) );
  XNOR2_X1 U799 ( .A(n665), .B(KEYINPUT86), .ZN(n740) );
  NOR2_X1 U800 ( .A1(n741), .A2(n740), .ZN(n742) );
  OR2_X1 U801 ( .A1(n742), .A2(KEYINPUT2), .ZN(n747) );
  INV_X1 U802 ( .A(n743), .ZN(n744) );
  NAND2_X1 U803 ( .A1(n744), .A2(KEYINPUT86), .ZN(n745) );
  NAND2_X1 U804 ( .A1(n745), .A2(KEYINPUT2), .ZN(n746) );
  NAND2_X1 U805 ( .A1(n747), .A2(n746), .ZN(n788) );
  NOR2_X1 U806 ( .A1(n749), .A2(n748), .ZN(n751) );
  NOR2_X1 U807 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U808 ( .A(KEYINPUT119), .B(n752), .Z(n756) );
  NOR2_X1 U809 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U810 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U811 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U812 ( .A(KEYINPUT50), .B(n760), .Z(n768) );
  NOR2_X1 U813 ( .A1(n762), .A2(n622), .ZN(n763) );
  XNOR2_X1 U814 ( .A(n763), .B(KEYINPUT49), .ZN(n766) );
  INV_X1 U815 ( .A(n764), .ZN(n765) );
  NAND2_X1 U816 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U817 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U818 ( .A(n769), .B(KEYINPUT117), .ZN(n771) );
  NAND2_X1 U819 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U820 ( .A(KEYINPUT51), .B(n772), .ZN(n773) );
  NOR2_X1 U821 ( .A1(n781), .A2(n773), .ZN(n774) );
  XNOR2_X1 U822 ( .A(n774), .B(KEYINPUT118), .ZN(n775) );
  NOR2_X1 U823 ( .A1(n416), .A2(n775), .ZN(n776) );
  XNOR2_X1 U824 ( .A(KEYINPUT120), .B(n776), .ZN(n777) );
  XNOR2_X1 U825 ( .A(KEYINPUT52), .B(n777), .ZN(n780) );
  NAND2_X1 U826 ( .A1(G952), .A2(n778), .ZN(n779) );
  NOR2_X1 U827 ( .A1(n780), .A2(n779), .ZN(n786) );
  INV_X1 U828 ( .A(n781), .ZN(n783) );
  NAND2_X1 U829 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U830 ( .A1(n784), .A2(n811), .ZN(n785) );
  NOR2_X1 U831 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U832 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U833 ( .A(KEYINPUT53), .B(n789), .Z(G75) );
  XOR2_X1 U834 ( .A(KEYINPUT29), .B(KEYINPUT115), .Z(n793) );
  INV_X1 U835 ( .A(n790), .ZN(n791) );
  NAND2_X1 U836 ( .A1(n797), .A2(n791), .ZN(n792) );
  XNOR2_X1 U837 ( .A(n793), .B(n792), .ZN(n794) );
  XOR2_X1 U838 ( .A(G128), .B(n794), .Z(G30) );
  INV_X1 U839 ( .A(n795), .ZN(n796) );
  NAND2_X1 U840 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U841 ( .A(n798), .B(KEYINPUT116), .ZN(n799) );
  XNOR2_X1 U842 ( .A(G146), .B(n799), .ZN(G48) );
  XNOR2_X1 U843 ( .A(n800), .B(G125), .ZN(n801) );
  XNOR2_X1 U844 ( .A(n801), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 U845 ( .A(n802), .ZN(n803) );
  XOR2_X1 U846 ( .A(G134), .B(n803), .Z(G36) );
  NOR2_X1 U847 ( .A1(n665), .A2(n409), .ZN(n808) );
  NAND2_X1 U848 ( .A1(n409), .A2(G224), .ZN(n804) );
  XNOR2_X1 U849 ( .A(KEYINPUT61), .B(n804), .ZN(n805) );
  NAND2_X1 U850 ( .A1(n805), .A2(G898), .ZN(n806) );
  XNOR2_X1 U851 ( .A(n806), .B(KEYINPUT123), .ZN(n807) );
  NOR2_X1 U852 ( .A1(n808), .A2(n807), .ZN(n817) );
  BUF_X1 U853 ( .A(n809), .Z(n810) );
  XOR2_X1 U854 ( .A(KEYINPUT125), .B(n810), .Z(n813) );
  NOR2_X1 U855 ( .A1(n811), .A2(G898), .ZN(n812) );
  NOR2_X1 U856 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U857 ( .A(n814), .B(KEYINPUT126), .Z(n815) );
  XNOR2_X1 U858 ( .A(KEYINPUT124), .B(n815), .ZN(n816) );
  XNOR2_X1 U859 ( .A(n817), .B(n816), .ZN(G69) );
  XOR2_X1 U860 ( .A(n818), .B(G131), .Z(G33) );
  XOR2_X1 U861 ( .A(G137), .B(n819), .Z(G39) );
endmodule

