

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(n713), .A2(G299), .ZN(n516) );
  OR2_X1 U550 ( .A1(n689), .A2(n698), .ZN(n691) );
  XNOR2_X1 U551 ( .A(n516), .B(KEYINPUT92), .ZN(n702) );
  NAND2_X1 U552 ( .A1(n946), .A2(n703), .ZN(n705) );
  NOR2_X2 U553 ( .A1(n751), .A2(n747), .ZN(n726) );
  XNOR2_X2 U554 ( .A(n533), .B(KEYINPUT66), .ZN(n613) );
  XNOR2_X1 U555 ( .A(n691), .B(n690), .ZN(n695) );
  NOR2_X2 U556 ( .A1(n815), .A2(n814), .ZN(n816) );
  INV_X1 U557 ( .A(KEYINPUT91), .ZN(n690) );
  NOR2_X1 U558 ( .A1(G1966), .A2(n778), .ZN(n751) );
  NOR2_X1 U559 ( .A1(G2084), .A2(n697), .ZN(n747) );
  NOR2_X2 U560 ( .A1(n782), .A2(n688), .ZN(n698) );
  AND2_X1 U561 ( .A1(n771), .A2(n770), .ZN(n772) );
  INV_X1 U562 ( .A(G2104), .ZN(n524) );
  XNOR2_X1 U563 ( .A(n522), .B(KEYINPUT67), .ZN(n531) );
  NOR2_X1 U564 ( .A1(n778), .A2(n767), .ZN(n517) );
  XOR2_X1 U565 ( .A(n535), .B(n534), .Z(n518) );
  AND2_X1 U566 ( .A1(n887), .A2(G138), .ZN(n519) );
  AND2_X1 U567 ( .A1(n551), .A2(n550), .ZN(n520) );
  OR2_X1 U568 ( .A1(n768), .A2(n778), .ZN(n521) );
  INV_X1 U569 ( .A(KEYINPUT27), .ZN(n692) );
  XNOR2_X1 U570 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U571 ( .A(KEYINPUT30), .B(KEYINPUT94), .ZN(n727) );
  NOR2_X1 U572 ( .A1(G168), .A2(n729), .ZN(n730) );
  XNOR2_X1 U573 ( .A(KEYINPUT31), .B(KEYINPUT96), .ZN(n734) );
  XNOR2_X1 U574 ( .A(n735), .B(n734), .ZN(n736) );
  INV_X1 U575 ( .A(KEYINPUT97), .ZN(n743) );
  AND2_X1 U576 ( .A1(n769), .A2(n521), .ZN(n770) );
  OR2_X2 U577 ( .A1(n725), .A2(n724), .ZN(n778) );
  INV_X1 U578 ( .A(G2105), .ZN(n523) );
  AND2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n884) );
  NOR2_X1 U580 ( .A1(G651), .A2(n634), .ZN(n652) );
  OR2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n536) );
  NOR2_X1 U582 ( .A1(n536), .A2(n518), .ZN(n685) );
  BUF_X1 U583 ( .A(n685), .Z(G160) );
  NAND2_X1 U584 ( .A1(G113), .A2(n884), .ZN(n522) );
  NAND2_X1 U585 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X2 U586 ( .A(n525), .B(KEYINPUT17), .ZN(n887) );
  NAND2_X1 U587 ( .A1(G137), .A2(n887), .ZN(n529) );
  XNOR2_X2 U588 ( .A(G2104), .B(KEYINPUT65), .ZN(n532) );
  INV_X1 U589 ( .A(n532), .ZN(n527) );
  INV_X1 U590 ( .A(G2105), .ZN(n526) );
  NOR2_X2 U591 ( .A1(n527), .A2(n526), .ZN(n549) );
  BUF_X2 U592 ( .A(n549), .Z(n883) );
  NAND2_X1 U593 ( .A1(G125), .A2(n883), .ZN(n528) );
  NAND2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X2 U595 ( .A1(n532), .A2(G2105), .ZN(n533) );
  NAND2_X1 U596 ( .A1(n613), .A2(G101), .ZN(n535) );
  INV_X1 U597 ( .A(KEYINPUT23), .ZN(n534) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U599 ( .A1(n649), .A2(G89), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n537), .B(KEYINPUT4), .ZN(n539) );
  XOR2_X1 U601 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  INV_X1 U602 ( .A(G651), .ZN(n541) );
  NOR2_X1 U603 ( .A1(n634), .A2(n541), .ZN(n645) );
  NAND2_X1 U604 ( .A1(G76), .A2(n645), .ZN(n538) );
  NAND2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n540), .B(KEYINPUT5), .ZN(n547) );
  NOR2_X1 U607 ( .A1(G543), .A2(n541), .ZN(n542) );
  XOR2_X1 U608 ( .A(KEYINPUT1), .B(n542), .Z(n647) );
  NAND2_X1 U609 ( .A1(G63), .A2(n647), .ZN(n544) );
  NAND2_X1 U610 ( .A1(G51), .A2(n652), .ZN(n543) );
  NAND2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U612 ( .A(KEYINPUT6), .B(n545), .Z(n546) );
  NAND2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n548), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U615 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U616 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U617 ( .A(G120), .ZN(G236) );
  INV_X1 U618 ( .A(G69), .ZN(G235) );
  INV_X1 U619 ( .A(G108), .ZN(G238) );
  NAND2_X1 U620 ( .A1(n613), .A2(G102), .ZN(n552) );
  NAND2_X1 U621 ( .A1(G126), .A2(n549), .ZN(n551) );
  NAND2_X1 U622 ( .A1(G114), .A2(n884), .ZN(n550) );
  NAND2_X1 U623 ( .A1(n552), .A2(n520), .ZN(n553) );
  NOR2_X1 U624 ( .A1(n553), .A2(n519), .ZN(n686) );
  BUF_X1 U625 ( .A(n686), .Z(G164) );
  NAND2_X1 U626 ( .A1(G88), .A2(n649), .ZN(n555) );
  NAND2_X1 U627 ( .A1(G75), .A2(n645), .ZN(n554) );
  NAND2_X1 U628 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U629 ( .A1(G62), .A2(n647), .ZN(n557) );
  NAND2_X1 U630 ( .A1(G50), .A2(n652), .ZN(n556) );
  NAND2_X1 U631 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U632 ( .A1(n559), .A2(n558), .ZN(G166) );
  NAND2_X1 U633 ( .A1(G91), .A2(n649), .ZN(n561) );
  NAND2_X1 U634 ( .A1(G78), .A2(n645), .ZN(n560) );
  NAND2_X1 U635 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U636 ( .A1(n647), .A2(G65), .ZN(n562) );
  XOR2_X1 U637 ( .A(KEYINPUT70), .B(n562), .Z(n563) );
  NOR2_X1 U638 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U639 ( .A1(n652), .A2(G53), .ZN(n565) );
  NAND2_X1 U640 ( .A1(n566), .A2(n565), .ZN(G299) );
  NAND2_X1 U641 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U642 ( .A(n567), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U643 ( .A(G223), .ZN(n832) );
  NAND2_X1 U644 ( .A1(n832), .A2(G567), .ZN(n568) );
  XOR2_X1 U645 ( .A(KEYINPUT11), .B(n568), .Z(G234) );
  NAND2_X1 U646 ( .A1(G56), .A2(n647), .ZN(n569) );
  XNOR2_X1 U647 ( .A(n569), .B(KEYINPUT14), .ZN(n576) );
  NAND2_X1 U648 ( .A1(n649), .A2(G81), .ZN(n570) );
  XNOR2_X1 U649 ( .A(n570), .B(KEYINPUT12), .ZN(n572) );
  NAND2_X1 U650 ( .A1(G68), .A2(n645), .ZN(n571) );
  NAND2_X1 U651 ( .A1(n572), .A2(n571), .ZN(n574) );
  XOR2_X1 U652 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n573) );
  XNOR2_X1 U653 ( .A(n574), .B(n573), .ZN(n575) );
  NAND2_X1 U654 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U655 ( .A1(n652), .A2(G43), .ZN(n577) );
  XOR2_X1 U656 ( .A(KEYINPUT72), .B(n577), .Z(n578) );
  NOR2_X1 U657 ( .A1(n579), .A2(n578), .ZN(n947) );
  INV_X1 U658 ( .A(n947), .ZN(n606) );
  XNOR2_X1 U659 ( .A(G860), .B(KEYINPUT73), .ZN(n602) );
  OR2_X1 U660 ( .A1(n606), .A2(n602), .ZN(G153) );
  NAND2_X1 U661 ( .A1(G64), .A2(n647), .ZN(n581) );
  NAND2_X1 U662 ( .A1(G52), .A2(n652), .ZN(n580) );
  NAND2_X1 U663 ( .A1(n581), .A2(n580), .ZN(n586) );
  NAND2_X1 U664 ( .A1(G90), .A2(n649), .ZN(n583) );
  NAND2_X1 U665 ( .A1(G77), .A2(n645), .ZN(n582) );
  NAND2_X1 U666 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U667 ( .A(KEYINPUT9), .B(n584), .Z(n585) );
  NOR2_X1 U668 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U669 ( .A(KEYINPUT69), .B(n587), .ZN(G301) );
  NAND2_X1 U670 ( .A1(G868), .A2(G301), .ZN(n597) );
  NAND2_X1 U671 ( .A1(G66), .A2(n647), .ZN(n589) );
  NAND2_X1 U672 ( .A1(G92), .A2(n649), .ZN(n588) );
  NAND2_X1 U673 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U674 ( .A1(G79), .A2(n645), .ZN(n591) );
  NAND2_X1 U675 ( .A1(G54), .A2(n652), .ZN(n590) );
  NAND2_X1 U676 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U677 ( .A1(n593), .A2(n592), .ZN(n595) );
  XNOR2_X1 U678 ( .A(KEYINPUT74), .B(KEYINPUT15), .ZN(n594) );
  XNOR2_X1 U679 ( .A(n595), .B(n594), .ZN(n946) );
  INV_X1 U680 ( .A(n946), .ZN(n621) );
  OR2_X1 U681 ( .A1(n621), .A2(G868), .ZN(n596) );
  NAND2_X1 U682 ( .A1(n597), .A2(n596), .ZN(G284) );
  XNOR2_X1 U683 ( .A(KEYINPUT75), .B(G868), .ZN(n598) );
  NOR2_X1 U684 ( .A1(G286), .A2(n598), .ZN(n600) );
  NOR2_X1 U685 ( .A1(G868), .A2(G299), .ZN(n599) );
  NOR2_X1 U686 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U687 ( .A(KEYINPUT76), .B(n601), .ZN(G297) );
  NAND2_X1 U688 ( .A1(n602), .A2(G559), .ZN(n603) );
  NAND2_X1 U689 ( .A1(n603), .A2(n621), .ZN(n604) );
  XNOR2_X1 U690 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U691 ( .A1(G868), .A2(n621), .ZN(n605) );
  NOR2_X1 U692 ( .A1(G559), .A2(n605), .ZN(n608) );
  NOR2_X1 U693 ( .A1(G868), .A2(n606), .ZN(n607) );
  NOR2_X1 U694 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U695 ( .A1(G123), .A2(n883), .ZN(n609) );
  XOR2_X1 U696 ( .A(KEYINPUT18), .B(n609), .Z(n610) );
  XNOR2_X1 U697 ( .A(n610), .B(KEYINPUT77), .ZN(n612) );
  NAND2_X1 U698 ( .A1(G111), .A2(n884), .ZN(n611) );
  NAND2_X1 U699 ( .A1(n612), .A2(n611), .ZN(n618) );
  NAND2_X1 U700 ( .A1(G135), .A2(n887), .ZN(n616) );
  BUF_X1 U701 ( .A(n613), .Z(n614) );
  NAND2_X1 U702 ( .A1(G99), .A2(n614), .ZN(n615) );
  NAND2_X1 U703 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U704 ( .A1(n618), .A2(n617), .ZN(n1008) );
  XNOR2_X1 U705 ( .A(G2096), .B(n1008), .ZN(n620) );
  INV_X1 U706 ( .A(G2100), .ZN(n619) );
  NAND2_X1 U707 ( .A1(n620), .A2(n619), .ZN(G156) );
  XOR2_X1 U708 ( .A(n947), .B(KEYINPUT78), .Z(n623) );
  NAND2_X1 U709 ( .A1(G559), .A2(n621), .ZN(n622) );
  XNOR2_X1 U710 ( .A(n623), .B(n622), .ZN(n663) );
  NOR2_X1 U711 ( .A1(G860), .A2(n663), .ZN(n630) );
  NAND2_X1 U712 ( .A1(G67), .A2(n647), .ZN(n625) );
  NAND2_X1 U713 ( .A1(G93), .A2(n649), .ZN(n624) );
  NAND2_X1 U714 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U715 ( .A1(G80), .A2(n645), .ZN(n627) );
  NAND2_X1 U716 ( .A1(G55), .A2(n652), .ZN(n626) );
  NAND2_X1 U717 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U718 ( .A1(n629), .A2(n628), .ZN(n666) );
  XNOR2_X1 U719 ( .A(n630), .B(n666), .ZN(G145) );
  NAND2_X1 U720 ( .A1(G49), .A2(n652), .ZN(n632) );
  NAND2_X1 U721 ( .A1(G74), .A2(G651), .ZN(n631) );
  NAND2_X1 U722 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U723 ( .A1(n647), .A2(n633), .ZN(n637) );
  NAND2_X1 U724 ( .A1(G87), .A2(n634), .ZN(n635) );
  XOR2_X1 U725 ( .A(KEYINPUT79), .B(n635), .Z(n636) );
  NAND2_X1 U726 ( .A1(n637), .A2(n636), .ZN(G288) );
  NAND2_X1 U727 ( .A1(G85), .A2(n649), .ZN(n639) );
  NAND2_X1 U728 ( .A1(G72), .A2(n645), .ZN(n638) );
  NAND2_X1 U729 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U730 ( .A1(G60), .A2(n647), .ZN(n641) );
  NAND2_X1 U731 ( .A1(G47), .A2(n652), .ZN(n640) );
  NAND2_X1 U732 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U733 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U734 ( .A(KEYINPUT68), .B(n644), .Z(G290) );
  NAND2_X1 U735 ( .A1(G73), .A2(n645), .ZN(n646) );
  XNOR2_X1 U736 ( .A(n646), .B(KEYINPUT2), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n647), .A2(G61), .ZN(n648) );
  XNOR2_X1 U738 ( .A(n648), .B(KEYINPUT80), .ZN(n651) );
  NAND2_X1 U739 ( .A1(G86), .A2(n649), .ZN(n650) );
  NAND2_X1 U740 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U741 ( .A1(G48), .A2(n652), .ZN(n653) );
  XNOR2_X1 U742 ( .A(KEYINPUT81), .B(n653), .ZN(n654) );
  NOR2_X1 U743 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U744 ( .A1(n657), .A2(n656), .ZN(G305) );
  XNOR2_X1 U745 ( .A(KEYINPUT19), .B(G288), .ZN(n662) );
  XNOR2_X1 U746 ( .A(G166), .B(n666), .ZN(n660) );
  XOR2_X1 U747 ( .A(G290), .B(G305), .Z(n658) );
  XNOR2_X1 U748 ( .A(G299), .B(n658), .ZN(n659) );
  XNOR2_X1 U749 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U750 ( .A(n662), .B(n661), .ZN(n904) );
  XNOR2_X1 U751 ( .A(n904), .B(n663), .ZN(n664) );
  NAND2_X1 U752 ( .A1(n664), .A2(G868), .ZN(n665) );
  XNOR2_X1 U753 ( .A(n665), .B(KEYINPUT82), .ZN(n668) );
  OR2_X1 U754 ( .A1(G868), .A2(n666), .ZN(n667) );
  NAND2_X1 U755 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U756 ( .A1(G2084), .A2(G2078), .ZN(n669) );
  XNOR2_X1 U757 ( .A(n669), .B(KEYINPUT20), .ZN(n670) );
  XNOR2_X1 U758 ( .A(KEYINPUT83), .B(n670), .ZN(n671) );
  NAND2_X1 U759 ( .A1(n671), .A2(G2090), .ZN(n672) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U761 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U763 ( .A1(G483), .A2(G661), .ZN(n683) );
  NOR2_X1 U764 ( .A1(G235), .A2(G236), .ZN(n674) );
  XNOR2_X1 U765 ( .A(n674), .B(KEYINPUT85), .ZN(n675) );
  NOR2_X1 U766 ( .A1(G238), .A2(n675), .ZN(n676) );
  NAND2_X1 U767 ( .A1(G57), .A2(n676), .ZN(n838) );
  NAND2_X1 U768 ( .A1(n838), .A2(G567), .ZN(n682) );
  NAND2_X1 U769 ( .A1(G132), .A2(G82), .ZN(n677) );
  XNOR2_X1 U770 ( .A(n677), .B(KEYINPUT22), .ZN(n678) );
  XNOR2_X1 U771 ( .A(n678), .B(KEYINPUT84), .ZN(n679) );
  NOR2_X1 U772 ( .A1(G218), .A2(n679), .ZN(n680) );
  NAND2_X1 U773 ( .A1(G96), .A2(n680), .ZN(n839) );
  NAND2_X1 U774 ( .A1(n839), .A2(G2106), .ZN(n681) );
  NAND2_X1 U775 ( .A1(n682), .A2(n681), .ZN(n861) );
  NOR2_X1 U776 ( .A1(n683), .A2(n861), .ZN(n684) );
  XNOR2_X1 U777 ( .A(n684), .B(KEYINPUT86), .ZN(n837) );
  NAND2_X1 U778 ( .A1(G36), .A2(n837), .ZN(G176) );
  INV_X1 U779 ( .A(G166), .ZN(G303) );
  INV_X1 U780 ( .A(G1956), .ZN(n689) );
  NAND2_X1 U781 ( .A1(n685), .A2(G40), .ZN(n782) );
  NOR2_X2 U782 ( .A1(n686), .A2(G1384), .ZN(n687) );
  XNOR2_X1 U783 ( .A(n687), .B(KEYINPUT64), .ZN(n781) );
  INV_X1 U784 ( .A(n781), .ZN(n688) );
  NAND2_X1 U785 ( .A1(n698), .A2(G2072), .ZN(n693) );
  NAND2_X1 U786 ( .A1(n695), .A2(n694), .ZN(n713) );
  INV_X1 U787 ( .A(n698), .ZN(n697) );
  NAND2_X1 U788 ( .A1(G1348), .A2(n697), .ZN(n700) );
  BUF_X2 U789 ( .A(n698), .Z(n724) );
  NAND2_X1 U790 ( .A1(G2067), .A2(n724), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n700), .A2(n699), .ZN(n703) );
  NOR2_X1 U792 ( .A1(n703), .A2(n946), .ZN(n701) );
  NOR2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n711) );
  NAND2_X1 U794 ( .A1(G1341), .A2(n697), .ZN(n704) );
  NAND2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n708) );
  NAND2_X1 U796 ( .A1(G1996), .A2(n724), .ZN(n706) );
  XOR2_X1 U797 ( .A(KEYINPUT26), .B(n706), .Z(n707) );
  NOR2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U799 ( .A1(n947), .A2(n709), .ZN(n710) );
  NAND2_X1 U800 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U801 ( .A(n712), .B(KEYINPUT93), .ZN(n717) );
  BUF_X1 U802 ( .A(n713), .Z(n714) );
  NAND2_X1 U803 ( .A1(G299), .A2(n714), .ZN(n715) );
  XOR2_X1 U804 ( .A(KEYINPUT28), .B(n715), .Z(n716) );
  NOR2_X2 U805 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U806 ( .A(n718), .B(KEYINPUT29), .ZN(n723) );
  XOR2_X1 U807 ( .A(G2078), .B(KEYINPUT25), .Z(n719) );
  XNOR2_X1 U808 ( .A(KEYINPUT90), .B(n719), .ZN(n934) );
  NOR2_X1 U809 ( .A1(n697), .A2(n934), .ZN(n721) );
  NOR2_X1 U810 ( .A1(n724), .A2(G1961), .ZN(n720) );
  NOR2_X1 U811 ( .A1(n721), .A2(n720), .ZN(n731) );
  OR2_X1 U812 ( .A1(n731), .A2(G301), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n737) );
  INV_X1 U814 ( .A(G8), .ZN(n725) );
  NAND2_X1 U815 ( .A1(G8), .A2(n726), .ZN(n728) );
  XNOR2_X1 U816 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U817 ( .A(n730), .B(KEYINPUT95), .ZN(n733) );
  NAND2_X1 U818 ( .A1(n731), .A2(G301), .ZN(n732) );
  NAND2_X1 U819 ( .A1(n733), .A2(n732), .ZN(n735) );
  NAND2_X1 U820 ( .A1(n737), .A2(n736), .ZN(n748) );
  NAND2_X1 U821 ( .A1(n748), .A2(G286), .ZN(n742) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n778), .ZN(n739) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n697), .ZN(n738) );
  NOR2_X1 U824 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U825 ( .A1(n740), .A2(G303), .ZN(n741) );
  NAND2_X1 U826 ( .A1(n742), .A2(n741), .ZN(n744) );
  XNOR2_X1 U827 ( .A(n744), .B(n743), .ZN(n745) );
  NAND2_X1 U828 ( .A1(n745), .A2(G8), .ZN(n746) );
  XNOR2_X1 U829 ( .A(n746), .B(KEYINPUT32), .ZN(n755) );
  NAND2_X1 U830 ( .A1(G8), .A2(n747), .ZN(n753) );
  BUF_X1 U831 ( .A(n748), .Z(n749) );
  INV_X1 U832 ( .A(n749), .ZN(n750) );
  NOR2_X1 U833 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U834 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U835 ( .A1(n755), .A2(n754), .ZN(n766) );
  NOR2_X1 U836 ( .A1(G2090), .A2(G303), .ZN(n756) );
  NAND2_X1 U837 ( .A1(G8), .A2(n756), .ZN(n757) );
  NAND2_X1 U838 ( .A1(n766), .A2(n757), .ZN(n759) );
  INV_X1 U839 ( .A(KEYINPUT99), .ZN(n758) );
  XNOR2_X1 U840 ( .A(n759), .B(n758), .ZN(n760) );
  NAND2_X1 U841 ( .A1(n760), .A2(n778), .ZN(n774) );
  NOR2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n950) );
  NOR2_X1 U843 ( .A1(G1971), .A2(G303), .ZN(n761) );
  NOR2_X1 U844 ( .A1(n950), .A2(n761), .ZN(n762) );
  XNOR2_X1 U845 ( .A(n762), .B(KEYINPUT98), .ZN(n764) );
  INV_X1 U846 ( .A(KEYINPUT33), .ZN(n763) );
  AND2_X1 U847 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U848 ( .A1(n766), .A2(n765), .ZN(n771) );
  NAND2_X1 U849 ( .A1(G1976), .A2(G288), .ZN(n953) );
  INV_X1 U850 ( .A(n953), .ZN(n767) );
  OR2_X1 U851 ( .A1(KEYINPUT33), .A2(n517), .ZN(n769) );
  NAND2_X1 U852 ( .A1(n950), .A2(KEYINPUT33), .ZN(n768) );
  XOR2_X1 U853 ( .A(G1981), .B(G305), .Z(n965) );
  NAND2_X1 U854 ( .A1(n772), .A2(n965), .ZN(n773) );
  NAND2_X1 U855 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U856 ( .A(n775), .B(KEYINPUT100), .ZN(n780) );
  NOR2_X1 U857 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U858 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  NOR2_X1 U859 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U860 ( .A1(n780), .A2(n779), .ZN(n815) );
  BUF_X1 U861 ( .A(n781), .Z(n783) );
  NOR2_X1 U862 ( .A1(n783), .A2(n782), .ZN(n827) );
  XNOR2_X1 U863 ( .A(KEYINPUT37), .B(G2067), .ZN(n825) );
  NAND2_X1 U864 ( .A1(G140), .A2(n887), .ZN(n785) );
  NAND2_X1 U865 ( .A1(G104), .A2(n614), .ZN(n784) );
  NAND2_X1 U866 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U867 ( .A(KEYINPUT34), .B(n786), .ZN(n791) );
  NAND2_X1 U868 ( .A1(G128), .A2(n883), .ZN(n788) );
  NAND2_X1 U869 ( .A1(G116), .A2(n884), .ZN(n787) );
  NAND2_X1 U870 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U871 ( .A(KEYINPUT35), .B(n789), .Z(n790) );
  NOR2_X1 U872 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U873 ( .A(KEYINPUT36), .B(n792), .ZN(n901) );
  NOR2_X1 U874 ( .A1(n825), .A2(n901), .ZN(n1015) );
  NAND2_X1 U875 ( .A1(n827), .A2(n1015), .ZN(n793) );
  XOR2_X1 U876 ( .A(KEYINPUT87), .B(n793), .Z(n823) );
  NAND2_X1 U877 ( .A1(G129), .A2(n883), .ZN(n795) );
  NAND2_X1 U878 ( .A1(G117), .A2(n884), .ZN(n794) );
  NAND2_X1 U879 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U880 ( .A(KEYINPUT88), .B(n796), .ZN(n799) );
  NAND2_X1 U881 ( .A1(G105), .A2(n614), .ZN(n797) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(n797), .Z(n798) );
  NOR2_X1 U883 ( .A1(n799), .A2(n798), .ZN(n801) );
  NAND2_X1 U884 ( .A1(n887), .A2(G141), .ZN(n800) );
  NAND2_X1 U885 ( .A1(n801), .A2(n800), .ZN(n900) );
  NAND2_X1 U886 ( .A1(G1996), .A2(n900), .ZN(n809) );
  NAND2_X1 U887 ( .A1(G131), .A2(n887), .ZN(n803) );
  NAND2_X1 U888 ( .A1(G119), .A2(n883), .ZN(n802) );
  NAND2_X1 U889 ( .A1(n803), .A2(n802), .ZN(n807) );
  NAND2_X1 U890 ( .A1(n884), .A2(G107), .ZN(n805) );
  NAND2_X1 U891 ( .A1(G95), .A2(n614), .ZN(n804) );
  NAND2_X1 U892 ( .A1(n805), .A2(n804), .ZN(n806) );
  OR2_X1 U893 ( .A1(n807), .A2(n806), .ZN(n872) );
  NAND2_X1 U894 ( .A1(G1991), .A2(n872), .ZN(n808) );
  NAND2_X1 U895 ( .A1(n809), .A2(n808), .ZN(n1011) );
  NAND2_X1 U896 ( .A1(n827), .A2(n1011), .ZN(n810) );
  NAND2_X1 U897 ( .A1(n823), .A2(n810), .ZN(n811) );
  XNOR2_X1 U898 ( .A(n811), .B(KEYINPUT89), .ZN(n813) );
  XNOR2_X1 U899 ( .A(G1986), .B(G290), .ZN(n956) );
  NAND2_X1 U900 ( .A1(n827), .A2(n956), .ZN(n812) );
  NAND2_X1 U901 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U902 ( .A(n816), .B(KEYINPUT101), .ZN(n830) );
  NOR2_X1 U903 ( .A1(n900), .A2(G1996), .ZN(n817) );
  XNOR2_X1 U904 ( .A(n817), .B(KEYINPUT102), .ZN(n1019) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n872), .ZN(n1009) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U907 ( .A1(n1009), .A2(n818), .ZN(n819) );
  NOR2_X1 U908 ( .A1(n819), .A2(n1011), .ZN(n820) );
  NOR2_X1 U909 ( .A1(n1019), .A2(n820), .ZN(n821) );
  XOR2_X1 U910 ( .A(n821), .B(KEYINPUT39), .Z(n822) );
  XNOR2_X1 U911 ( .A(KEYINPUT103), .B(n822), .ZN(n824) );
  NAND2_X1 U912 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U913 ( .A1(n825), .A2(n901), .ZN(n1022) );
  NAND2_X1 U914 ( .A1(n826), .A2(n1022), .ZN(n828) );
  NAND2_X1 U915 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U916 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U917 ( .A(n831), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n832), .ZN(G217) );
  INV_X1 U919 ( .A(G661), .ZN(n834) );
  NAND2_X1 U920 ( .A1(G2), .A2(G15), .ZN(n833) );
  NOR2_X1 U921 ( .A1(n834), .A2(n833), .ZN(n835) );
  XOR2_X1 U922 ( .A(KEYINPUT104), .B(n835), .Z(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U924 ( .A1(n837), .A2(n836), .ZN(G188) );
  NOR2_X1 U925 ( .A1(n839), .A2(n838), .ZN(G325) );
  XNOR2_X1 U926 ( .A(KEYINPUT105), .B(G325), .ZN(G261) );
  INV_X1 U928 ( .A(G132), .ZN(G219) );
  INV_X1 U929 ( .A(G82), .ZN(G220) );
  XOR2_X1 U930 ( .A(KEYINPUT108), .B(KEYINPUT106), .Z(n841) );
  XNOR2_X1 U931 ( .A(KEYINPUT107), .B(G2096), .ZN(n840) );
  XNOR2_X1 U932 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U933 ( .A(n842), .B(KEYINPUT42), .Z(n844) );
  XNOR2_X1 U934 ( .A(G2067), .B(G2090), .ZN(n843) );
  XNOR2_X1 U935 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U936 ( .A(G2100), .B(G2072), .Z(n846) );
  XNOR2_X1 U937 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U938 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U939 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U940 ( .A(KEYINPUT43), .B(G2678), .ZN(n849) );
  XNOR2_X1 U941 ( .A(n850), .B(n849), .ZN(G227) );
  XOR2_X1 U942 ( .A(G1971), .B(G1961), .Z(n852) );
  XNOR2_X1 U943 ( .A(G1986), .B(G1966), .ZN(n851) );
  XNOR2_X1 U944 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U945 ( .A(G1976), .B(G1956), .Z(n854) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1991), .ZN(n853) );
  XNOR2_X1 U947 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U948 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U949 ( .A(KEYINPUT109), .B(G2474), .ZN(n857) );
  XNOR2_X1 U950 ( .A(n858), .B(n857), .ZN(n860) );
  XOR2_X1 U951 ( .A(G1981), .B(KEYINPUT41), .Z(n859) );
  XNOR2_X1 U952 ( .A(n860), .B(n859), .ZN(G229) );
  INV_X1 U953 ( .A(n861), .ZN(G319) );
  NAND2_X1 U954 ( .A1(n887), .A2(G136), .ZN(n862) );
  XNOR2_X1 U955 ( .A(KEYINPUT110), .B(n862), .ZN(n865) );
  NAND2_X1 U956 ( .A1(n883), .A2(G124), .ZN(n863) );
  XNOR2_X1 U957 ( .A(KEYINPUT44), .B(n863), .ZN(n864) );
  NAND2_X1 U958 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U959 ( .A(n866), .B(KEYINPUT111), .ZN(n868) );
  NAND2_X1 U960 ( .A1(G112), .A2(n884), .ZN(n867) );
  NAND2_X1 U961 ( .A1(n868), .A2(n867), .ZN(n871) );
  NAND2_X1 U962 ( .A1(n614), .A2(G100), .ZN(n869) );
  XOR2_X1 U963 ( .A(KEYINPUT112), .B(n869), .Z(n870) );
  NOR2_X1 U964 ( .A1(n871), .A2(n870), .ZN(G162) );
  XNOR2_X1 U965 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n874) );
  XNOR2_X1 U966 ( .A(n872), .B(KEYINPUT46), .ZN(n873) );
  XNOR2_X1 U967 ( .A(n874), .B(n873), .ZN(n898) );
  XNOR2_X1 U968 ( .A(G160), .B(G162), .ZN(n882) );
  NAND2_X1 U969 ( .A1(G139), .A2(n887), .ZN(n876) );
  NAND2_X1 U970 ( .A1(G103), .A2(n614), .ZN(n875) );
  NAND2_X1 U971 ( .A1(n876), .A2(n875), .ZN(n881) );
  NAND2_X1 U972 ( .A1(G127), .A2(n883), .ZN(n878) );
  NAND2_X1 U973 ( .A1(G115), .A2(n884), .ZN(n877) );
  NAND2_X1 U974 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U975 ( .A(KEYINPUT47), .B(n879), .Z(n880) );
  NOR2_X1 U976 ( .A1(n881), .A2(n880), .ZN(n1004) );
  XNOR2_X1 U977 ( .A(n882), .B(n1004), .ZN(n894) );
  NAND2_X1 U978 ( .A1(G130), .A2(n883), .ZN(n886) );
  NAND2_X1 U979 ( .A1(G118), .A2(n884), .ZN(n885) );
  NAND2_X1 U980 ( .A1(n886), .A2(n885), .ZN(n892) );
  NAND2_X1 U981 ( .A1(G142), .A2(n887), .ZN(n889) );
  NAND2_X1 U982 ( .A1(G106), .A2(n614), .ZN(n888) );
  NAND2_X1 U983 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U984 ( .A(KEYINPUT45), .B(n890), .Z(n891) );
  NOR2_X1 U985 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U986 ( .A(n894), .B(n893), .Z(n896) );
  XNOR2_X1 U987 ( .A(G164), .B(n1008), .ZN(n895) );
  XNOR2_X1 U988 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U989 ( .A(n898), .B(n897), .Z(n899) );
  XNOR2_X1 U990 ( .A(n900), .B(n899), .ZN(n902) );
  XOR2_X1 U991 ( .A(n902), .B(n901), .Z(n903) );
  NOR2_X1 U992 ( .A1(G37), .A2(n903), .ZN(G395) );
  INV_X1 U993 ( .A(G301), .ZN(G171) );
  XOR2_X1 U994 ( .A(n904), .B(G286), .Z(n906) );
  XNOR2_X1 U995 ( .A(n947), .B(n946), .ZN(n905) );
  XNOR2_X1 U996 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U997 ( .A(G171), .B(n907), .ZN(n908) );
  NOR2_X1 U998 ( .A1(G37), .A2(n908), .ZN(G397) );
  NOR2_X1 U999 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1000 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(n910), .B(n909), .ZN(n921) );
  XOR2_X1 U1002 ( .A(G2451), .B(G2430), .Z(n912) );
  XNOR2_X1 U1003 ( .A(G2438), .B(G2443), .ZN(n911) );
  XNOR2_X1 U1004 ( .A(n912), .B(n911), .ZN(n918) );
  XOR2_X1 U1005 ( .A(G2435), .B(G2454), .Z(n914) );
  XNOR2_X1 U1006 ( .A(G1348), .B(G1341), .ZN(n913) );
  XNOR2_X1 U1007 ( .A(n914), .B(n913), .ZN(n916) );
  XOR2_X1 U1008 ( .A(G2446), .B(G2427), .Z(n915) );
  XNOR2_X1 U1009 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1010 ( .A(n918), .B(n917), .Z(n919) );
  NAND2_X1 U1011 ( .A1(G14), .A2(n919), .ZN(n924) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n924), .ZN(n920) );
  NOR2_X1 U1013 ( .A1(n921), .A2(n920), .ZN(n923) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1015 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G96), .ZN(G221) );
  INV_X1 U1018 ( .A(G57), .ZN(G237) );
  INV_X1 U1019 ( .A(n924), .ZN(G401) );
  XOR2_X1 U1020 ( .A(G2090), .B(G35), .Z(n927) );
  XOR2_X1 U1021 ( .A(G34), .B(KEYINPUT54), .Z(n925) );
  XNOR2_X1 U1022 ( .A(n925), .B(G2084), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n943) );
  XNOR2_X1 U1024 ( .A(G25), .B(G1991), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(n928), .B(KEYINPUT117), .ZN(n933) );
  XOR2_X1 U1026 ( .A(G2067), .B(G26), .Z(n929) );
  NAND2_X1 U1027 ( .A1(n929), .A2(G28), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(G33), .B(G2072), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n939) );
  XNOR2_X1 U1031 ( .A(n934), .B(G27), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(G32), .B(G1996), .ZN(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1034 ( .A(n937), .B(KEYINPUT118), .Z(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1036 ( .A(KEYINPUT53), .B(n940), .Z(n941) );
  XNOR2_X1 U1037 ( .A(n941), .B(KEYINPUT119), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1039 ( .A(KEYINPUT55), .B(n944), .Z(n945) );
  NOR2_X1 U1040 ( .A1(G29), .A2(n945), .ZN(n1001) );
  XNOR2_X1 U1041 ( .A(G16), .B(KEYINPUT56), .ZN(n971) );
  XOR2_X1 U1042 ( .A(n946), .B(G1348), .Z(n949) );
  XNOR2_X1 U1043 ( .A(n947), .B(G1341), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n963) );
  XNOR2_X1 U1045 ( .A(G171), .B(G1961), .ZN(n961) );
  XNOR2_X1 U1046 ( .A(G299), .B(G1956), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(n950), .B(KEYINPUT120), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(G166), .B(G1971), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(KEYINPUT121), .B(n959), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(KEYINPUT122), .B(n964), .ZN(n969) );
  XNOR2_X1 U1057 ( .A(G1966), .B(G168), .ZN(n966) );
  NAND2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(KEYINPUT57), .B(n967), .ZN(n968) );
  NAND2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1061 ( .A1(n971), .A2(n970), .ZN(n998) );
  INV_X1 U1062 ( .A(G16), .ZN(n996) );
  XNOR2_X1 U1063 ( .A(KEYINPUT123), .B(G1961), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(n972), .B(G5), .ZN(n986) );
  XNOR2_X1 U1065 ( .A(KEYINPUT125), .B(G1341), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(n973), .B(G19), .ZN(n978) );
  XOR2_X1 U1067 ( .A(G1348), .B(KEYINPUT59), .Z(n974) );
  XNOR2_X1 U1068 ( .A(G4), .B(n974), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(G6), .B(G1981), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(G20), .B(G1956), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(KEYINPUT124), .B(n979), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1075 ( .A(KEYINPUT60), .B(n982), .Z(n984) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G21), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n993) );
  XNOR2_X1 U1079 ( .A(G1971), .B(G22), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(G23), .B(G1976), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n990) );
  XOR2_X1 U1082 ( .A(G1986), .B(G24), .Z(n989) );
  NAND2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(KEYINPUT58), .B(n991), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(KEYINPUT61), .B(n994), .ZN(n995) );
  NAND2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(n999), .B(KEYINPUT126), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(G11), .A2(n1002), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(KEYINPUT127), .B(n1003), .Z(n1032) );
  XOR2_X1 U1093 ( .A(G2072), .B(n1004), .Z(n1006) );
  XOR2_X1 U1094 ( .A(G164), .B(G2078), .Z(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1007), .ZN(n1017) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1013) );
  XOR2_X1 U1098 ( .A(G160), .B(G2084), .Z(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1025) );
  XOR2_X1 U1103 ( .A(G2090), .B(G162), .Z(n1018) );
  NOR2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(KEYINPUT115), .B(n1020), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(n1021), .B(KEYINPUT51), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1109 ( .A(KEYINPUT52), .B(n1026), .ZN(n1028) );
  INV_X1 U1110 ( .A(KEYINPUT55), .ZN(n1027) );
  NAND2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1112 ( .A1(n1029), .A2(G29), .ZN(n1030) );
  XOR2_X1 U1113 ( .A(KEYINPUT116), .B(n1030), .Z(n1031) );
  NOR2_X1 U1114 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1033), .ZN(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

