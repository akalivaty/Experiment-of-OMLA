//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n557, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n603, new_n605,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1087, new_n1088,
    new_n1089;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT64), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT65), .Z(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  AND3_X1   g040(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT66), .ZN(new_n466));
  AOI21_X1  g041(.A(KEYINPUT66), .B1(new_n463), .B2(new_n465), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n461), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n464), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n472));
  NOR3_X1   g047(.A1(new_n471), .A2(new_n472), .A3(G2105), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n462), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT67), .ZN(new_n477));
  NOR3_X1   g052(.A1(new_n470), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT68), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n473), .A2(G136), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n463), .A2(new_n465), .A3(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n461), .B2(G112), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n481), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT69), .Z(G162));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT70), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G114), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n482), .A2(G126), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(KEYINPUT71), .B2(G2105), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(new_n471), .B2(new_n472), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT66), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n461), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n495), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT72), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n495), .B(new_n510), .C1(new_n505), .C2(new_n507), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(G164));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT73), .B1(new_n517), .B2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(new_n520), .A3(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n517), .A2(KEYINPUT5), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(new_n513), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n516), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(G62), .ZN(new_n529));
  NAND2_X1  g104(.A1(G75), .A2(G543), .ZN(new_n530));
  XOR2_X1   g105(.A(new_n530), .B(KEYINPUT74), .Z(new_n531));
  AOI21_X1  g106(.A(new_n528), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n527), .A2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  INV_X1    g109(.A(new_n525), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G89), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XOR2_X1   g113(.A(new_n538), .B(KEYINPUT7), .Z(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(G51), .B2(new_n515), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(G168));
  XOR2_X1   g117(.A(KEYINPUT75), .B(G52), .Z(new_n543));
  AOI22_X1  g118(.A1(new_n535), .A2(G90), .B1(new_n515), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n528), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  AOI22_X1  g123(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n528), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(KEYINPUT76), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n535), .A2(G81), .B1(G43), .B2(new_n515), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n550), .A2(KEYINPUT76), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n522), .A2(new_n523), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n535), .A2(G91), .B1(new_n565), .B2(G651), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n515), .A2(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n567), .B1(KEYINPUT77), .B2(KEYINPUT9), .ZN(new_n568));
  XOR2_X1   g143(.A(KEYINPUT77), .B(KEYINPUT9), .Z(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G299));
  XOR2_X1   g146(.A(new_n541), .B(KEYINPUT78), .Z(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G286));
  NAND2_X1  g148(.A1(new_n535), .A2(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n515), .A2(G49), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  AOI22_X1  g152(.A1(new_n524), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n578));
  OR3_X1    g153(.A1(new_n578), .A2(KEYINPUT79), .A3(new_n528), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT79), .B1(new_n578), .B2(new_n528), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n579), .A2(new_n580), .B1(G86), .B2(new_n535), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n515), .A2(G48), .ZN(new_n582));
  XOR2_X1   g157(.A(new_n582), .B(KEYINPUT80), .Z(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n535), .A2(G85), .B1(G47), .B2(new_n515), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n528), .B2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n535), .A2(G92), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n515), .A2(G54), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT81), .Z(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n524), .B2(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n591), .B1(new_n594), .B2(new_n528), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n588), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n588), .B1(new_n596), .B2(G868), .ZN(G321));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(G299), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(new_n572), .B2(new_n599), .ZN(G297));
  OAI21_X1  g176(.A(new_n600), .B1(new_n572), .B2(new_n599), .ZN(G280));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n596), .B1(new_n603), .B2(G860), .ZN(G148));
  NAND2_X1  g179(.A1(new_n554), .A2(new_n599), .ZN(new_n605));
  INV_X1    g180(.A(new_n596), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n605), .B1(new_n607), .B2(new_n599), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g184(.A(new_n475), .B1(new_n466), .B2(new_n467), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(G2100), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(G2100), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n473), .A2(G135), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n482), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(G99), .A2(G2105), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT83), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2096), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n614), .A2(new_n615), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT84), .Z(G156));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT85), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2427), .B(G2430), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT14), .ZN(new_n630));
  XOR2_X1   g205(.A(G2451), .B(G2454), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT86), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n630), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G14), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(G401));
  XOR2_X1   g215(.A(G2072), .B(G2078), .Z(new_n641));
  XOR2_X1   g216(.A(G2067), .B(G2678), .Z(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n641), .B1(new_n645), .B2(KEYINPUT18), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2096), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2100), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n645), .A2(KEYINPUT17), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n643), .A2(new_n644), .ZN(new_n650));
  AOI21_X1  g225(.A(KEYINPUT18), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n648), .B(new_n651), .Z(G227));
  XOR2_X1   g227(.A(G1956), .B(G2474), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT87), .ZN(new_n654));
  XOR2_X1   g229(.A(G1961), .B(G1966), .Z(new_n655));
  AND2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT20), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n654), .A2(new_n655), .ZN(new_n661));
  AOI22_X1  g236(.A1(new_n659), .A2(new_n660), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  OR3_X1    g237(.A1(new_n656), .A2(new_n661), .A3(new_n658), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n662), .B(new_n663), .C1(new_n660), .C2(new_n659), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(G1986), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1991), .B(G1996), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT22), .B(G1981), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G229));
  MUX2_X1   g245(.A(G6), .B(G305), .S(G16), .Z(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT32), .B(G1981), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G22), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(G166), .B2(new_n676), .ZN(new_n678));
  INV_X1    g253(.A(G1971), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(G16), .A2(G23), .ZN(new_n681));
  INV_X1    g256(.A(G288), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(G16), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT33), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n675), .A2(new_n680), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT91), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT34), .ZN(new_n688));
  MUX2_X1   g263(.A(G24), .B(G290), .S(G16), .Z(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(G1986), .Z(new_n690));
  INV_X1    g265(.A(KEYINPUT92), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT36), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(G25), .A2(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n473), .A2(G131), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n482), .A2(G119), .ZN(new_n696));
  NOR2_X1   g271(.A1(G95), .A2(G2105), .ZN(new_n697));
  OAI21_X1  g272(.A(G2104), .B1(new_n461), .B2(G107), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n695), .B(new_n696), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT88), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n694), .B1(new_n700), .B2(G29), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT35), .B(G1991), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n693), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n688), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n691), .A2(new_n692), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(G26), .ZN(new_n711));
  OAI21_X1  g286(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n712));
  INV_X1    g287(.A(G104), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n461), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT95), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n482), .A2(G128), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n473), .A2(G140), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n711), .B1(new_n718), .B2(G29), .ZN(new_n719));
  MUX2_X1   g294(.A(new_n711), .B(new_n719), .S(KEYINPUT28), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT96), .B(G2067), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT24), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(G34), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(G34), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n724), .A2(new_n725), .A3(new_n710), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n479), .B2(new_n710), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(G2084), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n676), .A2(G20), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT100), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT23), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G299), .B2(G16), .ZN(new_n732));
  INV_X1    g307(.A(G1956), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n676), .A2(G4), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n596), .B2(new_n676), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT93), .B(G1348), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G29), .A2(G35), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G162), .B2(G29), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT29), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n735), .B(new_n739), .C1(G2090), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n710), .A2(G32), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n473), .A2(G141), .B1(new_n482), .B2(G129), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n475), .A2(G105), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT26), .Z(new_n748));
  NAND3_X1  g323(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT99), .Z(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n744), .B1(new_n751), .B2(new_n710), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT27), .B(G1996), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G27), .A2(G29), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G164), .B2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2078), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(KEYINPUT97), .B1(G29), .B2(G33), .ZN(new_n759));
  OR3_X1    g334(.A1(KEYINPUT97), .A2(G29), .A3(G33), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n475), .A2(G103), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT25), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n473), .A2(G139), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT98), .Z(new_n765));
  INV_X1    g340(.A(G127), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n503), .B2(new_n504), .ZN(new_n767));
  AND2_X1   g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  OAI21_X1  g343(.A(G2105), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n759), .B(new_n760), .C1(new_n770), .C2(new_n710), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G2072), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n742), .A2(G2090), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT31), .B(G11), .Z(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT30), .B(G28), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n710), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n758), .A2(new_n772), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G21), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G168), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1966), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n620), .A2(new_n710), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n743), .A2(new_n777), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n708), .A2(new_n709), .A3(new_n722), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n676), .A2(G5), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G171), .B2(new_n676), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1961), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n676), .A2(G19), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n555), .B2(new_n676), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT94), .B(G1341), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n783), .A2(new_n786), .A3(new_n790), .ZN(G311));
  AND3_X1   g366(.A1(new_n708), .A2(new_n709), .A3(new_n782), .ZN(new_n792));
  INV_X1    g367(.A(new_n786), .ZN(new_n793));
  INV_X1    g368(.A(new_n790), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n792), .A2(new_n793), .A3(new_n794), .A4(new_n722), .ZN(G150));
  AOI22_X1  g370(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n796), .A2(new_n528), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n515), .A2(G55), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT103), .B(G93), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n525), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(G860), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT37), .Z(new_n802));
  NOR2_X1   g377(.A1(new_n606), .A2(new_n603), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n797), .A2(new_n800), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n554), .B(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n803), .B(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT102), .B(KEYINPUT104), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT39), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n808), .B(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n802), .B1(new_n811), .B2(G860), .ZN(G145));
  NAND2_X1  g387(.A1(new_n770), .A2(new_n749), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n750), .B2(new_n770), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n718), .B(new_n508), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n699), .B(KEYINPUT105), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n473), .A2(G142), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n482), .A2(G130), .ZN(new_n819));
  NOR2_X1   g394(.A1(G106), .A2(G2105), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n818), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n817), .B(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(new_n612), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n816), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT106), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n479), .B(new_n620), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G162), .ZN(new_n828));
  INV_X1    g403(.A(new_n816), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n824), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n826), .B(new_n828), .C1(KEYINPUT106), .C2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(G37), .ZN(new_n832));
  INV_X1    g407(.A(new_n825), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n831), .B(new_n832), .C1(new_n833), .C2(new_n828), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g410(.A(G303), .B(G288), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G290), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G305), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT42), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n596), .B(G299), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT41), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n607), .B(new_n805), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n840), .B(KEYINPUT107), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n839), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G868), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(G868), .B2(new_n804), .ZN(G295));
  OAI21_X1  g423(.A(new_n847), .B1(G868), .B2(new_n804), .ZN(G331));
  NAND2_X1  g424(.A1(G168), .A2(G301), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n572), .B2(G301), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(new_n805), .Z(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(new_n841), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n840), .B2(new_n852), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(new_n838), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n838), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n855), .A2(new_n832), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(KEYINPUT43), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n853), .B1(new_n844), .B2(new_n852), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n856), .B(new_n832), .C1(new_n838), .C2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT43), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(KEYINPUT44), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n857), .A2(KEYINPUT43), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n860), .A2(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n863), .B1(KEYINPUT44), .B2(new_n866), .ZN(G397));
  INV_X1    g442(.A(G40), .ZN(new_n868));
  NOR4_X1   g443(.A1(new_n470), .A2(new_n868), .A3(new_n474), .A4(new_n477), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(G1384), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n508), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT45), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(G1996), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n751), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT108), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n875), .B(KEYINPUT109), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G2067), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n718), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n749), .A2(G1996), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n879), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n699), .B(new_n702), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n880), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(G290), .B(G1986), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n891), .B1(new_n875), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n872), .A2(KEYINPUT50), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n870), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n509), .A2(new_n871), .A3(new_n511), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT50), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT117), .ZN(new_n899));
  INV_X1    g474(.A(G1348), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT117), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n895), .A2(new_n901), .A3(new_n897), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n870), .A2(new_n872), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n882), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(KEYINPUT60), .A3(new_n905), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n906), .A2(KEYINPUT124), .A3(new_n606), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n606), .B1(new_n906), .B2(KEYINPUT124), .ZN(new_n908));
  OAI22_X1  g483(.A1(new_n907), .A2(new_n908), .B1(KEYINPUT124), .B2(new_n906), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n903), .A2(new_n905), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n909), .B1(KEYINPUT60), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n566), .B(KEYINPUT115), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n912), .A2(new_n570), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT116), .B1(new_n913), .B2(KEYINPUT57), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT57), .ZN(new_n915));
  NOR2_X1   g490(.A1(G299), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n912), .A2(new_n570), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT116), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n915), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n914), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n872), .A2(KEYINPUT50), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n869), .B(new_n922), .C1(new_n896), .C2(KEYINPUT50), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n733), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n896), .A2(new_n873), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n871), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT110), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n508), .A2(new_n928), .A3(KEYINPUT45), .A4(new_n871), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n869), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(KEYINPUT56), .B(G2072), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n921), .A2(new_n924), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n924), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n914), .A2(new_n935), .A3(new_n917), .A4(new_n920), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT61), .ZN(new_n938));
  XNOR2_X1  g513(.A(KEYINPUT119), .B(G1996), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n925), .A2(new_n930), .A3(new_n939), .ZN(new_n940));
  XOR2_X1   g515(.A(KEYINPUT58), .B(G1341), .Z(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n870), .B2(new_n872), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT120), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n930), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n896), .A2(new_n873), .ZN(new_n946));
  INV_X1    g521(.A(new_n939), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT120), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n949), .A3(new_n942), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n944), .A2(new_n555), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT121), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT121), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n944), .A2(new_n950), .A3(new_n953), .A4(new_n555), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(KEYINPUT59), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT59), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n944), .A2(new_n950), .A3(new_n956), .A4(new_n555), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n957), .A2(KEYINPUT122), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT123), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT122), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n952), .A2(new_n961), .A3(KEYINPUT59), .A4(new_n954), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n960), .B1(new_n959), .B2(new_n962), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n911), .B(new_n938), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT125), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n936), .B1(new_n910), .B2(new_n606), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n934), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT118), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n965), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n966), .B1(new_n965), .B2(new_n969), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n869), .B(new_n874), .C1(new_n896), .C2(new_n873), .ZN(new_n972));
  INV_X1    g547(.A(G1966), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT113), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(G2084), .B2(new_n898), .ZN(new_n976));
  OAI21_X1  g551(.A(G8), .B1(new_n976), .B2(new_n541), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT51), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n979), .B1(new_n976), .B2(new_n541), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G2078), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT53), .B1(new_n931), .B2(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n899), .A2(new_n902), .ZN(new_n984));
  INV_X1    g559(.A(G1961), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n982), .A2(KEYINPUT53), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n986), .B1(new_n972), .B2(new_n987), .ZN(new_n988));
  OR2_X1    g563(.A1(G171), .A2(KEYINPUT54), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT126), .B(KEYINPUT54), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n988), .B(new_n989), .C1(G301), .C2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n981), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(G305), .A2(G1981), .ZN(new_n993));
  INV_X1    g568(.A(G1981), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n581), .A2(new_n994), .A3(new_n583), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT49), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G8), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n904), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n993), .A2(KEYINPUT49), .A3(new_n995), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1976), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1000), .B1(new_n1003), .B2(G288), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT52), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT111), .B(G1976), .Z(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT52), .B1(G288), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1000), .B(new_n1007), .C1(new_n1003), .C2(G288), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1002), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n898), .A2(G2090), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n679), .B1(new_n925), .B2(new_n930), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(G8), .ZN(new_n1013));
  NAND2_X1  g588(.A1(G303), .A2(G8), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT55), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1011), .B1(G2090), .B2(new_n923), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(G8), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1018), .A2(new_n1015), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1009), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(G171), .A2(new_n990), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n874), .A2(KEYINPUT53), .A3(new_n982), .ZN(new_n1022));
  OAI221_X1 g597(.A(new_n986), .B1(KEYINPUT54), .B2(G301), .C1(new_n930), .C2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1020), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n992), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n970), .A2(new_n971), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1009), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n1016), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1002), .A2(new_n1003), .A3(new_n682), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n995), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT112), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1030), .A2(new_n1033), .A3(new_n995), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1000), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n976), .A2(G8), .A3(new_n572), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT63), .B1(new_n1020), .B2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1009), .A2(new_n1016), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT63), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(new_n1037), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1029), .B(new_n1035), .C1(new_n1038), .C2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1016), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1019), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1028), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1040), .B1(new_n1049), .B2(new_n1036), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n1042), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1051), .A2(KEYINPUT114), .A3(new_n1029), .A4(new_n1035), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1046), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(G301), .B1(new_n981), .B2(KEYINPUT62), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT62), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n978), .B(new_n1055), .C1(new_n977), .C2(new_n980), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1054), .A2(new_n988), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n1020), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1053), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n893), .B1(new_n1027), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT127), .ZN(new_n1061));
  INV_X1    g636(.A(new_n702), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n888), .A2(new_n1062), .A3(new_n700), .ZN(new_n1063));
  OR2_X1    g638(.A1(new_n718), .A2(G2067), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n880), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n876), .A2(G1986), .A3(G290), .ZN(new_n1066));
  XOR2_X1   g641(.A(new_n1066), .B(KEYINPUT48), .Z(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n891), .A2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n877), .B(KEYINPUT46), .ZN(new_n1070));
  OR2_X1    g645(.A1(new_n884), .A2(new_n749), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n881), .B2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1072), .B(KEYINPUT47), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1065), .A2(new_n1069), .A3(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1060), .A2(new_n1061), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n893), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n965), .A2(new_n969), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT125), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n965), .A2(new_n966), .A3(new_n969), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(new_n1025), .A3(new_n1079), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1046), .A2(new_n1052), .B1(new_n1057), .B2(new_n1020), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1076), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1074), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT127), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1075), .A2(new_n1084), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g660(.A1(new_n864), .A2(G319), .A3(new_n834), .A4(new_n865), .ZN(new_n1087));
  NOR3_X1   g661(.A1(G229), .A2(G401), .A3(G227), .ZN(new_n1088));
  INV_X1    g662(.A(new_n1088), .ZN(new_n1089));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1089), .ZN(G308));
  INV_X1    g664(.A(G308), .ZN(G225));
endmodule


