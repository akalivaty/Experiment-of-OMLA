// Benchmark "locked_c1355" written by ABC on Sat Dec 16 10:33:07 2023

module locked_c1355 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat,
    G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat,
    G85gat, G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat,
    G141gat, G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat,
    G197gat, G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat,
    G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat,
    G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat,
    G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat, G120gat,
    G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat, G176gat,
    G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat, G226gat,
    G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n138, new_n139, new_n140, new_n141, new_n142, new_n143, new_n144,
    new_n145, new_n146, new_n147, new_n148, new_n149, new_n150, new_n151,
    new_n152, new_n153, new_n154, new_n155, new_n156, new_n157, new_n158,
    new_n159, new_n160, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n508, new_n509, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n647, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n138));
  INV_X1    g001(.A(G1gat), .ZN(new_n139));
  NAND3_X1  g002(.A1(new_n138), .A2(KEYINPUT16), .A3(new_n139), .ZN(new_n140));
  OAI21_X1  g003(.A(new_n140), .B1(new_n139), .B2(new_n138), .ZN(new_n141));
  XNOR2_X1  g004(.A(new_n141), .B(G8gat), .ZN(new_n142));
  INV_X1    g005(.A(KEYINPUT17), .ZN(new_n143));
  INV_X1    g006(.A(G29gat), .ZN(new_n144));
  INV_X1    g007(.A(G36gat), .ZN(new_n145));
  NAND3_X1  g008(.A1(new_n144), .A2(new_n145), .A3(KEYINPUT14), .ZN(new_n146));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n147));
  OAI21_X1  g010(.A(new_n147), .B1(G29gat), .B2(G36gat), .ZN(new_n148));
  NAND2_X1  g011(.A1(G29gat), .A2(G36gat), .ZN(new_n149));
  NAND3_X1  g012(.A1(new_n146), .A2(new_n148), .A3(new_n149), .ZN(new_n150));
  AND2_X1   g013(.A1(G43gat), .A2(G50gat), .ZN(new_n151));
  NOR2_X1   g014(.A1(G43gat), .A2(G50gat), .ZN(new_n152));
  NOR2_X1   g015(.A1(new_n151), .A2(new_n152), .ZN(new_n153));
  OAI21_X1  g016(.A(KEYINPUT15), .B1(new_n150), .B2(new_n153), .ZN(new_n154));
  AND2_X1   g017(.A1(G29gat), .A2(G36gat), .ZN(new_n155));
  NOR2_X1   g018(.A1(G29gat), .A2(G36gat), .ZN(new_n156));
  AOI21_X1  g019(.A(new_n155), .B1(KEYINPUT14), .B2(new_n156), .ZN(new_n157));
  INV_X1    g020(.A(KEYINPUT15), .ZN(new_n158));
  XNOR2_X1  g021(.A(G43gat), .B(G50gat), .ZN(new_n159));
  NAND4_X1  g022(.A1(new_n157), .A2(new_n158), .A3(new_n148), .A4(new_n159), .ZN(new_n160));
  AOI221_X4 g023(.A(new_n143), .B1(new_n150), .B2(new_n153), .C1(new_n154), .C2(new_n160), .ZN(new_n161));
  NAND2_X1  g024(.A1(new_n154), .A2(new_n160), .ZN(new_n162));
  NAND2_X1  g025(.A1(new_n150), .A2(new_n153), .ZN(new_n163));
  AOI21_X1  g026(.A(KEYINPUT17), .B1(new_n162), .B2(new_n163), .ZN(new_n164));
  OAI21_X1  g027(.A(new_n142), .B1(new_n161), .B2(new_n164), .ZN(new_n165));
  INV_X1    g028(.A(G8gat), .ZN(new_n166));
  XNOR2_X1  g029(.A(new_n141), .B(new_n166), .ZN(new_n167));
  NAND3_X1  g030(.A1(new_n167), .A2(new_n162), .A3(new_n163), .ZN(new_n168));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n169));
  NAND3_X1  g032(.A1(new_n165), .A2(new_n168), .A3(new_n169), .ZN(new_n170));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n171));
  NAND2_X1  g034(.A1(new_n170), .A2(new_n171), .ZN(new_n172));
  NAND2_X1  g035(.A1(new_n162), .A2(new_n163), .ZN(new_n173));
  NAND2_X1  g036(.A1(new_n142), .A2(new_n173), .ZN(new_n174));
  NAND2_X1  g037(.A1(new_n168), .A2(new_n174), .ZN(new_n175));
  XOR2_X1   g038(.A(new_n169), .B(KEYINPUT13), .Z(new_n176));
  NAND2_X1  g039(.A1(new_n175), .A2(new_n176), .ZN(new_n177));
  NAND4_X1  g040(.A1(new_n165), .A2(new_n168), .A3(KEYINPUT18), .A4(new_n169), .ZN(new_n178));
  NAND3_X1  g041(.A1(new_n172), .A2(new_n177), .A3(new_n178), .ZN(new_n179));
  XOR2_X1   g042(.A(G113gat), .B(G141gat), .Z(new_n180));
  XNOR2_X1  g043(.A(new_n180), .B(KEYINPUT11), .ZN(new_n181));
  XNOR2_X1  g044(.A(G169gat), .B(G197gat), .ZN(new_n182));
  XNOR2_X1  g045(.A(new_n181), .B(new_n182), .ZN(new_n183));
  XNOR2_X1  g046(.A(new_n183), .B(KEYINPUT12), .ZN(new_n184));
  XNOR2_X1  g047(.A(new_n179), .B(new_n184), .ZN(new_n185));
  INV_X1    g048(.A(KEYINPUT36), .ZN(new_n186));
  NAND2_X1  g049(.A1(G227gat), .A2(G233gat), .ZN(new_n187));
  NAND2_X1  g050(.A1(G183gat), .A2(G190gat), .ZN(new_n188));
  INV_X1    g051(.A(KEYINPUT24), .ZN(new_n189));
  NAND2_X1  g052(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  OR2_X1    g053(.A1(G183gat), .A2(G190gat), .ZN(new_n191));
  NAND3_X1  g054(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n192));
  NAND3_X1  g055(.A1(new_n190), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  INV_X1    g056(.A(KEYINPUT23), .ZN(new_n194));
  INV_X1    g057(.A(G169gat), .ZN(new_n195));
  INV_X1    g058(.A(G176gat), .ZN(new_n196));
  NAND3_X1  g059(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  OAI21_X1  g060(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n198));
  NAND2_X1  g061(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n200));
  NAND3_X1  g063(.A1(new_n193), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  INV_X1    g064(.A(KEYINPUT25), .ZN(new_n202));
  NAND2_X1  g065(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND4_X1  g066(.A1(new_n193), .A2(new_n199), .A3(KEYINPUT25), .A4(new_n200), .ZN(new_n204));
  NAND2_X1  g067(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XOR2_X1   g068(.A(G127gat), .B(G134gat), .Z(new_n206));
  XNOR2_X1  g069(.A(G113gat), .B(G120gat), .ZN(new_n207));
  OAI21_X1  g070(.A(new_n206), .B1(KEYINPUT1), .B2(new_n207), .ZN(new_n208));
  XOR2_X1   g071(.A(G113gat), .B(G120gat), .Z(new_n209));
  INV_X1    g072(.A(KEYINPUT1), .ZN(new_n210));
  XNOR2_X1  g073(.A(G127gat), .B(G134gat), .ZN(new_n211));
  NAND3_X1  g074(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g075(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g076(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n214));
  NAND2_X1  g077(.A1(new_n214), .A2(new_n200), .ZN(new_n215));
  NOR3_X1   g078(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n216));
  NOR2_X1   g079(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g080(.A(new_n217), .ZN(new_n218));
  XNOR2_X1  g081(.A(KEYINPUT27), .B(G183gat), .ZN(new_n219));
  INV_X1    g082(.A(G190gat), .ZN(new_n220));
  AOI21_X1  g083(.A(KEYINPUT28), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g084(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n222));
  NOR2_X1   g085(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n223));
  OAI211_X1 g086(.A(KEYINPUT28), .B(new_n220), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g087(.A(new_n224), .ZN(new_n225));
  OAI211_X1 g088(.A(new_n218), .B(new_n188), .C1(new_n221), .C2(new_n225), .ZN(new_n226));
  AND3_X1   g089(.A1(new_n205), .A2(new_n213), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g090(.A(new_n213), .B1(new_n205), .B2(new_n226), .ZN(new_n228));
  OAI21_X1  g091(.A(new_n187), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n230));
  NAND2_X1  g093(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g094(.A(KEYINPUT32), .B(new_n187), .C1(new_n227), .C2(new_n228), .ZN(new_n232));
  OR3_X1    g095(.A1(new_n227), .A2(new_n228), .A3(new_n187), .ZN(new_n233));
  NAND3_X1  g096(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g097(.A1(new_n234), .A2(KEYINPUT34), .ZN(new_n235));
  XNOR2_X1  g098(.A(G15gat), .B(G43gat), .ZN(new_n236));
  XNOR2_X1  g099(.A(G71gat), .B(G99gat), .ZN(new_n237));
  XOR2_X1   g100(.A(new_n236), .B(new_n237), .Z(new_n238));
  INV_X1    g101(.A(new_n238), .ZN(new_n239));
  INV_X1    g102(.A(KEYINPUT33), .ZN(new_n240));
  AOI21_X1  g103(.A(new_n239), .B1(new_n233), .B2(new_n240), .ZN(new_n241));
  INV_X1    g104(.A(KEYINPUT34), .ZN(new_n242));
  NAND4_X1  g105(.A1(new_n231), .A2(new_n233), .A3(new_n242), .A4(new_n232), .ZN(new_n243));
  AND3_X1   g106(.A1(new_n235), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g107(.A(new_n241), .B1(new_n235), .B2(new_n243), .ZN(new_n245));
  OAI21_X1  g108(.A(new_n186), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g109(.A1(new_n235), .A2(new_n243), .ZN(new_n247));
  INV_X1    g110(.A(new_n241), .ZN(new_n248));
  NAND2_X1  g111(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g112(.A1(new_n235), .A2(new_n241), .A3(new_n243), .ZN(new_n250));
  NAND3_X1  g113(.A1(new_n249), .A2(KEYINPUT36), .A3(new_n250), .ZN(new_n251));
  AND2_X1   g114(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g115(.A(G78gat), .B(G106gat), .ZN(new_n253));
  XNOR2_X1  g116(.A(new_n253), .B(KEYINPUT31), .ZN(new_n254));
  XOR2_X1   g117(.A(G22gat), .B(G50gat), .Z(new_n255));
  XNOR2_X1  g118(.A(G197gat), .B(G204gat), .ZN(new_n256));
  INV_X1    g119(.A(KEYINPUT22), .ZN(new_n257));
  INV_X1    g120(.A(G211gat), .ZN(new_n258));
  INV_X1    g121(.A(G218gat), .ZN(new_n259));
  OAI21_X1  g122(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g123(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g124(.A(G211gat), .B(G218gat), .ZN(new_n262));
  INV_X1    g125(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g126(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g127(.A1(new_n262), .A2(new_n256), .A3(new_n260), .ZN(new_n265));
  NAND2_X1  g128(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n267));
  NAND2_X1  g130(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XOR2_X1   g131(.A(G155gat), .B(G162gat), .Z(new_n269));
  INV_X1    g132(.A(G141gat), .ZN(new_n270));
  INV_X1    g133(.A(G148gat), .ZN(new_n271));
  NAND2_X1  g134(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g135(.A1(G141gat), .A2(G148gat), .ZN(new_n273));
  NAND2_X1  g136(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g137(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g138(.A(G155gat), .B(G162gat), .ZN(new_n276));
  NOR2_X1   g139(.A1(new_n276), .A2(KEYINPUT2), .ZN(new_n277));
  INV_X1    g140(.A(G155gat), .ZN(new_n278));
  INV_X1    g141(.A(G162gat), .ZN(new_n279));
  NAND3_X1  g142(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT2), .ZN(new_n280));
  NAND3_X1  g143(.A1(new_n280), .A2(new_n272), .A3(new_n273), .ZN(new_n281));
  OAI21_X1  g144(.A(new_n275), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g145(.A1(new_n282), .A2(KEYINPUT3), .ZN(new_n283));
  AND2_X1   g146(.A1(new_n272), .A2(new_n273), .ZN(new_n284));
  OAI211_X1 g147(.A(new_n284), .B(new_n280), .C1(KEYINPUT2), .C2(new_n276), .ZN(new_n285));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n286));
  NAND3_X1  g149(.A1(new_n285), .A2(new_n286), .A3(new_n275), .ZN(new_n287));
  NAND3_X1  g150(.A1(new_n264), .A2(KEYINPUT29), .A3(new_n265), .ZN(new_n288));
  NAND4_X1  g151(.A1(new_n268), .A2(new_n283), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g152(.A1(G228gat), .A2(G233gat), .ZN(new_n290));
  INV_X1    g153(.A(KEYINPUT2), .ZN(new_n291));
  NAND2_X1  g154(.A1(new_n269), .A2(new_n291), .ZN(new_n292));
  INV_X1    g155(.A(new_n281), .ZN(new_n293));
  AOI22_X1  g156(.A1(new_n292), .A2(new_n293), .B1(new_n269), .B2(new_n274), .ZN(new_n294));
  NAND2_X1  g157(.A1(new_n294), .A2(new_n266), .ZN(new_n295));
  NAND3_X1  g158(.A1(new_n289), .A2(new_n290), .A3(new_n295), .ZN(new_n296));
  INV_X1    g159(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g160(.A(new_n290), .B1(new_n289), .B2(new_n295), .ZN(new_n298));
  OAI21_X1  g161(.A(new_n255), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g162(.A1(new_n289), .A2(new_n295), .ZN(new_n300));
  INV_X1    g163(.A(new_n290), .ZN(new_n301));
  NAND2_X1  g164(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g165(.A(new_n255), .ZN(new_n303));
  NAND3_X1  g166(.A1(new_n302), .A2(new_n296), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g167(.A(new_n254), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  INV_X1    g168(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g169(.A1(new_n299), .A2(new_n304), .A3(new_n254), .ZN(new_n307));
  NAND2_X1  g170(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g171(.A1(new_n283), .A2(new_n213), .A3(new_n287), .ZN(new_n309));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n310));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n311));
  OAI21_X1  g174(.A(new_n311), .B1(new_n213), .B2(new_n282), .ZN(new_n312));
  AND2_X1   g175(.A1(new_n208), .A2(new_n212), .ZN(new_n313));
  NAND3_X1  g176(.A1(new_n313), .A2(KEYINPUT4), .A3(new_n294), .ZN(new_n314));
  NAND4_X1  g177(.A1(new_n309), .A2(new_n310), .A3(new_n312), .A4(new_n314), .ZN(new_n315));
  XNOR2_X1  g178(.A(new_n315), .B(KEYINPUT5), .ZN(new_n316));
  INV_X1    g179(.A(KEYINPUT6), .ZN(new_n317));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n318));
  XNOR2_X1  g181(.A(new_n318), .B(KEYINPUT0), .ZN(new_n319));
  XNOR2_X1  g182(.A(G57gat), .B(G85gat), .ZN(new_n320));
  XNOR2_X1  g183(.A(new_n319), .B(new_n320), .ZN(new_n321));
  XNOR2_X1  g184(.A(new_n294), .B(new_n213), .ZN(new_n322));
  OR2_X1    g185(.A1(new_n322), .A2(new_n310), .ZN(new_n323));
  NAND4_X1  g186(.A1(new_n316), .A2(new_n317), .A3(new_n321), .A4(new_n323), .ZN(new_n324));
  AND2_X1   g187(.A1(new_n314), .A2(new_n312), .ZN(new_n325));
  NAND4_X1  g188(.A1(new_n325), .A2(KEYINPUT5), .A3(new_n310), .A4(new_n309), .ZN(new_n326));
  INV_X1    g189(.A(KEYINPUT5), .ZN(new_n327));
  NAND2_X1  g190(.A1(new_n315), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g191(.A1(new_n326), .A2(new_n328), .A3(new_n323), .A4(new_n321), .ZN(new_n329));
  NAND2_X1  g192(.A1(new_n329), .A2(KEYINPUT6), .ZN(new_n330));
  NAND3_X1  g193(.A1(new_n326), .A2(new_n328), .A3(new_n323), .ZN(new_n331));
  INV_X1    g194(.A(new_n321), .ZN(new_n332));
  NAND2_X1  g195(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g196(.A1(new_n324), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  AND3_X1   g197(.A1(new_n205), .A2(new_n226), .A3(new_n266), .ZN(new_n335));
  AOI21_X1  g198(.A(new_n266), .B1(new_n205), .B2(new_n226), .ZN(new_n336));
  OAI211_X1 g199(.A(G226gat), .B(G233gat), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND3_X1  g200(.A1(new_n205), .A2(new_n226), .A3(new_n266), .ZN(new_n338));
  NAND2_X1  g201(.A1(G226gat), .A2(G233gat), .ZN(new_n339));
  NAND2_X1  g202(.A1(new_n219), .A2(new_n220), .ZN(new_n340));
  INV_X1    g203(.A(KEYINPUT28), .ZN(new_n341));
  NAND2_X1  g204(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g205(.A(new_n217), .B1(new_n342), .B2(new_n224), .ZN(new_n343));
  AOI22_X1  g206(.A1(new_n343), .A2(new_n188), .B1(new_n203), .B2(new_n204), .ZN(new_n344));
  NAND2_X1  g207(.A1(new_n268), .A2(new_n288), .ZN(new_n345));
  OAI211_X1 g208(.A(new_n338), .B(new_n339), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  XNOR2_X1  g209(.A(G8gat), .B(G36gat), .ZN(new_n347));
  XNOR2_X1  g210(.A(G64gat), .B(G92gat), .ZN(new_n348));
  XNOR2_X1  g211(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g212(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g213(.A1(new_n337), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  INV_X1    g214(.A(KEYINPUT37), .ZN(new_n352));
  INV_X1    g215(.A(new_n346), .ZN(new_n353));
  NAND2_X1  g216(.A1(new_n205), .A2(new_n226), .ZN(new_n354));
  INV_X1    g217(.A(new_n266), .ZN(new_n355));
  NAND2_X1  g218(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g219(.A(new_n339), .B1(new_n356), .B2(new_n338), .ZN(new_n357));
  OAI21_X1  g220(.A(new_n352), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g221(.A1(new_n337), .A2(KEYINPUT37), .A3(new_n346), .ZN(new_n359));
  NAND2_X1  g222(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g223(.A(KEYINPUT38), .B1(new_n360), .B2(new_n349), .ZN(new_n361));
  INV_X1    g224(.A(KEYINPUT38), .ZN(new_n362));
  AOI211_X1 g225(.A(new_n362), .B(new_n350), .C1(new_n358), .C2(new_n359), .ZN(new_n363));
  OAI211_X1 g226(.A(new_n334), .B(new_n351), .C1(new_n361), .C2(new_n363), .ZN(new_n364));
  AOI21_X1  g227(.A(new_n350), .B1(new_n337), .B2(new_n346), .ZN(new_n365));
  INV_X1    g228(.A(new_n351), .ZN(new_n366));
  AOI21_X1  g229(.A(new_n365), .B1(new_n366), .B2(KEYINPUT30), .ZN(new_n367));
  INV_X1    g230(.A(KEYINPUT30), .ZN(new_n368));
  NAND2_X1  g231(.A1(new_n351), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g232(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g233(.A1(new_n309), .A2(new_n312), .A3(new_n314), .ZN(new_n371));
  INV_X1    g234(.A(new_n310), .ZN(new_n372));
  NAND2_X1  g235(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g236(.A(KEYINPUT39), .ZN(new_n374));
  NAND2_X1  g237(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g238(.A1(new_n322), .A2(new_n310), .ZN(new_n376));
  NAND3_X1  g239(.A1(new_n371), .A2(KEYINPUT39), .A3(new_n372), .ZN(new_n377));
  NAND3_X1  g240(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g241(.A1(new_n378), .A2(new_n332), .ZN(new_n379));
  INV_X1    g242(.A(KEYINPUT40), .ZN(new_n380));
  NAND2_X1  g243(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g244(.A1(new_n378), .A2(KEYINPUT40), .A3(new_n332), .ZN(new_n382));
  NAND4_X1  g245(.A1(new_n370), .A2(new_n381), .A3(new_n329), .A4(new_n382), .ZN(new_n383));
  AOI21_X1  g246(.A(new_n308), .B1(new_n364), .B2(new_n383), .ZN(new_n384));
  INV_X1    g247(.A(new_n307), .ZN(new_n385));
  NOR2_X1   g248(.A1(new_n385), .A2(new_n305), .ZN(new_n386));
  NOR3_X1   g249(.A1(new_n386), .A2(new_n334), .A3(new_n370), .ZN(new_n387));
  OAI21_X1  g250(.A(new_n252), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  AND2_X1   g251(.A1(new_n367), .A2(new_n369), .ZN(new_n389));
  OAI21_X1  g252(.A(new_n389), .B1(new_n244), .B2(new_n245), .ZN(new_n390));
  INV_X1    g253(.A(new_n334), .ZN(new_n391));
  NAND2_X1  g254(.A1(new_n391), .A2(new_n386), .ZN(new_n392));
  OAI21_X1  g255(.A(KEYINPUT35), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g256(.A1(new_n308), .A2(new_n334), .ZN(new_n394));
  NAND2_X1  g257(.A1(new_n249), .A2(new_n250), .ZN(new_n395));
  INV_X1    g258(.A(KEYINPUT35), .ZN(new_n396));
  NAND4_X1  g259(.A1(new_n394), .A2(new_n395), .A3(new_n396), .A4(new_n389), .ZN(new_n397));
  NAND2_X1  g260(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g261(.A(new_n185), .B1(new_n388), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g262(.A1(new_n173), .A2(new_n143), .ZN(new_n400));
  NAND3_X1  g263(.A1(new_n162), .A2(KEYINPUT17), .A3(new_n163), .ZN(new_n401));
  NAND2_X1  g264(.A1(G85gat), .A2(G92gat), .ZN(new_n402));
  NAND2_X1  g265(.A1(new_n402), .A2(KEYINPUT7), .ZN(new_n403));
  INV_X1    g266(.A(KEYINPUT7), .ZN(new_n404));
  NAND3_X1  g267(.A1(new_n404), .A2(G85gat), .A3(G92gat), .ZN(new_n405));
  NAND2_X1  g268(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  OR2_X1    g269(.A1(G85gat), .A2(G92gat), .ZN(new_n407));
  NAND2_X1  g270(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g271(.A(G99gat), .ZN(new_n409));
  INV_X1    g272(.A(G106gat), .ZN(new_n410));
  NAND2_X1  g273(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g274(.A1(G99gat), .A2(G106gat), .ZN(new_n412));
  NAND2_X1  g275(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g276(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g277(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  INV_X1    g278(.A(KEYINPUT8), .ZN(new_n416));
  NAND3_X1  g279(.A1(new_n411), .A2(new_n416), .A3(new_n412), .ZN(new_n417));
  NAND3_X1  g280(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT8), .ZN(new_n418));
  NAND4_X1  g281(.A1(new_n406), .A2(new_n417), .A3(new_n407), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g282(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g283(.A1(new_n400), .A2(new_n401), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g284(.A1(G232gat), .A2(G233gat), .ZN(new_n422));
  INV_X1    g285(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g286(.A(new_n420), .B1(new_n162), .B2(new_n163), .ZN(new_n424));
  INV_X1    g287(.A(new_n424), .ZN(new_n425));
  AND3_X1   g288(.A1(new_n421), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  INV_X1    g289(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g290(.A1(new_n421), .A2(new_n425), .ZN(new_n428));
  AOI21_X1  g291(.A(KEYINPUT41), .B1(new_n428), .B2(new_n422), .ZN(new_n429));
  INV_X1    g292(.A(KEYINPUT41), .ZN(new_n430));
  AOI211_X1 g293(.A(new_n430), .B(new_n423), .C1(new_n421), .C2(new_n425), .ZN(new_n431));
  OAI21_X1  g294(.A(new_n427), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  XOR2_X1   g295(.A(G134gat), .B(G162gat), .Z(new_n433));
  NAND2_X1  g296(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g297(.A1(new_n161), .A2(new_n164), .ZN(new_n435));
  AOI21_X1  g298(.A(new_n424), .B1(new_n435), .B2(new_n420), .ZN(new_n436));
  OAI21_X1  g299(.A(new_n430), .B1(new_n436), .B2(new_n423), .ZN(new_n437));
  NAND3_X1  g300(.A1(new_n428), .A2(KEYINPUT41), .A3(new_n422), .ZN(new_n438));
  NAND2_X1  g301(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g302(.A(new_n433), .ZN(new_n440));
  NAND3_X1  g303(.A1(new_n439), .A2(new_n427), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g304(.A(G190gat), .B(G218gat), .ZN(new_n442));
  AND3_X1   g305(.A1(new_n434), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g306(.A(new_n442), .B1(new_n434), .B2(new_n441), .ZN(new_n444));
  NOR2_X1   g307(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  XOR2_X1   g308(.A(G57gat), .B(G64gat), .Z(new_n446));
  INV_X1    g309(.A(G71gat), .ZN(new_n447));
  INV_X1    g310(.A(G78gat), .ZN(new_n448));
  NAND2_X1  g311(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g312(.A1(G71gat), .A2(G78gat), .ZN(new_n450));
  NAND3_X1  g313(.A1(new_n449), .A2(KEYINPUT9), .A3(new_n450), .ZN(new_n451));
  OR3_X1    g314(.A1(KEYINPUT9), .A2(G71gat), .A3(G78gat), .ZN(new_n452));
  NAND3_X1  g315(.A1(new_n446), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  XNOR2_X1  g316(.A(G57gat), .B(G64gat), .ZN(new_n454));
  NAND3_X1  g317(.A1(new_n454), .A2(new_n449), .A3(new_n450), .ZN(new_n455));
  NAND2_X1  g318(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g319(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g320(.A(new_n457), .B1(new_n167), .B2(KEYINPUT21), .ZN(new_n458));
  XNOR2_X1  g321(.A(G127gat), .B(G155gat), .ZN(new_n459));
  XOR2_X1   g322(.A(new_n459), .B(KEYINPUT19), .Z(new_n460));
  XNOR2_X1  g323(.A(G183gat), .B(G211gat), .ZN(new_n461));
  XNOR2_X1  g324(.A(new_n461), .B(KEYINPUT20), .ZN(new_n462));
  XNOR2_X1  g325(.A(new_n460), .B(new_n462), .ZN(new_n463));
  XNOR2_X1  g326(.A(new_n458), .B(new_n463), .ZN(new_n464));
  NOR2_X1   g327(.A1(new_n167), .A2(KEYINPUT21), .ZN(new_n465));
  NAND2_X1  g328(.A1(G231gat), .A2(G233gat), .ZN(new_n466));
  XNOR2_X1  g329(.A(new_n465), .B(new_n466), .ZN(new_n467));
  XOR2_X1   g330(.A(new_n464), .B(new_n467), .Z(new_n468));
  INV_X1    g331(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g332(.A1(new_n445), .A2(new_n469), .ZN(new_n470));
  AND4_X1   g333(.A1(new_n407), .A2(new_n406), .A3(new_n417), .A4(new_n418), .ZN(new_n471));
  AOI21_X1  g334(.A(new_n413), .B1(new_n406), .B2(new_n407), .ZN(new_n472));
  OAI21_X1  g335(.A(new_n456), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g336(.A(KEYINPUT10), .ZN(new_n474));
  NAND4_X1  g337(.A1(new_n415), .A2(new_n455), .A3(new_n419), .A4(new_n453), .ZN(new_n475));
  NAND3_X1  g338(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NOR2_X1   g339(.A1(new_n471), .A2(new_n472), .ZN(new_n477));
  NAND3_X1  g340(.A1(new_n477), .A2(KEYINPUT10), .A3(new_n457), .ZN(new_n478));
  NAND2_X1  g341(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g342(.A1(G230gat), .A2(G233gat), .ZN(new_n480));
  NAND2_X1  g343(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g344(.A1(new_n473), .A2(new_n475), .ZN(new_n482));
  INV_X1    g345(.A(new_n480), .ZN(new_n483));
  NAND2_X1  g346(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g347(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g348(.A(G120gat), .B(G148gat), .ZN(new_n486));
  XNOR2_X1  g349(.A(G176gat), .B(G204gat), .ZN(new_n487));
  XNOR2_X1  g350(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND2_X1  g351(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g352(.A(new_n488), .ZN(new_n490));
  NAND3_X1  g353(.A1(new_n481), .A2(new_n484), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g354(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g355(.A1(new_n470), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g356(.A1(new_n399), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g357(.A1(new_n494), .A2(new_n391), .ZN(new_n495));
  XNOR2_X1  g358(.A(new_n495), .B(new_n139), .ZN(G1324gat));
  INV_X1    g359(.A(new_n494), .ZN(new_n497));
  NAND2_X1  g360(.A1(new_n497), .A2(new_n370), .ZN(new_n498));
  XNOR2_X1  g361(.A(KEYINPUT16), .B(G8gat), .ZN(new_n499));
  NOR2_X1   g362(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OR2_X1    g363(.A1(new_n500), .A2(KEYINPUT42), .ZN(new_n501));
  NAND2_X1  g364(.A1(new_n498), .A2(G8gat), .ZN(new_n502));
  NAND2_X1  g365(.A1(new_n500), .A2(KEYINPUT42), .ZN(new_n503));
  NAND3_X1  g366(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(G1325gat));
  OAI21_X1  g367(.A(G15gat), .B1(new_n494), .B2(new_n252), .ZN(new_n505));
  NAND2_X1  g368(.A1(new_n497), .A2(new_n395), .ZN(new_n506));
  OAI21_X1  g369(.A(new_n505), .B1(new_n506), .B2(G15gat), .ZN(G1326gat));
  NOR2_X1   g370(.A1(new_n494), .A2(new_n386), .ZN(new_n508));
  XOR2_X1   g371(.A(KEYINPUT43), .B(G22gat), .Z(new_n509));
  XNOR2_X1  g372(.A(new_n508), .B(new_n509), .ZN(G1327gat));
  INV_X1    g373(.A(new_n492), .ZN(new_n511));
  NOR2_X1   g374(.A1(new_n445), .A2(new_n469), .ZN(new_n512));
  NAND3_X1  g375(.A1(new_n399), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NOR3_X1   g376(.A1(new_n513), .A2(G29gat), .A3(new_n391), .ZN(new_n514));
  XOR2_X1   g377(.A(new_n514), .B(KEYINPUT45), .Z(new_n515));
  INV_X1    g378(.A(KEYINPUT44), .ZN(new_n516));
  NAND2_X1  g379(.A1(new_n388), .A2(new_n398), .ZN(new_n517));
  INV_X1    g380(.A(new_n442), .ZN(new_n518));
  AOI21_X1  g381(.A(new_n440), .B1(new_n439), .B2(new_n427), .ZN(new_n519));
  AOI211_X1 g382(.A(new_n426), .B(new_n433), .C1(new_n437), .C2(new_n438), .ZN(new_n520));
  OAI21_X1  g383(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g384(.A1(new_n434), .A2(new_n441), .A3(new_n442), .ZN(new_n522));
  NAND2_X1  g385(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g386(.A(new_n516), .B1(new_n517), .B2(new_n523), .ZN(new_n524));
  AOI211_X1 g387(.A(KEYINPUT44), .B(new_n445), .C1(new_n388), .C2(new_n398), .ZN(new_n525));
  OAI211_X1 g388(.A(new_n511), .B(new_n468), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NOR3_X1   g389(.A1(new_n526), .A2(new_n391), .A3(new_n185), .ZN(new_n527));
  OAI21_X1  g390(.A(new_n515), .B1(new_n144), .B2(new_n527), .ZN(G1328gat));
  NOR3_X1   g391(.A1(new_n513), .A2(G36gat), .A3(new_n389), .ZN(new_n529));
  XNOR2_X1  g392(.A(new_n529), .B(KEYINPUT46), .ZN(new_n530));
  NOR3_X1   g393(.A1(new_n526), .A2(new_n185), .A3(new_n389), .ZN(new_n531));
  OAI21_X1  g394(.A(new_n530), .B1(new_n145), .B2(new_n531), .ZN(G1329gat));
  INV_X1    g395(.A(G43gat), .ZN(new_n533));
  NOR4_X1   g396(.A1(new_n526), .A2(new_n533), .A3(new_n185), .A4(new_n252), .ZN(new_n534));
  INV_X1    g397(.A(new_n395), .ZN(new_n535));
  OAI21_X1  g398(.A(new_n533), .B1(new_n513), .B2(new_n535), .ZN(new_n536));
  INV_X1    g399(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g400(.A(KEYINPUT47), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  INV_X1    g401(.A(KEYINPUT47), .ZN(new_n539));
  INV_X1    g402(.A(new_n387), .ZN(new_n540));
  AND3_X1   g403(.A1(new_n337), .A2(KEYINPUT37), .A3(new_n346), .ZN(new_n541));
  AOI21_X1  g404(.A(KEYINPUT37), .B1(new_n337), .B2(new_n346), .ZN(new_n542));
  OAI21_X1  g405(.A(new_n349), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g406(.A1(new_n543), .A2(new_n362), .ZN(new_n544));
  NAND3_X1  g407(.A1(new_n360), .A2(KEYINPUT38), .A3(new_n349), .ZN(new_n545));
  AOI21_X1  g408(.A(new_n366), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g409(.A1(new_n367), .A2(new_n369), .B1(new_n379), .B2(new_n380), .ZN(new_n547));
  AND2_X1   g410(.A1(new_n382), .A2(new_n329), .ZN(new_n548));
  AOI22_X1  g411(.A1(new_n546), .A2(new_n334), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g412(.A(new_n540), .B1(new_n549), .B2(new_n308), .ZN(new_n550));
  AOI22_X1  g413(.A1(new_n550), .A2(new_n252), .B1(new_n393), .B2(new_n397), .ZN(new_n551));
  OAI21_X1  g414(.A(KEYINPUT44), .B1(new_n551), .B2(new_n445), .ZN(new_n552));
  NAND3_X1  g415(.A1(new_n517), .A2(new_n516), .A3(new_n523), .ZN(new_n553));
  AOI21_X1  g416(.A(new_n469), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g417(.A(new_n185), .ZN(new_n555));
  INV_X1    g418(.A(new_n252), .ZN(new_n556));
  NAND4_X1  g419(.A1(new_n554), .A2(new_n555), .A3(new_n556), .A4(new_n511), .ZN(new_n557));
  OAI211_X1 g420(.A(new_n539), .B(new_n536), .C1(new_n557), .C2(new_n533), .ZN(new_n558));
  NAND2_X1  g421(.A1(new_n538), .A2(new_n558), .ZN(G1330gat));
  INV_X1    g422(.A(G50gat), .ZN(new_n560));
  NOR4_X1   g423(.A1(new_n526), .A2(new_n560), .A3(new_n185), .A4(new_n386), .ZN(new_n561));
  OAI21_X1  g424(.A(new_n560), .B1(new_n513), .B2(new_n386), .ZN(new_n562));
  INV_X1    g425(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g426(.A(KEYINPUT48), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  INV_X1    g427(.A(KEYINPUT48), .ZN(new_n565));
  NAND4_X1  g428(.A1(new_n554), .A2(new_n555), .A3(new_n308), .A4(new_n511), .ZN(new_n566));
  OAI211_X1 g429(.A(new_n565), .B(new_n562), .C1(new_n566), .C2(new_n560), .ZN(new_n567));
  NAND2_X1  g430(.A1(new_n564), .A2(new_n567), .ZN(G1331gat));
  NOR4_X1   g431(.A1(new_n551), .A2(new_n555), .A3(new_n511), .A4(new_n470), .ZN(new_n569));
  NAND2_X1  g432(.A1(new_n569), .A2(new_n334), .ZN(new_n570));
  XNOR2_X1  g433(.A(new_n570), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g434(.A(new_n555), .B1(new_n388), .B2(new_n398), .ZN(new_n572));
  NAND4_X1  g435(.A1(new_n572), .A2(new_n492), .A3(new_n469), .A4(new_n445), .ZN(new_n573));
  AOI211_X1 g436(.A(new_n389), .B(new_n573), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n574));
  NOR2_X1   g437(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n575));
  XNOR2_X1  g438(.A(new_n574), .B(new_n575), .ZN(G1333gat));
  AOI21_X1  g439(.A(new_n447), .B1(new_n569), .B2(new_n556), .ZN(new_n577));
  NOR3_X1   g440(.A1(new_n573), .A2(G71gat), .A3(new_n535), .ZN(new_n578));
  NOR2_X1   g441(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g442(.A(new_n579), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g443(.A1(new_n573), .A2(new_n386), .ZN(new_n581));
  XNOR2_X1  g444(.A(new_n581), .B(new_n448), .ZN(G1335gat));
  NAND3_X1  g445(.A1(new_n517), .A2(new_n185), .A3(new_n512), .ZN(new_n583));
  INV_X1    g446(.A(KEYINPUT51), .ZN(new_n584));
  NAND2_X1  g447(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g448(.A1(new_n572), .A2(KEYINPUT51), .A3(new_n512), .ZN(new_n586));
  AOI21_X1  g449(.A(new_n511), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g450(.A(G85gat), .B1(new_n587), .B2(new_n334), .ZN(new_n588));
  OAI211_X1 g451(.A(new_n185), .B(new_n468), .C1(new_n524), .C2(new_n525), .ZN(new_n589));
  NOR3_X1   g452(.A1(new_n589), .A2(new_n391), .A3(new_n511), .ZN(new_n590));
  AOI21_X1  g453(.A(new_n588), .B1(G85gat), .B2(new_n590), .ZN(G1336gat));
  INV_X1    g454(.A(KEYINPUT52), .ZN(new_n592));
  INV_X1    g455(.A(G92gat), .ZN(new_n593));
  NOR4_X1   g456(.A1(new_n589), .A2(new_n593), .A3(new_n389), .A4(new_n511), .ZN(new_n594));
  AOI21_X1  g457(.A(G92gat), .B1(new_n587), .B2(new_n370), .ZN(new_n595));
  OAI21_X1  g458(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g459(.A1(new_n583), .A2(new_n584), .ZN(new_n597));
  AOI21_X1  g460(.A(KEYINPUT51), .B1(new_n572), .B2(new_n512), .ZN(new_n598));
  OAI211_X1 g461(.A(new_n370), .B(new_n492), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  NAND2_X1  g462(.A1(new_n599), .A2(new_n593), .ZN(new_n600));
  NAND4_X1  g463(.A1(new_n554), .A2(new_n185), .A3(new_n370), .A4(new_n492), .ZN(new_n601));
  OAI211_X1 g464(.A(new_n600), .B(KEYINPUT52), .C1(new_n593), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g465(.A1(new_n596), .A2(new_n602), .ZN(G1337gat));
  AOI21_X1  g466(.A(G99gat), .B1(new_n587), .B2(new_n395), .ZN(new_n604));
  NOR3_X1   g467(.A1(new_n589), .A2(new_n252), .A3(new_n511), .ZN(new_n605));
  AOI21_X1  g468(.A(new_n604), .B1(G99gat), .B2(new_n605), .ZN(G1338gat));
  INV_X1    g469(.A(KEYINPUT53), .ZN(new_n607));
  NOR4_X1   g470(.A1(new_n589), .A2(new_n410), .A3(new_n386), .A4(new_n511), .ZN(new_n608));
  AOI21_X1  g471(.A(G106gat), .B1(new_n587), .B2(new_n308), .ZN(new_n609));
  OAI21_X1  g472(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI211_X1 g473(.A(new_n308), .B(new_n492), .C1(new_n597), .C2(new_n598), .ZN(new_n611));
  NAND2_X1  g474(.A1(new_n611), .A2(new_n410), .ZN(new_n612));
  NAND4_X1  g475(.A1(new_n554), .A2(new_n185), .A3(new_n308), .A4(new_n492), .ZN(new_n613));
  OAI211_X1 g476(.A(new_n612), .B(KEYINPUT53), .C1(new_n410), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g477(.A1(new_n610), .A2(new_n614), .ZN(G1339gat));
  NOR4_X1   g478(.A1(new_n523), .A2(new_n555), .A3(new_n492), .A4(new_n468), .ZN(new_n616));
  NAND4_X1  g479(.A1(new_n172), .A2(new_n177), .A3(new_n178), .A4(new_n184), .ZN(new_n617));
  NOR2_X1   g480(.A1(new_n175), .A2(new_n176), .ZN(new_n618));
  AOI21_X1  g481(.A(new_n169), .B1(new_n165), .B2(new_n168), .ZN(new_n619));
  OAI21_X1  g482(.A(new_n183), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g483(.A(KEYINPUT54), .B1(new_n479), .B2(new_n480), .ZN(new_n621));
  INV_X1    g484(.A(KEYINPUT54), .ZN(new_n622));
  AOI211_X1 g485(.A(new_n622), .B(new_n483), .C1(new_n476), .C2(new_n478), .ZN(new_n623));
  NAND3_X1  g486(.A1(new_n476), .A2(new_n483), .A3(new_n478), .ZN(new_n624));
  INV_X1    g487(.A(new_n624), .ZN(new_n625));
  NOR3_X1   g488(.A1(new_n621), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  NOR3_X1   g489(.A1(new_n626), .A2(KEYINPUT55), .A3(new_n490), .ZN(new_n627));
  INV_X1    g490(.A(KEYINPUT55), .ZN(new_n628));
  NAND2_X1  g491(.A1(new_n481), .A2(new_n622), .ZN(new_n629));
  NAND3_X1  g492(.A1(new_n479), .A2(KEYINPUT54), .A3(new_n480), .ZN(new_n630));
  NAND3_X1  g493(.A1(new_n629), .A2(new_n624), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g494(.A(new_n628), .B1(new_n631), .B2(new_n488), .ZN(new_n632));
  OAI21_X1  g495(.A(new_n491), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  INV_X1    g496(.A(new_n633), .ZN(new_n634));
  NAND4_X1  g497(.A1(new_n523), .A2(new_n617), .A3(new_n620), .A4(new_n634), .ZN(new_n635));
  NAND3_X1  g498(.A1(new_n492), .A2(new_n617), .A3(new_n620), .ZN(new_n636));
  OAI21_X1  g499(.A(new_n636), .B1(new_n633), .B2(new_n185), .ZN(new_n637));
  NAND2_X1  g500(.A1(new_n445), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g501(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g502(.A(new_n616), .B1(new_n639), .B2(new_n468), .ZN(new_n640));
  NOR2_X1   g503(.A1(new_n640), .A2(new_n535), .ZN(new_n641));
  NAND4_X1  g504(.A1(new_n641), .A2(new_n334), .A3(new_n389), .A4(new_n386), .ZN(new_n642));
  NOR2_X1   g505(.A1(new_n642), .A2(new_n185), .ZN(new_n643));
  XOR2_X1   g506(.A(new_n643), .B(G113gat), .Z(G1340gat));
  NOR2_X1   g507(.A1(new_n642), .A2(new_n511), .ZN(new_n645));
  XOR2_X1   g508(.A(new_n645), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g509(.A1(new_n642), .A2(new_n468), .ZN(new_n647));
  XOR2_X1   g510(.A(new_n647), .B(G127gat), .Z(G1342gat));
  AND2_X1   g511(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n649));
  NOR3_X1   g512(.A1(new_n642), .A2(new_n445), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g513(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n651));
  XNOR2_X1  g514(.A(new_n650), .B(new_n651), .ZN(G1343gat));
  INV_X1    g515(.A(KEYINPUT57), .ZN(new_n653));
  OAI21_X1  g516(.A(new_n653), .B1(new_n640), .B2(new_n386), .ZN(new_n654));
  AOI21_X1  g517(.A(new_n469), .B1(new_n635), .B2(new_n638), .ZN(new_n655));
  OAI211_X1 g518(.A(KEYINPUT57), .B(new_n308), .C1(new_n655), .C2(new_n616), .ZN(new_n656));
  AOI21_X1  g519(.A(new_n556), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g520(.A1(new_n391), .A2(new_n370), .ZN(new_n658));
  NAND4_X1  g521(.A1(new_n657), .A2(G141gat), .A3(new_n555), .A4(new_n658), .ZN(new_n659));
  NOR2_X1   g522(.A1(new_n640), .A2(new_n386), .ZN(new_n660));
  NAND4_X1  g523(.A1(new_n660), .A2(new_n555), .A3(new_n252), .A4(new_n658), .ZN(new_n661));
  NAND2_X1  g524(.A1(new_n661), .A2(new_n270), .ZN(new_n662));
  NAND2_X1  g525(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g526(.A(KEYINPUT58), .ZN(new_n664));
  NAND2_X1  g527(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g528(.A1(new_n659), .A2(KEYINPUT58), .A3(new_n662), .ZN(new_n666));
  NAND2_X1  g529(.A1(new_n665), .A2(new_n666), .ZN(G1344gat));
  NAND2_X1  g530(.A1(new_n654), .A2(new_n656), .ZN(new_n668));
  NAND4_X1  g531(.A1(new_n668), .A2(new_n252), .A3(new_n492), .A4(new_n658), .ZN(new_n669));
  INV_X1    g532(.A(KEYINPUT59), .ZN(new_n670));
  AND3_X1   g533(.A1(new_n669), .A2(new_n670), .A3(G148gat), .ZN(new_n671));
  AOI21_X1  g534(.A(new_n670), .B1(new_n669), .B2(G148gat), .ZN(new_n672));
  NAND2_X1  g535(.A1(new_n660), .A2(new_n252), .ZN(new_n673));
  INV_X1    g536(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g537(.A1(new_n674), .A2(new_n658), .ZN(new_n675));
  NAND2_X1  g538(.A1(new_n492), .A2(new_n271), .ZN(new_n676));
  OAI22_X1  g539(.A1(new_n671), .A2(new_n672), .B1(new_n675), .B2(new_n676), .ZN(G1345gat));
  OAI21_X1  g540(.A(new_n278), .B1(new_n675), .B2(new_n468), .ZN(new_n678));
  NAND4_X1  g541(.A1(new_n657), .A2(G155gat), .A3(new_n469), .A4(new_n658), .ZN(new_n679));
  AND2_X1   g542(.A1(new_n678), .A2(new_n679), .ZN(G1346gat));
  OAI21_X1  g543(.A(new_n279), .B1(new_n675), .B2(new_n445), .ZN(new_n681));
  NAND4_X1  g544(.A1(new_n657), .A2(G162gat), .A3(new_n523), .A4(new_n658), .ZN(new_n682));
  AND2_X1   g545(.A1(new_n681), .A2(new_n682), .ZN(G1347gat));
  NOR2_X1   g546(.A1(new_n392), .A2(new_n389), .ZN(new_n684));
  NAND2_X1  g547(.A1(new_n641), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g548(.A1(new_n685), .A2(new_n185), .ZN(new_n686));
  XNOR2_X1  g549(.A(new_n686), .B(new_n195), .ZN(G1348gat));
  NOR2_X1   g550(.A1(new_n685), .A2(new_n511), .ZN(new_n688));
  XNOR2_X1  g551(.A(new_n688), .B(new_n196), .ZN(G1349gat));
  INV_X1    g552(.A(new_n685), .ZN(new_n690));
  NAND3_X1  g553(.A1(new_n690), .A2(new_n219), .A3(new_n469), .ZN(new_n691));
  OAI21_X1  g554(.A(G183gat), .B1(new_n685), .B2(new_n468), .ZN(new_n692));
  NAND2_X1  g555(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g556(.A1(new_n693), .A2(KEYINPUT60), .ZN(new_n694));
  INV_X1    g557(.A(KEYINPUT60), .ZN(new_n695));
  NAND3_X1  g558(.A1(new_n691), .A2(new_n695), .A3(new_n692), .ZN(new_n696));
  NAND2_X1  g559(.A1(new_n694), .A2(new_n696), .ZN(G1350gat));
  NAND2_X1  g560(.A1(new_n690), .A2(new_n523), .ZN(new_n698));
  NAND2_X1  g561(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n699));
  NOR2_X1   g562(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g563(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  OR2_X1    g564(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n702));
  AOI21_X1  g565(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(G1351gat));
  NOR3_X1   g566(.A1(new_n673), .A2(new_n334), .A3(new_n389), .ZN(new_n704));
  AOI21_X1  g567(.A(G197gat), .B1(new_n704), .B2(new_n555), .ZN(new_n705));
  NOR2_X1   g568(.A1(new_n389), .A2(new_n334), .ZN(new_n706));
  AND3_X1   g569(.A1(new_n657), .A2(new_n555), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g570(.A(new_n705), .B1(G197gat), .B2(new_n707), .ZN(G1352gat));
  NAND3_X1  g571(.A1(new_n657), .A2(new_n492), .A3(new_n706), .ZN(new_n709));
  NAND2_X1  g572(.A1(new_n709), .A2(G204gat), .ZN(new_n710));
  NOR2_X1   g573(.A1(new_n511), .A2(G204gat), .ZN(new_n711));
  AND3_X1   g574(.A1(new_n704), .A2(KEYINPUT62), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g575(.A(KEYINPUT62), .B1(new_n704), .B2(new_n711), .ZN(new_n713));
  OAI21_X1  g576(.A(new_n710), .B1(new_n712), .B2(new_n713), .ZN(G1353gat));
  NAND3_X1  g577(.A1(new_n704), .A2(new_n258), .A3(new_n469), .ZN(new_n715));
  NAND4_X1  g578(.A1(new_n668), .A2(new_n252), .A3(new_n469), .A4(new_n706), .ZN(new_n716));
  AND3_X1   g579(.A1(new_n716), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n717));
  AOI21_X1  g580(.A(KEYINPUT63), .B1(new_n716), .B2(G211gat), .ZN(new_n718));
  OAI21_X1  g581(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(G1354gat));
  NAND3_X1  g582(.A1(new_n704), .A2(new_n259), .A3(new_n523), .ZN(new_n720));
  AND3_X1   g583(.A1(new_n657), .A2(new_n523), .A3(new_n706), .ZN(new_n721));
  OAI21_X1  g584(.A(new_n720), .B1(new_n721), .B2(new_n259), .ZN(G1355gat));
endmodule


