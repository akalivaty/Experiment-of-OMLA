//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1204, new_n1205, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0002(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n203));
  INV_X1    g0003(.A(G87), .ZN(new_n204));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G257), .ZN(new_n207));
  OAI221_X1 g0007(.A(new_n203), .B1(new_n204), .B2(new_n205), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(KEYINPUT66), .ZN(new_n209));
  XOR2_X1   g0009(.A(KEYINPUT65), .B(G238), .Z(new_n210));
  AOI21_X1  g0010(.A(new_n209), .B1(G68), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(KEYINPUT66), .ZN(new_n212));
  INV_X1    g0012(.A(G116), .ZN(new_n213));
  INV_X1    g0013(.A(G270), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n211), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G77), .B2(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G1), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n220), .A2(new_n221), .ZN(new_n224));
  INV_X1    g0024(.A(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n205), .B(new_n226), .C1(new_n207), .C2(new_n227), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n228), .A2(KEYINPUT0), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n221), .ZN(new_n231));
  INV_X1    g0031(.A(G58), .ZN(new_n232));
  INV_X1    g0032(.A(G68), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n231), .A2(G50), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n228), .A2(KEYINPUT0), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n229), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT64), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n223), .A2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G264), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n214), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G358));
  XNOR2_X1  g0048(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(G68), .B(G77), .Z(new_n254));
  XNOR2_X1  g0054(.A(G50), .B(G58), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  OAI21_X1  g0057(.A(G20), .B1(new_n234), .B2(G50), .ZN(new_n258));
  INV_X1    g0058(.A(G150), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n221), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n221), .A2(G33), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  OAI221_X1 g0063(.A(new_n258), .B1(new_n259), .B2(new_n261), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n230), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n225), .A2(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G20), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n264), .A2(new_n266), .B1(new_n217), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n266), .B1(new_n220), .B2(G20), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n270), .B1(new_n217), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT9), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G222), .ZN(new_n280));
  INV_X1    g0080(.A(G223), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n278), .B(new_n280), .C1(new_n281), .C2(new_n279), .ZN(new_n282));
  AND2_X1   g0082(.A1(G1), .A2(G13), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n282), .B(new_n286), .C1(G77), .C2(new_n278), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n220), .B1(G41), .B2(G45), .ZN(new_n288));
  INV_X1    g0088(.A(G274), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n285), .A2(new_n288), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n287), .B(new_n291), .C1(new_n218), .C2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(KEYINPUT72), .B1(new_n293), .B2(G200), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n293), .A2(KEYINPUT72), .A3(G200), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n274), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT10), .ZN(new_n300));
  INV_X1    g0100(.A(G77), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n263), .A2(new_n261), .B1(new_n221), .B2(new_n301), .ZN(new_n302));
  XOR2_X1   g0102(.A(new_n302), .B(KEYINPUT71), .Z(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT15), .B(G87), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(new_n262), .B2(new_n304), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n305), .A2(new_n266), .B1(new_n301), .B2(new_n269), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n301), .B2(new_n272), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n210), .A2(G1698), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(new_n278), .C1(new_n241), .C2(G1698), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n309), .B(new_n286), .C1(G107), .C2(new_n278), .ZN(new_n310));
  INV_X1    g0110(.A(new_n292), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G244), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n291), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n307), .B1(G190), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G200), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(new_n314), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n307), .B(new_n319), .C1(G179), .C2(new_n313), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n293), .A2(new_n318), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n273), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT69), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n293), .A2(G179), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT70), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n300), .A2(new_n317), .A3(new_n320), .A4(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT73), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(new_n328), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G97), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n241), .A2(G1698), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(G226), .B2(G1698), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n276), .A2(new_n277), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n290), .B1(new_n335), .B2(new_n286), .ZN(new_n336));
  INV_X1    g0136(.A(G238), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n292), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n338), .A2(KEYINPUT13), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(KEYINPUT13), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(KEYINPUT74), .A3(new_n340), .ZN(new_n341));
  OR3_X1    g0141(.A1(new_n338), .A2(KEYINPUT74), .A3(KEYINPUT13), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G190), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n261), .A2(new_n217), .B1(new_n262), .B2(new_n301), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n221), .A2(G68), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n266), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT11), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n347), .A2(new_n348), .B1(G68), .B2(new_n271), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n267), .A2(new_n346), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT75), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT12), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n352), .B2(new_n353), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n349), .A2(new_n350), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n339), .A2(new_n340), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G200), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n344), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G179), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n341), .B2(new_n342), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT14), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n359), .B2(G169), .ZN(new_n365));
  AOI211_X1 g0165(.A(KEYINPUT14), .B(new_n318), .C1(new_n339), .C2(new_n340), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n361), .B1(new_n367), .B2(new_n358), .ZN(new_n368));
  XNOR2_X1  g0168(.A(G58), .B(G68), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G20), .ZN(new_n370));
  INV_X1    g0170(.A(G159), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(new_n261), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AND2_X1   g0173(.A1(KEYINPUT76), .A2(G33), .ZN(new_n374));
  NOR2_X1   g0174(.A1(KEYINPUT76), .A2(G33), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT3), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n276), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT78), .B(KEYINPUT7), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n221), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT77), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n376), .A2(new_n381), .A3(new_n276), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n381), .B1(new_n376), .B2(new_n276), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n221), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI211_X1 g0186(.A(KEYINPUT16), .B(new_n373), .C1(new_n386), .C2(new_n233), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT16), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT76), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n260), .ZN(new_n390));
  NAND2_X1  g0190(.A1(KEYINPUT76), .A2(G33), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n277), .B1(new_n392), .B2(KEYINPUT3), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(KEYINPUT7), .A3(new_n221), .ZN(new_n394));
  INV_X1    g0194(.A(new_n378), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n278), .B2(G20), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n233), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n388), .B1(new_n397), .B2(new_n372), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n387), .A2(new_n266), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n281), .A2(new_n279), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n218), .A2(G1698), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n376), .A2(new_n276), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G87), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n285), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n290), .B1(new_n311), .B2(G232), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(G190), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n263), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(new_n268), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n271), .B2(new_n408), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n399), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n406), .ZN(new_n412));
  OAI21_X1  g0212(.A(G200), .B1(new_n412), .B2(new_n404), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(KEYINPUT17), .A3(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n399), .A2(new_n413), .A3(new_n407), .A4(new_n410), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT17), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n318), .B1(new_n405), .B2(new_n406), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n412), .A2(new_n404), .A3(new_n362), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n399), .B2(new_n410), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(KEYINPUT18), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT18), .ZN(new_n423));
  AOI211_X1 g0223(.A(new_n423), .B(new_n420), .C1(new_n399), .C2(new_n410), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n414), .B(new_n417), .C1(new_n422), .C2(new_n424), .ZN(new_n425));
  NOR4_X1   g0225(.A1(new_n329), .A2(new_n330), .A3(new_n368), .A4(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT24), .ZN(new_n427));
  XNOR2_X1  g0227(.A(KEYINPUT89), .B(KEYINPUT22), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n278), .A2(new_n221), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n376), .A2(new_n221), .A3(G87), .A4(new_n276), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n429), .A2(G87), .B1(new_n430), .B2(KEYINPUT22), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n392), .A2(new_n213), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n221), .ZN(new_n433));
  INV_X1    g0233(.A(G107), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G20), .ZN(new_n435));
  XOR2_X1   g0235(.A(new_n435), .B(KEYINPUT23), .Z(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n427), .B1(new_n431), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n430), .A2(KEYINPUT22), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n278), .A2(new_n221), .A3(G87), .A4(new_n428), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n441), .A2(KEYINPUT24), .A3(new_n433), .A4(new_n436), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n438), .A2(new_n442), .A3(new_n266), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n265), .A2(new_n230), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(new_n268), .C1(G1), .C2(new_n260), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G107), .ZN(new_n447));
  INV_X1    g0247(.A(new_n267), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(new_n435), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT25), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n443), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n205), .A2(new_n279), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n207), .A2(G1698), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n376), .A2(new_n276), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n374), .A2(new_n375), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G294), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n285), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G41), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(KEYINPUT5), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n220), .A2(G45), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT83), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT5), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G41), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT83), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(new_n220), .A4(G45), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n458), .A2(KEYINPUT5), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n289), .B1(new_n283), .B2(new_n284), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n461), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  OR2_X1    g0268(.A1(new_n468), .A2(KEYINPUT84), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(KEYINPUT84), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n457), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n461), .A2(new_n466), .A3(new_n465), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(G264), .A3(new_n285), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT90), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n472), .A2(KEYINPUT90), .A3(G264), .A4(new_n285), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n471), .A2(new_n477), .A3(G179), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n454), .A2(new_n456), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n286), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n468), .A2(KEYINPUT84), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n468), .A2(KEYINPUT84), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n480), .B(new_n473), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G169), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n478), .A2(new_n484), .A3(KEYINPUT91), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT91), .B1(new_n478), .B2(new_n484), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n451), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT92), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT92), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n489), .B(new_n451), .C1(new_n485), .C2(new_n486), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT93), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n471), .A2(new_n477), .ZN(new_n492));
  INV_X1    g0292(.A(new_n483), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n316), .A2(new_n492), .B1(new_n493), .B2(new_n295), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n491), .B1(new_n494), .B2(new_n451), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n443), .A2(new_n447), .A3(new_n450), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n492), .A2(new_n316), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n493), .A2(new_n295), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n496), .A2(new_n499), .A3(KEYINPUT93), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n488), .A2(new_n490), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT87), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n446), .A2(G116), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n269), .A2(new_n213), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n505), .B(new_n221), .C1(G33), .C2(new_n206), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n506), .B(new_n266), .C1(new_n221), .C2(G116), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT20), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n507), .A2(new_n508), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n503), .B(new_n504), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n207), .A2(new_n279), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n227), .A2(G1698), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n376), .A2(new_n276), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n334), .A2(G303), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n286), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n472), .A2(G270), .A3(new_n285), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n518), .B(new_n519), .C1(new_n481), .C2(new_n482), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n512), .B1(new_n295), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(G200), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n502), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n520), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G190), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n526), .A2(KEYINPUT87), .A3(new_n512), .A4(new_n522), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n520), .A2(new_n511), .A3(G169), .ZN(new_n529));
  NOR2_X1   g0329(.A1(KEYINPUT86), .A2(KEYINPUT21), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n525), .A2(G179), .A3(new_n511), .ZN(new_n532));
  INV_X1    g0332(.A(new_n530), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n520), .A2(new_n511), .A3(G169), .A4(new_n533), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT88), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT88), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n528), .A2(new_n538), .A3(new_n535), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n376), .A2(new_n221), .A3(G68), .A4(new_n276), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT19), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n262), .B2(new_n206), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n221), .B1(new_n331), .B2(new_n542), .ZN(new_n544));
  NOR2_X1   g0344(.A1(G97), .A2(G107), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n204), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n541), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(new_n266), .B1(new_n304), .B2(new_n269), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n304), .B2(new_n445), .ZN(new_n550));
  INV_X1    g0350(.A(new_n432), .ZN(new_n551));
  NOR2_X1   g0351(.A1(G238), .A2(G1698), .ZN(new_n552));
  INV_X1    g0352(.A(G244), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n553), .B2(G1698), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(new_n376), .A3(new_n276), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n285), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n460), .A2(G274), .ZN(new_n557));
  AOI21_X1  g0357(.A(G250), .B1(new_n220), .B2(G45), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n286), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n362), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n550), .B(new_n561), .C1(G169), .C2(new_n560), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(G190), .ZN(new_n563));
  OAI21_X1  g0363(.A(G200), .B1(new_n556), .B2(new_n559), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n446), .A2(G87), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n549), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n553), .A2(G1698), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n376), .A2(new_n276), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT81), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT4), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT81), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n376), .A2(new_n572), .A3(new_n276), .A4(new_n568), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n568), .A2(KEYINPUT4), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n205), .B2(new_n279), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(new_n278), .B1(G33), .B2(G283), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n286), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT82), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n469), .A2(new_n470), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n472), .A2(G257), .A3(new_n285), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n285), .B1(new_n574), .B2(new_n577), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT82), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n581), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n582), .A2(new_n583), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(new_n585), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n587), .A2(G200), .B1(G190), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n445), .A2(new_n206), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n268), .A2(G97), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n434), .A2(G97), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT79), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n596), .A2(KEYINPUT6), .B1(new_n434), .B2(G97), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT6), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(KEYINPUT79), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n597), .A2(KEYINPUT80), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT80), .ZN(new_n601));
  AOI22_X1  g0401(.A1(KEYINPUT79), .A2(new_n598), .B1(new_n206), .B2(G107), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n596), .A2(KEYINPUT6), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n595), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT80), .B1(new_n597), .B2(new_n599), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n602), .A2(new_n601), .A3(new_n603), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(G97), .A4(new_n434), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n221), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n434), .B1(new_n394), .B2(new_n396), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n261), .A2(new_n301), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n592), .B(new_n594), .C1(new_n612), .C2(new_n444), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n581), .A2(new_n362), .A3(new_n584), .A4(new_n586), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n318), .B1(new_n588), .B2(new_n585), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n616), .A3(new_n613), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT85), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n615), .A2(new_n613), .A3(KEYINPUT85), .A4(new_n616), .ZN(new_n620));
  AOI221_X4 g0420(.A(new_n567), .B1(new_n590), .B2(new_n614), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n426), .A2(new_n501), .A3(new_n540), .A4(new_n621), .ZN(G372));
  NAND2_X1  g0422(.A1(new_n619), .A2(new_n620), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n564), .A2(new_n549), .A3(new_n565), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT94), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT94), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n564), .A2(new_n549), .A3(new_n626), .A4(new_n565), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n563), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n562), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n500), .B2(new_n495), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n590), .A2(new_n614), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n623), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT95), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n478), .A2(new_n484), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n451), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n535), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g0436(.A(new_n636), .B(KEYINPUT96), .Z(new_n637));
  INV_X1    g0437(.A(KEYINPUT95), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n623), .A2(new_n630), .A3(new_n638), .A4(new_n631), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n633), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n615), .A2(new_n616), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT97), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n615), .A2(KEYINPUT97), .A3(new_n616), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n614), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  INV_X1    g0446(.A(new_n629), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n567), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n619), .A2(new_n649), .A3(new_n620), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT26), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n648), .A2(new_n562), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n640), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n426), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n367), .A2(new_n358), .ZN(new_n655));
  INV_X1    g0455(.A(new_n361), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n655), .B1(new_n656), .B2(new_n320), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(new_n417), .A3(new_n414), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n422), .A2(new_n424), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n660), .A2(new_n300), .B1(new_n325), .B2(new_n323), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n654), .A2(new_n661), .ZN(G369));
  INV_X1    g0462(.A(new_n535), .ZN(new_n663));
  OR3_X1    g0463(.A1(new_n448), .A2(KEYINPUT27), .A3(G20), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT27), .B1(new_n448), .B2(G20), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n512), .A2(new_n669), .ZN(new_n670));
  MUX2_X1   g0470(.A(new_n540), .B(new_n663), .S(new_n670), .Z(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n501), .B1(new_n496), .B2(new_n669), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n487), .B2(new_n669), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n535), .A2(new_n668), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n501), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n451), .A2(new_n634), .A3(new_n669), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT98), .Z(G399));
  NOR2_X1   g0483(.A1(new_n226), .A2(G41), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G1), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n545), .A2(new_n204), .A3(new_n213), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n234), .A2(G50), .ZN(new_n688));
  OAI22_X1  g0488(.A1(new_n686), .A2(new_n687), .B1(new_n688), .B2(new_n685), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n621), .A2(new_n540), .A3(new_n501), .A4(new_n669), .ZN(new_n691));
  INV_X1    g0491(.A(new_n492), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n520), .A2(new_n362), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n589), .A2(new_n692), .A3(new_n693), .A4(new_n560), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT30), .Z(new_n695));
  XNOR2_X1  g0495(.A(new_n560), .B(KEYINPUT99), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n587), .A2(new_n520), .A3(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n697), .A2(G179), .A3(new_n692), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n668), .B1(new_n695), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n699), .A2(KEYINPUT31), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n645), .A2(KEYINPUT100), .A3(KEYINPUT26), .A4(new_n647), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n663), .B1(new_n488), .B2(new_n490), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n704), .B(new_n562), .C1(new_n632), .C2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n650), .A2(new_n646), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n643), .A2(new_n644), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(KEYINPUT26), .A3(new_n613), .A4(new_n647), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT100), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  OAI211_X1 g0511(.A(KEYINPUT29), .B(new_n669), .C1(new_n706), .C2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n668), .B1(new_n640), .B2(new_n652), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(KEYINPUT29), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n703), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n690), .B1(new_n716), .B2(G1), .ZN(G364));
  NOR2_X1   g0517(.A1(G13), .A2(G33), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G20), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n671), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n221), .A2(G179), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(new_n295), .A3(new_n316), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n295), .A2(new_n316), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n723), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n725), .A2(G329), .B1(new_n728), .B2(G303), .ZN(new_n729));
  INV_X1    g0529(.A(G294), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n295), .A2(G179), .A3(G200), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n221), .ZN(new_n732));
  INV_X1    g0532(.A(G322), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n221), .A2(new_n362), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n735), .A2(new_n295), .A3(G200), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI221_X1 g0537(.A(new_n729), .B1(new_n730), .B2(new_n732), .C1(new_n733), .C2(new_n737), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n735), .A2(new_n316), .A3(G190), .ZN(new_n739));
  XNOR2_X1  g0539(.A(KEYINPUT33), .B(G317), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n734), .A2(new_n726), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G326), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n723), .A2(new_n295), .A3(G200), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT101), .Z(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G283), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n735), .A2(G190), .A3(G200), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n278), .B1(new_n749), .B2(G311), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n741), .A2(new_n744), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n732), .A2(new_n206), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT32), .B1(new_n724), .B2(new_n371), .ZN(new_n753));
  INV_X1    g0553(.A(new_n749), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n753), .B1(new_n217), .B2(new_n742), .C1(new_n754), .C2(new_n301), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n752), .B(new_n755), .C1(G68), .C2(new_n739), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n727), .A2(new_n204), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n334), .B(new_n757), .C1(new_n747), .C2(G107), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n725), .A2(G159), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n756), .B(new_n758), .C1(KEYINPUT32), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n737), .A2(new_n232), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n751), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n230), .B1(G20), .B2(new_n318), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n226), .A2(new_n334), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G355), .ZN(new_n766));
  INV_X1    g0566(.A(new_n226), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n382), .A2(new_n383), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n226), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(G45), .B2(new_n688), .ZN(new_n770));
  INV_X1    g0570(.A(G45), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n256), .A2(new_n771), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n766), .B1(G116), .B2(new_n767), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n720), .A2(new_n763), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n225), .A2(G20), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n686), .B1(G45), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n722), .A2(new_n764), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n671), .A2(G330), .ZN(new_n779));
  INV_X1    g0579(.A(new_n777), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n672), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n778), .B1(new_n779), .B2(new_n781), .ZN(G396));
  OR2_X1    g0582(.A1(new_n320), .A2(new_n668), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n307), .A2(new_n668), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n317), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n784), .B1(new_n320), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n653), .A2(new_n669), .A3(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT102), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n703), .B(new_n790), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n713), .A2(new_n787), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n780), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n787), .A2(new_n719), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n763), .A2(new_n718), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n301), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n752), .B1(G303), .B2(new_n743), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n730), .B2(new_n737), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n278), .B(new_n799), .C1(G283), .C2(new_n739), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n749), .A2(G116), .B1(G311), .B2(new_n725), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n800), .B(new_n801), .C1(new_n434), .C2(new_n727), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G87), .B2(new_n747), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n768), .B1(new_n217), .B2(new_n727), .C1(new_n746), .C2(new_n233), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G143), .A2(new_n736), .B1(new_n749), .B2(G159), .ZN(new_n805));
  INV_X1    g0605(.A(G137), .ZN(new_n806));
  INV_X1    g0606(.A(new_n739), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n805), .B1(new_n806), .B2(new_n742), .C1(new_n259), .C2(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT34), .Z(new_n809));
  INV_X1    g0609(.A(new_n732), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n804), .B(new_n809), .C1(G58), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n725), .A2(G132), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n803), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n763), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n797), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n777), .B1(new_n795), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n794), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT103), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n817), .B(new_n818), .ZN(G384));
  INV_X1    g0619(.A(KEYINPUT40), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n358), .A2(new_n669), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n368), .B(new_n821), .ZN(new_n822));
  AND4_X1   g0622(.A1(new_n700), .A2(new_n701), .A3(new_n822), .A4(new_n787), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n820), .B1(new_n823), .B2(KEYINPUT107), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n700), .A2(new_n701), .A3(new_n822), .A4(new_n787), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT107), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n399), .A2(new_n410), .ZN(new_n828));
  INV_X1    g0628(.A(new_n666), .ZN(new_n829));
  AOI21_X1  g0629(.A(KEYINPUT105), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT105), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n831), .B(new_n666), .C1(new_n399), .C2(new_n410), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n828), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n415), .B1(new_n834), .B2(new_n420), .ZN(new_n835));
  OAI21_X1  g0635(.A(KEYINPUT37), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n421), .B1(new_n411), .B2(new_n413), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT37), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n837), .B(new_n838), .C1(new_n830), .C2(new_n832), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n836), .A2(KEYINPUT106), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n425), .A2(new_n833), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n833), .A2(new_n835), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT106), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n842), .A2(new_n843), .A3(new_n838), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n840), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT38), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n410), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n275), .B1(new_n390), .B2(new_n391), .ZN(new_n849));
  INV_X1    g0649(.A(new_n276), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT77), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n376), .A2(new_n381), .A3(new_n276), .ZN(new_n852));
  AOI21_X1  g0652(.A(G20), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n379), .B1(new_n853), .B2(KEYINPUT7), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n372), .B1(new_n854), .B2(G68), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n444), .B1(new_n855), .B2(KEYINPUT16), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n373), .B1(new_n386), .B2(new_n233), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n388), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n848), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n859), .A2(new_n666), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n425), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n415), .B1(new_n859), .B2(new_n420), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n860), .B1(new_n862), .B2(KEYINPUT104), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT104), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n415), .B(new_n864), .C1(new_n859), .C2(new_n420), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n838), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n833), .A2(KEYINPUT37), .A3(new_n835), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n861), .B(KEYINPUT38), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n847), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT108), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n847), .A2(KEYINPUT108), .A3(new_n868), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n824), .A2(new_n827), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n861), .B1(new_n866), .B2(new_n867), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n846), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n868), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n820), .B1(new_n877), .B2(new_n825), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n426), .A2(new_n702), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n879), .B(new_n880), .Z(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(G330), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n655), .A2(new_n668), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n875), .A2(KEYINPUT39), .A3(new_n868), .ZN(new_n884));
  INV_X1    g0684(.A(new_n868), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n846), .B2(new_n845), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n883), .B(new_n884), .C1(new_n886), .C2(KEYINPUT39), .ZN(new_n887));
  INV_X1    g0687(.A(new_n822), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n788), .B2(new_n783), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n876), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n659), .A2(new_n829), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n887), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n426), .B(new_n712), .C1(new_n713), .C2(KEYINPUT29), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n661), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n892), .B(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n882), .B(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n220), .B2(new_n776), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n605), .A2(new_n608), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n213), .B1(new_n898), .B2(KEYINPUT35), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n899), .B(new_n231), .C1(KEYINPUT35), .C2(new_n898), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT36), .ZN(new_n901));
  OAI21_X1  g0701(.A(G77), .B1(new_n232), .B2(new_n233), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n688), .A2(new_n902), .B1(G50), .B2(new_n233), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(G1), .A3(new_n225), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n897), .A2(new_n901), .A3(new_n904), .ZN(G367));
  INV_X1    g0705(.A(KEYINPUT111), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n623), .A2(new_n631), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n614), .A2(new_n669), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n645), .A2(new_n668), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n906), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n910), .B(KEYINPUT111), .C1(new_n907), .C2(new_n908), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n678), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT42), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n916), .B(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n914), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n488), .A2(new_n490), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n623), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n669), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n549), .A2(new_n565), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n668), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n647), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT109), .Z(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n562), .B2(new_n925), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT110), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT43), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n923), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n918), .A2(new_n930), .A3(new_n922), .A4(new_n929), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n676), .A2(new_n919), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT112), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n933), .A2(new_n934), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n676), .B2(new_n919), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n684), .B(KEYINPUT41), .Z(new_n940));
  NAND2_X1  g0740(.A1(new_n919), .A2(new_n680), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n941), .A2(KEYINPUT44), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(KEYINPUT44), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT45), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n919), .A2(new_n945), .A3(new_n680), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT45), .B1(new_n914), .B2(new_n681), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n673), .B(new_n675), .C1(new_n944), .C2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n948), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n950), .A2(new_n676), .A3(new_n943), .A4(new_n942), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n678), .B1(new_n675), .B2(new_n677), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(new_n672), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n715), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n949), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n940), .B1(new_n955), .B2(new_n716), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n776), .A2(G45), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(G1), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT113), .Z(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n937), .B(new_n939), .C1(new_n956), .C2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n929), .A2(new_n720), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n732), .A2(new_n233), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(G150), .B2(new_n736), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT114), .Z(new_n965));
  OAI22_X1  g0765(.A1(new_n724), .A2(new_n806), .B1(new_n745), .B2(new_n301), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n334), .B(new_n966), .C1(G143), .C2(new_n743), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n217), .B2(new_n754), .C1(new_n232), .C2(new_n727), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n807), .A2(new_n371), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n732), .A2(new_n434), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n728), .A2(G116), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT46), .Z(new_n973));
  INV_X1    g0773(.A(new_n768), .ZN(new_n974));
  INV_X1    g0774(.A(G317), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n975), .B2(new_n724), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n743), .A2(G311), .ZN(new_n977));
  INV_X1    g0777(.A(G283), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n977), .B1(new_n807), .B2(new_n730), .C1(new_n978), .C2(new_n754), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n736), .A2(G303), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n206), .B2(new_n745), .ZN(new_n981));
  OR4_X1    g0781(.A1(new_n973), .A2(new_n976), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n969), .A2(new_n970), .B1(new_n971), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT47), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n763), .ZN(new_n985));
  INV_X1    g0785(.A(new_n769), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n774), .B1(new_n767), .B2(new_n304), .C1(new_n986), .C2(new_n247), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n962), .A2(new_n777), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n961), .A2(new_n988), .ZN(G387));
  INV_X1    g0789(.A(new_n954), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n685), .B1(new_n715), .B2(new_n953), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n974), .B1(new_n213), .B2(new_n745), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G303), .A2(new_n749), .B1(new_n739), .B2(G311), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n975), .B2(new_n737), .C1(new_n733), .C2(new_n742), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT48), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n978), .B2(new_n732), .C1(new_n730), .C2(new_n727), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT49), .Z(new_n998));
  AOI211_X1 g0798(.A(new_n993), .B(new_n998), .C1(G326), .C2(new_n725), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n408), .A2(new_n739), .B1(new_n749), .B2(G68), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n732), .A2(new_n304), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G159), .B2(new_n743), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n736), .A2(G50), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1000), .A2(new_n1002), .A3(new_n768), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n728), .A2(G77), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n259), .B2(new_n724), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT115), .Z(new_n1007));
  AOI211_X1 g0807(.A(new_n1004), .B(new_n1007), .C1(G97), .C2(new_n747), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n763), .B1(new_n999), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n986), .B1(new_n244), .B2(G45), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n687), .B2(new_n765), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n408), .A2(new_n217), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT50), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n233), .A2(new_n301), .ZN(new_n1014));
  NOR4_X1   g0814(.A1(new_n1013), .A2(G45), .A3(new_n1014), .A4(new_n687), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1011), .A2(new_n1015), .B1(G107), .B2(new_n767), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n780), .B1(new_n1016), .B2(new_n774), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1009), .B(new_n1017), .C1(new_n675), .C2(new_n721), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n992), .B(new_n1018), .C1(new_n953), .C2(new_n959), .ZN(G393));
  NAND2_X1  g0819(.A1(new_n919), .A2(new_n720), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n774), .B1(new_n206), .B2(new_n767), .C1(new_n986), .C2(new_n253), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n754), .A2(new_n730), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n736), .A2(G311), .B1(new_n743), .B2(G317), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT52), .Z(new_n1024));
  NAND2_X1  g0824(.A1(new_n728), .A2(G283), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n747), .A2(G107), .B1(G303), .B2(new_n739), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n278), .B1(new_n725), .B2(G322), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1022), .B(new_n1028), .C1(G116), .C2(new_n810), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n736), .A2(G159), .B1(new_n743), .B2(G150), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT51), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G77), .B2(new_n810), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n725), .A2(G143), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n747), .A2(G87), .B1(G50), .B2(new_n739), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n974), .B1(G68), .B2(new_n728), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n408), .B2(new_n749), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n763), .B1(new_n1029), .B2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1020), .A2(new_n777), .A3(new_n1021), .A4(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n949), .A2(new_n951), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1039), .B1(new_n1040), .B2(new_n959), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n685), .B1(new_n1040), .B2(new_n990), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1041), .B1(new_n955), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(G390));
  INV_X1    g0844(.A(KEYINPUT116), .ZN(new_n1045));
  AOI21_X1  g0845(.A(KEYINPUT39), .B1(new_n847), .B2(new_n868), .ZN(new_n1046));
  AND3_X1   g0846(.A1(new_n875), .A2(KEYINPUT39), .A3(new_n868), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n889), .A2(new_n883), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n786), .A2(new_n320), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n669), .B(new_n1049), .C1(new_n706), .C2(new_n711), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n783), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n822), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n883), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n871), .A2(new_n1052), .A3(new_n872), .A4(new_n1053), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n700), .A2(G330), .A3(new_n701), .A4(new_n787), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1055), .A2(new_n888), .ZN(new_n1056));
  AND3_X1   g0856(.A1(new_n1048), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1056), .B1(new_n1048), .B2(new_n1054), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n426), .A2(new_n702), .A3(G330), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n893), .A2(new_n661), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n788), .A2(new_n783), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1055), .A2(new_n888), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1055), .A2(new_n888), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1056), .A2(new_n783), .A3(new_n1063), .A4(new_n1050), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1061), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1045), .B1(new_n1059), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1048), .A2(new_n1054), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n1065), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1048), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1071), .A2(new_n1068), .A3(new_n1045), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n684), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT117), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1068), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1071), .A2(new_n1068), .A3(new_n1072), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(KEYINPUT116), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1073), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1083), .A2(KEYINPUT117), .A3(new_n684), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1077), .A2(new_n1080), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1059), .A2(new_n960), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT118), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1086), .B(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n718), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n796), .A2(new_n263), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT54), .B(G143), .Z(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n754), .A2(new_n1092), .B1(new_n371), .B2(new_n732), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G137), .B2(new_n739), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT119), .Z(new_n1095));
  NAND2_X1  g0895(.A1(new_n728), .A2(G150), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT53), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n278), .B1(new_n745), .B2(new_n217), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n1095), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n725), .A2(G125), .ZN(new_n1100));
  INV_X1    g0900(.A(G128), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1099), .B(new_n1100), .C1(new_n1101), .C2(new_n742), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G132), .B2(new_n736), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n807), .A2(new_n434), .B1(new_n730), .B2(new_n724), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n757), .B(new_n1104), .C1(G97), .C2(new_n749), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n278), .B1(new_n743), .B2(G283), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n747), .A2(G68), .B1(G77), .B2(new_n810), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G116), .B2(new_n736), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n763), .B1(new_n1103), .B2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1089), .A2(new_n777), .A3(new_n1090), .A4(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1088), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1085), .A2(new_n1112), .ZN(G378));
  NAND3_X1  g0913(.A1(new_n871), .A2(new_n827), .A3(new_n872), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT40), .B1(new_n825), .B2(new_n826), .ZN(new_n1115));
  OAI211_X1 g0915(.A(G330), .B(new_n878), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n892), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n300), .A2(new_n326), .ZN(new_n1118));
  XOR2_X1   g0918(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1119));
  XNOR2_X1  g0919(.A(new_n1118), .B(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n273), .A2(new_n829), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT122), .Z(new_n1122));
  XOR2_X1   g0922(.A(new_n1120), .B(new_n1122), .Z(new_n1123));
  NAND3_X1  g0923(.A1(new_n887), .A2(new_n890), .A3(new_n891), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1124), .A2(new_n873), .A3(G330), .A4(new_n878), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1117), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1123), .B1(new_n1117), .B2(new_n1125), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n960), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n780), .B1(new_n1123), .B2(new_n718), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n796), .A2(new_n217), .ZN(new_n1130));
  INV_X1    g0930(.A(G124), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n260), .B1(new_n724), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n739), .A2(G132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n754), .B2(new_n806), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1092), .A2(new_n727), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT120), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1134), .B(new_n1136), .C1(G150), .C2(new_n810), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n743), .A2(G125), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1137), .B(new_n1138), .C1(new_n1101), .C2(new_n737), .ZN(new_n1139));
  AOI211_X1 g0939(.A(G41), .B(new_n1132), .C1(new_n1139), .C2(KEYINPUT59), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1140), .B1(KEYINPUT59), .B2(new_n1139), .C1(new_n371), .C2(new_n745), .ZN(new_n1141));
  AOI21_X1  g0941(.A(G41), .B1(new_n768), .B2(G33), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1141), .B1(G50), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n745), .A2(new_n232), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n754), .A2(new_n304), .B1(new_n742), .B2(new_n213), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(G283), .C2(new_n725), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n458), .B1(new_n807), .B2(new_n206), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n963), .B(new_n1147), .C1(G107), .C2(new_n736), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1146), .A2(new_n1148), .A3(new_n974), .A4(new_n1005), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT58), .Z(new_n1150));
  OAI21_X1  g0950(.A(new_n763), .B1(new_n1143), .B2(new_n1150), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT121), .Z(new_n1152));
  NAND3_X1  g0952(.A1(new_n1129), .A2(new_n1130), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1061), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1083), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1127), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1117), .A2(new_n1125), .A3(new_n1123), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT57), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1061), .B1(new_n1082), .B2(new_n1073), .ZN(new_n1160));
  OAI21_X1  g0960(.A(KEYINPUT57), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n684), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1128), .B(new_n1153), .C1(new_n1159), .C2(new_n1162), .ZN(G375));
  NAND3_X1  g0963(.A1(new_n1061), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n940), .B(KEYINPUT123), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1079), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n334), .B1(new_n206), .B2(new_n727), .C1(new_n737), .C2(new_n978), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1001), .B(new_n1167), .C1(G116), .C2(new_n739), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G294), .A2(new_n743), .B1(new_n725), .B2(G303), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n301), .B2(new_n746), .C1(new_n434), .C2(new_n754), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n737), .A2(new_n806), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n725), .A2(G128), .B1(new_n728), .B2(G159), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n259), .B2(new_n754), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1144), .B(new_n1174), .C1(G50), .C2(new_n810), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n743), .A2(G132), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n974), .B1(new_n739), .B2(new_n1091), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1171), .B1(new_n1172), .B2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT124), .Z(new_n1180));
  OAI221_X1 g0980(.A(new_n777), .B1(new_n822), .B2(new_n719), .C1(new_n1180), .C2(new_n814), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n233), .B2(new_n796), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1182), .B1(new_n1183), .B2(new_n960), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1166), .A2(new_n1184), .ZN(G381));
  NAND3_X1  g0985(.A1(new_n961), .A2(new_n988), .A3(new_n1043), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n817), .B(KEYINPUT103), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n1189), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1088), .A2(new_n1111), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT117), .B1(new_n1083), .B2(new_n684), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1076), .B(new_n685), .C1(new_n1082), .C2(new_n1073), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1191), .B1(new_n1194), .B2(new_n1080), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1128), .A2(new_n1153), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT57), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n685), .B1(new_n1155), .B2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1197), .B1(new_n1160), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1196), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1190), .A2(new_n1195), .A3(new_n1202), .ZN(G407));
  NOR2_X1   g1003(.A1(new_n1190), .A2(new_n667), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1195), .A2(new_n1202), .ZN(new_n1205));
  OAI21_X1  g1005(.A(G213), .B1(new_n1204), .B2(new_n1205), .ZN(G409));
  XNOR2_X1  g1006(.A(G393), .B(G396), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1043), .B1(new_n961), .B2(new_n988), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1208), .B1(new_n1187), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1209), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1211), .A2(new_n1186), .A3(new_n1207), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1160), .A2(new_n1200), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1196), .B1(new_n1214), .B2(new_n1165), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(new_n1085), .A3(new_n1112), .ZN(new_n1216));
  INV_X1    g1016(.A(G213), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1217), .A2(G343), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1216), .B(new_n1219), .C1(new_n1195), .C2(new_n1202), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT125), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT60), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1164), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1164), .A2(new_n1223), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1224), .A2(new_n684), .A3(new_n1079), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1184), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(G384), .B(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(G2897), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1219), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1188), .A2(new_n1227), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1188), .A2(new_n1227), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1232), .A2(new_n1233), .B1(new_n1229), .B2(new_n1219), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1218), .B1(G375), .B2(G378), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(KEYINPUT125), .A3(new_n1216), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1222), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT61), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT62), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1236), .A2(new_n1240), .A3(new_n1228), .A4(new_n1216), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1222), .A2(new_n1237), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1240), .B1(new_n1243), .B2(new_n1228), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1213), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(KEYINPUT63), .A3(new_n1228), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1231), .A2(new_n1234), .B1(new_n1236), .B2(new_n1216), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT63), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1228), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n1247), .A2(new_n1248), .B1(new_n1249), .B2(new_n1220), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1213), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1246), .A2(new_n1250), .A3(new_n1239), .A4(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1245), .A2(new_n1252), .ZN(G405));
  NAND3_X1  g1053(.A1(new_n1210), .A2(new_n1212), .A3(KEYINPUT126), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT127), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1254), .B(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G375), .A2(G378), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1205), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1228), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1249), .A2(new_n1205), .A3(new_n1257), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1259), .B(new_n1260), .C1(new_n1251), .C2(KEYINPUT126), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1256), .B(new_n1261), .ZN(G402));
endmodule


