//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT89), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G224), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n190), .B(KEYINPUT87), .Z(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT86), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n201), .B1(new_n196), .B2(G143), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n198), .A2(KEYINPUT64), .A3(G146), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n202), .A2(new_n203), .B1(G143), .B2(new_n196), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n194), .B1(new_n197), .B2(KEYINPUT1), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n193), .B(new_n200), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(new_n203), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n197), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n197), .A2(new_n199), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n208), .A2(new_n211), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n206), .B1(new_n213), .B2(new_n193), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n192), .B(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G110), .B(G122), .ZN(new_n217));
  XOR2_X1   g031(.A(new_n217), .B(KEYINPUT84), .Z(new_n218));
  INV_X1    g032(.A(G119), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G116), .ZN(new_n220));
  OR3_X1    g034(.A1(new_n220), .A2(KEYINPUT83), .A3(KEYINPUT5), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT83), .B1(new_n220), .B2(KEYINPUT5), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n221), .A2(G113), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G116), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G119), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT68), .ZN(new_n227));
  XNOR2_X1  g041(.A(G116), .B(G119), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT5), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n223), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT2), .A2(G113), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT2), .ZN(new_n235));
  INV_X1    g049(.A(G113), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT67), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n238), .A2(KEYINPUT2), .A3(G113), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n228), .B(new_n234), .C1(new_n237), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT69), .ZN(new_n241));
  INV_X1    g055(.A(new_n234), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT67), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n238), .B1(KEYINPUT2), .B2(G113), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(new_n228), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n241), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n233), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n250));
  INV_X1    g064(.A(G104), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(G107), .ZN(new_n252));
  INV_X1    g066(.A(G107), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT3), .A3(G104), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G101), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT79), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n257), .B1(new_n253), .B2(G104), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n251), .A2(KEYINPUT79), .A3(G107), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n255), .A2(new_n256), .A3(new_n258), .A4(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n251), .A2(G107), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n253), .A2(G104), .ZN(new_n262));
  OAI21_X1  g076(.A(G101), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n249), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n253), .A2(KEYINPUT3), .A3(G104), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT3), .B1(new_n253), .B2(G104), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n258), .B(new_n259), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(G101), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT80), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n269), .A2(KEYINPUT80), .A3(new_n270), .A4(G101), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n270), .B1(new_n269), .B2(G101), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n273), .A2(new_n274), .B1(new_n260), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n243), .A2(new_n244), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n234), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(new_n227), .A3(new_n230), .ZN(new_n279));
  AND4_X1   g093(.A1(new_n246), .A2(new_n277), .A3(new_n234), .A4(new_n228), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n246), .B1(new_n245), .B2(new_n228), .ZN(new_n281));
  OAI211_X1 g095(.A(KEYINPUT70), .B(new_n279), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT70), .B1(new_n248), .B2(new_n279), .ZN(new_n284));
  OAI211_X1 g098(.A(KEYINPUT82), .B(new_n276), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT70), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n282), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT82), .B1(new_n290), .B2(new_n276), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n218), .B(new_n266), .C1(new_n286), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT85), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT6), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n266), .B1(new_n286), .B2(new_n291), .ZN(new_n297));
  INV_X1    g111(.A(new_n218), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n298), .A3(new_n295), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n216), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT8), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n218), .B(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n249), .A2(new_n264), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n223), .B1(new_n232), .B2(new_n226), .ZN(new_n306));
  INV_X1    g120(.A(new_n264), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n248), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n304), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n191), .A2(KEYINPUT7), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n214), .A2(KEYINPUT88), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n311), .B1(new_n214), .B2(new_n310), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT88), .B1(new_n214), .B2(new_n310), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n309), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n292), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G902), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n188), .B1(new_n302), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n317), .ZN(new_n319));
  INV_X1    g133(.A(new_n188), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n276), .B1(new_n283), .B2(new_n284), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT82), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n265), .B1(new_n323), .B2(new_n285), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n324), .A2(new_n218), .A3(new_n294), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n299), .B2(new_n296), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n319), .B(new_n320), .C1(new_n326), .C2(new_n216), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n318), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(G214), .B1(G237), .B2(G902), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT9), .B(G234), .ZN(new_n330));
  OAI21_X1  g144(.A(G221), .B1(new_n330), .B2(G902), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n200), .B1(new_n204), .B2(new_n205), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n332), .A2(KEYINPUT10), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n200), .B1(new_n212), .B2(new_n205), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n260), .A3(new_n263), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT10), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n333), .A2(new_n307), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n275), .A2(new_n260), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n258), .A2(new_n259), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n256), .B1(new_n339), .B2(new_n255), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT80), .B1(new_n340), .B2(new_n270), .ZN(new_n341));
  INV_X1    g155(.A(new_n274), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n213), .B(new_n338), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT11), .ZN(new_n344));
  INV_X1    g158(.A(G134), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n344), .B1(new_n345), .B2(G137), .ZN(new_n346));
  INV_X1    g160(.A(G137), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT11), .A3(G134), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(G137), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G131), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT66), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT66), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n350), .A2(new_n353), .A3(G131), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n348), .A2(new_n349), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT65), .ZN(new_n356));
  INV_X1    g170(.A(G131), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n355), .A2(new_n356), .A3(new_n357), .A4(new_n346), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n346), .A2(new_n348), .A3(new_n357), .A4(new_n349), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT65), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n352), .A2(new_n354), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n337), .A2(new_n343), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n335), .B1(new_n307), .B2(new_n332), .ZN(new_n363));
  INV_X1    g177(.A(new_n361), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT12), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT12), .B1(new_n363), .B2(new_n364), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n362), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G110), .B(G140), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n189), .A2(G227), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  XOR2_X1   g184(.A(new_n370), .B(KEYINPUT78), .Z(new_n371));
  NAND2_X1  g185(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n361), .B1(new_n337), .B2(new_n343), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n370), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(new_n362), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n376), .A3(G469), .ZN(new_n377));
  NAND2_X1  g191(.A1(G469), .A2(G902), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n337), .A2(new_n343), .A3(new_n361), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n370), .B1(new_n380), .B2(new_n373), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n362), .B(new_n375), .C1(new_n365), .C2(new_n366), .ZN(new_n382));
  AOI211_X1 g196(.A(G469), .B(G902), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n331), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(KEYINPUT81), .B(new_n331), .C1(new_n379), .C2(new_n383), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n328), .A2(new_n329), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G472), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT71), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n283), .A2(new_n284), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n358), .A2(new_n360), .ZN(new_n393));
  INV_X1    g207(.A(new_n349), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n345), .A2(G137), .ZN(new_n395));
  OAI21_X1  g209(.A(G131), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n332), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n208), .A2(new_n211), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n212), .A2(new_n209), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n397), .B1(new_n361), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT30), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT30), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n397), .B(new_n403), .C1(new_n361), .C2(new_n400), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n392), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n350), .A2(new_n353), .A3(G131), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n353), .B1(new_n350), .B2(G131), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n359), .B(new_n356), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n213), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n410), .A2(new_n289), .A3(new_n282), .A4(new_n397), .ZN(new_n411));
  INV_X1    g225(.A(G237), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n189), .A3(G210), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT27), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT26), .B(G101), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n391), .B1(new_n405), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n404), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n403), .B1(new_n410), .B2(new_n397), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n290), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n416), .ZN(new_n422));
  INV_X1    g236(.A(new_n401), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n422), .B1(new_n423), .B2(new_n392), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n421), .A2(new_n424), .A3(KEYINPUT71), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n418), .A2(new_n425), .A3(KEYINPUT31), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT28), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n290), .A2(new_n401), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n427), .B1(new_n428), .B2(new_n411), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT28), .B1(new_n423), .B2(new_n392), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n422), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT31), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n421), .A2(new_n432), .A3(new_n424), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n390), .B(new_n316), .C1(new_n426), .C2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT32), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT72), .ZN(new_n438));
  INV_X1    g252(.A(new_n434), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n418), .A2(new_n425), .A3(KEYINPUT31), .ZN(new_n440));
  AOI21_X1  g254(.A(G902), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT32), .A3(new_n390), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT29), .ZN(new_n443));
  NOR4_X1   g257(.A1(new_n429), .A2(new_n430), .A3(new_n443), .A4(new_n422), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT74), .B1(new_n444), .B2(G902), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT74), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n290), .A2(new_n401), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n410), .A2(new_n397), .B1(new_n289), .B2(new_n282), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT28), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n411), .A2(new_n427), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n416), .A3(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n446), .B(new_n316), .C1(new_n451), .C2(new_n443), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(KEYINPUT73), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n421), .A2(new_n411), .ZN(new_n454));
  AOI21_X1  g268(.A(KEYINPUT29), .B1(new_n454), .B2(new_n422), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n451), .A2(KEYINPUT73), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n445), .B(new_n452), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G472), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT72), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n435), .A2(new_n460), .A3(new_n436), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n438), .A2(new_n442), .A3(new_n459), .A4(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G217), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(G234), .B2(new_n316), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n219), .A2(G128), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n194), .A2(G119), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT24), .B(G110), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n219), .A2(G128), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n472), .B(new_n466), .C1(new_n473), .C2(KEYINPUT23), .ZN(new_n474));
  OAI22_X1  g288(.A1(new_n469), .A2(new_n471), .B1(new_n474), .B2(G110), .ZN(new_n475));
  INV_X1    g289(.A(G140), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G125), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n193), .A2(G140), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT76), .B1(new_n479), .B2(G146), .ZN(new_n480));
  XNOR2_X1  g294(.A(G125), .B(G140), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT76), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(new_n196), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT16), .ZN(new_n485));
  OR3_X1    g299(.A1(new_n193), .A2(KEYINPUT16), .A3(G140), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(G146), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n475), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n474), .A2(KEYINPUT75), .A3(G110), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT75), .B1(new_n474), .B2(G110), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n469), .A2(new_n471), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n485), .A2(G146), .A3(new_n486), .ZN(new_n493));
  AOI21_X1  g307(.A(G146), .B1(new_n485), .B2(new_n486), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n488), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT22), .B(G137), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  OAI221_X1 g315(.A(new_n492), .B1(new_n493), .B2(new_n494), .C1(new_n489), .C2(new_n490), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(new_n488), .A3(new_n499), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n503), .A3(new_n316), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT77), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n505), .A2(KEYINPUT25), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n506), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n501), .A2(new_n503), .A3(new_n316), .A4(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n465), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n501), .A2(new_n503), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n511), .A2(G902), .A3(new_n464), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n514));
  XNOR2_X1  g328(.A(G113), .B(G122), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(new_n251), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT19), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n479), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n481), .A2(KEYINPUT19), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(KEYINPUT91), .B(new_n487), .C1(new_n520), .C2(G146), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n412), .A2(new_n189), .A3(G214), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n198), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n412), .A2(new_n189), .A3(G143), .A4(G214), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G131), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n357), .A3(new_n524), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT91), .ZN(new_n529));
  AOI21_X1  g343(.A(G146), .B1(new_n518), .B2(new_n519), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n529), .B1(new_n530), .B2(new_n493), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n521), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n484), .B1(new_n196), .B2(new_n481), .ZN(new_n533));
  INV_X1    g347(.A(new_n525), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n534), .A2(KEYINPUT90), .B1(KEYINPUT18), .B2(G131), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT90), .ZN(new_n536));
  NAND2_X1  g350(.A1(KEYINPUT18), .A2(G131), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n525), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n533), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n516), .B1(new_n532), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n493), .A2(new_n494), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n525), .A2(KEYINPUT17), .A3(G131), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n541), .B(new_n542), .C1(new_n528), .C2(KEYINPUT17), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n539), .A2(new_n543), .A3(new_n516), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(G475), .A2(G902), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  OAI211_X1 g361(.A(KEYINPUT92), .B(new_n514), .C1(new_n545), .C2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n516), .B1(new_n539), .B2(new_n543), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n316), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G475), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(G234), .A2(G237), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(G952), .A3(new_n189), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(G902), .A3(G953), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT21), .B(G898), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G478), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(KEYINPUT15), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G122), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G116), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT93), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n224), .A2(G122), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n567), .B1(KEYINPUT14), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(KEYINPUT14), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT95), .ZN(new_n571));
  OAI21_X1  g385(.A(G107), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n567), .A2(new_n253), .A3(new_n568), .ZN(new_n573));
  XNOR2_X1  g387(.A(G128), .B(G143), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(new_n345), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n567), .A2(new_n568), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(G107), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n253), .B1(new_n567), .B2(new_n568), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT94), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT13), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n580), .A2(new_n581), .B1(new_n194), .B2(G143), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n580), .B2(new_n581), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G134), .ZN(new_n584));
  INV_X1    g398(.A(new_n574), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n574), .B1(new_n583), .B2(G134), .ZN(new_n587));
  OAI22_X1  g401(.A1(new_n578), .A2(new_n579), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n576), .A2(new_n588), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n330), .A2(new_n463), .A3(G953), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n576), .A2(new_n588), .A3(new_n590), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n564), .B1(new_n594), .B2(new_n316), .ZN(new_n595));
  AOI211_X1 g409(.A(G902), .B(new_n563), .C1(new_n592), .C2(new_n593), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT92), .B1(new_n545), .B2(new_n547), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT92), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n599), .B(new_n546), .C1(new_n540), .C2(new_n544), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(KEYINPUT20), .A3(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n553), .A2(new_n561), .A3(new_n597), .A4(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n389), .A2(new_n462), .A3(new_n513), .A4(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n606), .B(new_n187), .C1(new_n302), .C2(new_n317), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n607), .A2(new_n329), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n606), .B1(new_n302), .B2(new_n317), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n294), .B1(new_n324), .B2(new_n218), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n324), .A2(new_n218), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n301), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n215), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(KEYINPUT98), .A3(new_n319), .ZN(new_n614));
  INV_X1    g428(.A(new_n187), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n609), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n601), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n552), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n562), .A2(G902), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n592), .A2(new_n620), .A3(new_n593), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n620), .B1(new_n592), .B2(new_n593), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT99), .B(G478), .ZN(new_n624));
  INV_X1    g438(.A(new_n594), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(G902), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n618), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n608), .A2(new_n561), .A3(new_n616), .A4(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT97), .ZN(new_n631));
  OAI21_X1  g445(.A(G472), .B1(new_n441), .B2(KEYINPUT96), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n316), .B1(new_n426), .B2(new_n434), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT96), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n631), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n441), .A2(KEYINPUT96), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n633), .A2(new_n634), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n637), .A2(new_n638), .A3(KEYINPUT97), .A4(G472), .ZN(new_n639));
  INV_X1    g453(.A(new_n513), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n386), .B2(new_n387), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n636), .A2(new_n435), .A3(new_n639), .A4(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n630), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G104), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  INV_X1    g460(.A(new_n597), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n553), .A3(new_n601), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n560), .B(KEYINPUT101), .Z(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n608), .A2(new_n616), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n642), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT35), .B(G107), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  INV_X1    g469(.A(new_n435), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n637), .A2(new_n638), .A3(G472), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n656), .B1(new_n657), .B2(new_n631), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n507), .A2(new_n509), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n464), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n502), .B2(new_n488), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n488), .B(new_n662), .C1(new_n491), .C2(new_n495), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  OAI22_X1  g479(.A1(new_n663), .A2(new_n665), .B1(KEYINPUT36), .B2(new_n500), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n464), .A2(G902), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n496), .A2(KEYINPUT102), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n500), .A2(KEYINPUT36), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n669), .A3(new_n664), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n666), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n659), .B1(new_n661), .B2(new_n671), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n666), .A2(new_n667), .A3(new_n670), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n510), .A2(new_n673), .A3(KEYINPUT103), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n602), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n389), .A2(new_n639), .A3(new_n658), .A4(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT37), .B(G110), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  OR2_X1    g493(.A1(new_n557), .A2(G900), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n555), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n647), .A2(new_n553), .A3(new_n601), .A4(new_n681), .ZN(new_n682));
  AOI211_X1 g496(.A(new_n675), .B(new_n682), .C1(new_n386), .C2(new_n387), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n462), .A2(new_n683), .A3(new_n616), .A4(new_n608), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  INV_X1    g499(.A(KEYINPUT38), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n328), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n418), .A2(new_n425), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n416), .B1(new_n428), .B2(new_n411), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n316), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G472), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n438), .A2(new_n442), .A3(new_n691), .A4(new_n461), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n618), .A2(new_n597), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n329), .A3(new_n675), .ZN(new_n695));
  OR3_X1    g509(.A1(new_n687), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n696), .A2(KEYINPUT104), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(KEYINPUT104), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT105), .B(KEYINPUT39), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n681), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n388), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(KEYINPUT40), .Z(new_n702));
  NAND3_X1  g516(.A1(new_n697), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G143), .ZN(G45));
  OAI211_X1 g518(.A(new_n627), .B(new_n681), .C1(new_n617), .C2(new_n552), .ZN(new_n705));
  AOI211_X1 g519(.A(new_n675), .B(new_n705), .C1(new_n386), .C2(new_n387), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n462), .A2(new_n706), .A3(new_n616), .A4(new_n608), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  INV_X1    g522(.A(new_n383), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n381), .A2(new_n382), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n316), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G469), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n709), .A2(new_n712), .A3(new_n331), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n462), .A2(new_n513), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n630), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT41), .B(G113), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  NOR2_X1   g531(.A1(new_n714), .A2(new_n652), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n224), .ZN(G18));
  AND2_X1   g533(.A1(new_n676), .A2(new_n713), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n462), .A2(new_n720), .A3(new_n616), .A4(new_n608), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  NAND2_X1  g536(.A1(new_n435), .A2(KEYINPUT106), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n633), .A2(G472), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n440), .A2(new_n431), .A3(new_n433), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(new_n726), .A3(new_n390), .A4(new_n316), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n723), .A2(new_n724), .A3(new_n513), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n713), .A2(new_n649), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(new_n616), .A3(new_n608), .A4(new_n694), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  OR2_X1    g546(.A1(new_n672), .A2(new_n674), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n723), .A2(new_n724), .A3(new_n733), .A4(new_n727), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n705), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n735), .A2(new_n616), .A3(new_n608), .A4(new_n713), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT107), .B(G125), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G27));
  INV_X1    g552(.A(new_n331), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n378), .B(KEYINPUT108), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n377), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n739), .B1(new_n741), .B2(new_n709), .ZN(new_n742));
  AND4_X1   g556(.A1(new_n329), .A2(new_n318), .A3(new_n327), .A4(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n459), .A2(new_n442), .A3(new_n437), .ZN(new_n745));
  INV_X1    g559(.A(new_n705), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n513), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT42), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n705), .A2(KEYINPUT42), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n462), .A2(new_n743), .A3(new_n513), .A4(new_n749), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  INV_X1    g566(.A(new_n682), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n462), .A2(new_n743), .A3(new_n513), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  NAND2_X1  g569(.A1(new_n618), .A2(new_n627), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT43), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n675), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n636), .A2(new_n435), .A3(new_n639), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n320), .B1(new_n613), .B2(new_n319), .ZN(new_n763));
  AOI211_X1 g577(.A(new_n188), .B(new_n317), .C1(new_n612), .C2(new_n215), .ZN(new_n764));
  INV_X1    g578(.A(new_n329), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n758), .A2(KEYINPUT44), .A3(new_n759), .ZN(new_n767));
  INV_X1    g581(.A(G469), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n372), .A2(new_n376), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n770), .B2(new_n769), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT46), .B1(new_n772), .B2(new_n740), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n383), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n740), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n739), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n700), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n762), .A2(new_n766), .A3(new_n767), .A4(new_n778), .ZN(new_n779));
  XOR2_X1   g593(.A(KEYINPUT109), .B(G137), .Z(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(G39));
  NAND2_X1  g595(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g597(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n784));
  OAI21_X1  g598(.A(new_n783), .B1(new_n776), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n766), .A2(new_n640), .A3(new_n746), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n786), .A2(new_n462), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT111), .Z(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  NAND2_X1  g604(.A1(new_n709), .A2(new_n712), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT112), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT49), .Z(new_n793));
  NOR4_X1   g607(.A1(new_n756), .A2(new_n640), .A3(new_n765), .A4(new_n739), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n793), .A2(new_n687), .A3(new_n693), .A4(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n731), .B(new_n721), .C1(new_n652), .C2(new_n714), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n462), .A2(new_n513), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n765), .B1(new_n318), .B2(new_n327), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n388), .A3(new_n603), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n388), .A3(new_n676), .ZN(new_n802));
  OAI22_X1  g616(.A1(new_n799), .A2(new_n801), .B1(new_n759), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n715), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n648), .A2(KEYINPUT113), .A3(new_n650), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n805), .B(new_n329), .C1(new_n763), .C2(new_n764), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n648), .A2(KEYINPUT113), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n629), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n800), .B2(new_n649), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n808), .A2(new_n642), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n798), .A2(new_n804), .A3(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n553), .A2(new_n597), .A3(new_n601), .A4(new_n681), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n814), .B(new_n675), .C1(new_n386), .C2(new_n387), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n462), .A2(new_n766), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n735), .A2(new_n743), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n754), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT114), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n754), .A2(new_n820), .A3(new_n816), .A4(new_n817), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n751), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n796), .B1(new_n813), .B2(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n604), .B(new_n677), .C1(new_n630), .C2(new_n714), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n824), .A2(new_n797), .A3(new_n811), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n821), .A2(new_n748), .A3(new_n750), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n825), .A2(KEYINPUT115), .A3(new_n819), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n736), .A2(new_n684), .A3(new_n707), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n661), .A2(new_n742), .A3(new_n671), .A4(new_n681), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n692), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n608), .A2(new_n616), .A3(new_n694), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n828), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n608), .A2(new_n616), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n835), .B(new_n462), .C1(new_n683), .C2(new_n706), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n831), .A2(new_n832), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n837), .A3(KEYINPUT52), .A4(new_n736), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n823), .A2(new_n827), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n811), .A2(new_n803), .A3(new_n715), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n826), .A2(new_n845), .A3(new_n798), .A4(new_n819), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n846), .A2(new_n839), .A3(new_n842), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n843), .A2(new_n844), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n839), .B1(new_n846), .B2(new_n796), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(KEYINPUT53), .A3(new_n827), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n843), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n841), .A2(new_n853), .A3(new_n842), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n850), .B1(new_n856), .B2(KEYINPUT54), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n785), .B1(new_n331), .B2(new_n792), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n757), .A2(new_n555), .A3(new_n728), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n766), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n687), .A3(new_n765), .A4(new_n713), .ZN(new_n861));
  OR3_X1    g675(.A1(new_n861), .A2(KEYINPUT117), .A3(KEYINPUT50), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n766), .A2(new_n713), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n757), .A2(new_n555), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n865), .A2(new_n734), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n513), .A2(new_n863), .A3(new_n556), .A4(new_n693), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n627), .A2(new_n617), .A3(new_n552), .ZN(new_n868));
  XOR2_X1   g682(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n869));
  AOI22_X1  g683(.A1(new_n867), .A2(new_n868), .B1(new_n861), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n860), .A2(new_n862), .A3(new_n866), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n745), .A2(new_n513), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n864), .A2(new_n875), .A3(new_n863), .ZN(new_n876));
  XOR2_X1   g690(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n877));
  OAI211_X1 g691(.A(G952), .B(new_n189), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n867), .A2(new_n629), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT48), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n876), .A2(KEYINPUT118), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n859), .A2(new_n835), .A3(new_n713), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NOR4_X1   g697(.A1(new_n873), .A2(new_n874), .A3(new_n878), .A4(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n857), .A2(KEYINPUT119), .A3(new_n884), .ZN(new_n885));
  OR2_X1    g699(.A1(G952), .A2(G953), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT119), .B1(new_n857), .B2(new_n884), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n795), .B1(new_n887), .B2(new_n888), .ZN(G75));
  INV_X1    g703(.A(KEYINPUT56), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT53), .B1(new_n851), .B2(new_n827), .ZN(new_n891));
  OAI21_X1  g705(.A(G902), .B1(new_n891), .B2(new_n847), .ZN(new_n892));
  INV_X1    g706(.A(G210), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n326), .A2(new_n216), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n613), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT55), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n894), .A2(new_n897), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n189), .A2(G952), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(G51));
  OAI21_X1  g715(.A(KEYINPUT54), .B1(new_n891), .B2(new_n847), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n903), .A3(new_n849), .ZN(new_n904));
  OAI211_X1 g718(.A(KEYINPUT120), .B(KEYINPUT54), .C1(new_n891), .C2(new_n847), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n740), .B(KEYINPUT57), .Z(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n710), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n892), .A2(new_n772), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n900), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(KEYINPUT121), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n909), .B1(new_n907), .B2(new_n710), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n915), .B2(new_n900), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n913), .A2(new_n916), .ZN(G54));
  INV_X1    g731(.A(KEYINPUT122), .ZN(new_n918));
  NAND2_X1  g732(.A1(KEYINPUT58), .A2(G475), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n892), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n918), .B1(new_n920), .B2(new_n545), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n900), .B1(new_n920), .B2(new_n545), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n920), .A2(new_n918), .A3(new_n545), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(G60));
  OR2_X1    g739(.A1(new_n621), .A2(new_n622), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT59), .Z(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n904), .A2(new_n905), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n912), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n857), .A2(new_n929), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(new_n927), .ZN(G63));
  XNOR2_X1  g748(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n935));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n935), .B(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n843), .B2(new_n848), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n938), .A2(new_n670), .A3(new_n666), .ZN(new_n939));
  INV_X1    g753(.A(new_n511), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n939), .B(new_n912), .C1(new_n940), .C2(new_n938), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g758(.A(new_n559), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n189), .B1(new_n945), .B2(G224), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n813), .B2(new_n189), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n326), .B1(G898), .B2(new_n189), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT125), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n947), .B(new_n949), .ZN(G69));
  AOI21_X1  g764(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n402), .A2(new_n404), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(new_n520), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT126), .Z(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n789), .A2(new_n779), .ZN(new_n957));
  INV_X1    g771(.A(new_n629), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n701), .B1(new_n958), .B2(new_n648), .ZN(new_n959));
  AND4_X1   g773(.A1(new_n462), .A2(new_n959), .A3(new_n513), .A4(new_n766), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n829), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n703), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n961), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n956), .B1(new_n966), .B2(new_n189), .ZN(new_n967));
  AND2_X1   g781(.A1(G900), .A2(G953), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n778), .A2(new_n835), .A3(new_n694), .A4(new_n875), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n751), .A2(new_n969), .A3(new_n754), .A4(new_n962), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n957), .A2(new_n970), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n968), .B(new_n954), .C1(new_n971), .C2(new_n189), .ZN(new_n972));
  OAI21_X1  g786(.A(KEYINPUT127), .B1(new_n967), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n967), .A2(new_n972), .A3(KEYINPUT127), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n952), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n975), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n977), .A2(new_n951), .A3(new_n973), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(G72));
  NAND2_X1  g793(.A1(G472), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT63), .Z(new_n981));
  INV_X1    g795(.A(new_n454), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n982), .A2(new_n416), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n856), .B(new_n981), .C1(new_n688), .C2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n981), .B1(new_n966), .B2(new_n813), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n985), .A2(new_n416), .A3(new_n454), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n971), .A2(new_n825), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n981), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(new_n422), .A3(new_n982), .ZN(new_n989));
  AND4_X1   g803(.A1(new_n912), .A2(new_n984), .A3(new_n986), .A4(new_n989), .ZN(G57));
endmodule


