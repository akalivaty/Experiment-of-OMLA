

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735;

  INV_X1 U369 ( .A(n406), .ZN(n529) );
  NOR2_X1 U370 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U371 ( .A(n383), .B(KEYINPUT110), .ZN(n537) );
  AND2_X2 U372 ( .A1(n380), .A2(n377), .ZN(n376) );
  NOR2_X2 U373 ( .A1(n586), .A2(n585), .ZN(n588) );
  NOR2_X1 U374 ( .A1(n735), .A2(n731), .ZN(n540) );
  XNOR2_X1 U375 ( .A(n355), .B(n354), .ZN(n735) );
  XNOR2_X2 U376 ( .A(n400), .B(n350), .ZN(n382) );
  XNOR2_X2 U377 ( .A(n723), .B(G146), .ZN(n437) );
  XNOR2_X2 U378 ( .A(n457), .B(n456), .ZN(n662) );
  XNOR2_X2 U379 ( .A(n474), .B(n422), .ZN(n723) );
  XNOR2_X2 U380 ( .A(n529), .B(KEYINPUT38), .ZN(n650) );
  OR2_X1 U381 ( .A1(n551), .A2(n550), .ZN(n373) );
  INV_X4 U382 ( .A(G128), .ZN(n356) );
  AND2_X2 U383 ( .A1(n692), .A2(n691), .ZN(n702) );
  NAND2_X1 U384 ( .A1(n371), .A2(n351), .ZN(n692) );
  NAND2_X1 U385 ( .A1(n373), .A2(n372), .ZN(n371) );
  XNOR2_X1 U386 ( .A(n570), .B(n569), .ZN(n599) );
  XNOR2_X1 U387 ( .A(n409), .B(n519), .ZN(n530) );
  XNOR2_X1 U388 ( .A(n384), .B(KEYINPUT1), .ZN(n552) );
  OR2_X1 U389 ( .A1(n687), .A2(G902), .ZN(n430) );
  INV_X2 U390 ( .A(G953), .ZN(n388) );
  XNOR2_X1 U391 ( .A(G122), .B(G104), .ZN(n491) );
  INV_X1 U392 ( .A(G902), .ZN(n483) );
  XNOR2_X1 U393 ( .A(G137), .B(G140), .ZN(n440) );
  XNOR2_X1 U394 ( .A(n428), .B(G101), .ZN(n432) );
  INV_X1 U395 ( .A(KEYINPUT65), .ZN(n428) );
  XNOR2_X1 U396 ( .A(n455), .B(n454), .ZN(n456) );
  INV_X1 U397 ( .A(KEYINPUT25), .ZN(n454) );
  XNOR2_X1 U398 ( .A(n432), .B(G110), .ZN(n475) );
  XNOR2_X1 U399 ( .A(KEYINPUT70), .B(KEYINPUT16), .ZN(n477) );
  NAND2_X1 U400 ( .A1(n530), .A2(n650), .ZN(n353) );
  NOR2_X1 U401 ( .A1(n571), .A2(n580), .ZN(n572) );
  XNOR2_X1 U402 ( .A(n361), .B(n360), .ZN(n571) );
  INV_X1 U403 ( .A(KEYINPUT104), .ZN(n360) );
  INV_X1 U404 ( .A(n627), .ZN(n368) );
  XNOR2_X1 U405 ( .A(KEYINPUT15), .B(G902), .ZN(n607) );
  XNOR2_X1 U406 ( .A(G131), .B(G134), .ZN(n422) );
  XNOR2_X1 U407 ( .A(n478), .B(G107), .ZN(n502) );
  INV_X1 U408 ( .A(G116), .ZN(n478) );
  NAND2_X2 U409 ( .A1(n376), .A2(n374), .ZN(n605) );
  NAND2_X1 U410 ( .A1(n375), .A2(KEYINPUT84), .ZN(n374) );
  XNOR2_X1 U411 ( .A(G119), .B(G110), .ZN(n441) );
  XNOR2_X1 U412 ( .A(n492), .B(n440), .ZN(n722) );
  XNOR2_X1 U413 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n447) );
  XNOR2_X1 U414 ( .A(KEYINPUT99), .B(KEYINPUT12), .ZN(n487) );
  XNOR2_X1 U415 ( .A(n490), .B(n397), .ZN(n396) );
  XNOR2_X1 U416 ( .A(n491), .B(KEYINPUT98), .ZN(n397) );
  XNOR2_X1 U417 ( .A(G131), .B(G143), .ZN(n493) );
  XOR2_X1 U418 ( .A(G140), .B(G113), .Z(n494) );
  XNOR2_X1 U419 ( .A(n473), .B(KEYINPUT10), .ZN(n492) );
  XOR2_X1 U420 ( .A(KEYINPUT89), .B(KEYINPUT77), .Z(n424) );
  XNOR2_X1 U421 ( .A(G107), .B(G104), .ZN(n423) );
  XNOR2_X1 U422 ( .A(n426), .B(n440), .ZN(n362) );
  NAND2_X1 U423 ( .A1(n546), .A2(n395), .ZN(n394) );
  NAND2_X1 U424 ( .A1(n666), .A2(n392), .ZN(n391) );
  NAND2_X1 U425 ( .A1(n637), .A2(n649), .ZN(n399) );
  INV_X1 U426 ( .A(KEYINPUT76), .ZN(n519) );
  NOR2_X1 U427 ( .A1(n579), .A2(n518), .ZN(n412) );
  BUF_X1 U428 ( .A(n552), .Z(n666) );
  INV_X1 U429 ( .A(G472), .ZN(n438) );
  NOR2_X1 U430 ( .A1(n618), .A2(G902), .ZN(n439) );
  XNOR2_X1 U431 ( .A(n348), .B(n498), .ZN(n532) );
  XNOR2_X1 U432 ( .A(n404), .B(n562), .ZN(n580) );
  XNOR2_X1 U433 ( .A(n482), .B(n708), .ZN(n610) );
  XNOR2_X1 U434 ( .A(n403), .B(n476), .ZN(n482) );
  XNOR2_X1 U435 ( .A(n474), .B(n475), .ZN(n403) );
  AND2_X1 U436 ( .A1(n613), .A2(G953), .ZN(n707) );
  INV_X1 U437 ( .A(KEYINPUT74), .ZN(n401) );
  INV_X1 U438 ( .A(KEYINPUT85), .ZN(n587) );
  XNOR2_X1 U439 ( .A(n432), .B(n433), .ZN(n418) );
  XNOR2_X1 U440 ( .A(n347), .B(n434), .ZN(n416) );
  INV_X1 U441 ( .A(KEYINPUT73), .ZN(n434) );
  NOR2_X1 U442 ( .A1(n379), .A2(n378), .ZN(n377) );
  INV_X1 U443 ( .A(n643), .ZN(n378) );
  NOR2_X1 U444 ( .A1(n414), .A2(n413), .ZN(n379) );
  XNOR2_X1 U445 ( .A(KEYINPUT23), .B(KEYINPUT80), .ZN(n443) );
  XNOR2_X1 U446 ( .A(n386), .B(KEYINPUT75), .ZN(n486) );
  NAND2_X1 U447 ( .A1(n388), .A2(n387), .ZN(n386) );
  XNOR2_X1 U448 ( .A(n431), .B(G113), .ZN(n480) );
  XNOR2_X1 U449 ( .A(KEYINPUT3), .B(G119), .ZN(n431) );
  INV_X1 U450 ( .A(KEYINPUT30), .ZN(n411) );
  XNOR2_X1 U451 ( .A(n366), .B(n349), .ZN(n406) );
  NAND2_X1 U452 ( .A1(n610), .A2(n607), .ZN(n366) );
  XNOR2_X1 U453 ( .A(n437), .B(n436), .ZN(n618) );
  XNOR2_X1 U454 ( .A(n417), .B(n415), .ZN(n436) );
  XNOR2_X1 U455 ( .A(n480), .B(n416), .ZN(n415) );
  XNOR2_X1 U456 ( .A(n435), .B(n418), .ZN(n417) );
  XNOR2_X1 U457 ( .A(G122), .B(G134), .ZN(n501) );
  INV_X1 U458 ( .A(KEYINPUT66), .ZN(n420) );
  XNOR2_X1 U459 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n471) );
  XNOR2_X1 U460 ( .A(n575), .B(KEYINPUT106), .ZN(n554) );
  NAND2_X1 U461 ( .A1(G234), .A2(G237), .ZN(n461) );
  XNOR2_X1 U462 ( .A(n534), .B(KEYINPUT41), .ZN(n535) );
  XNOR2_X1 U463 ( .A(n405), .B(KEYINPUT19), .ZN(n561) );
  NAND2_X1 U464 ( .A1(n406), .A2(n649), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n469), .B(KEYINPUT28), .ZN(n385) );
  NOR2_X1 U466 ( .A1(n670), .A2(n513), .ZN(n469) );
  XNOR2_X1 U467 ( .A(n618), .B(KEYINPUT62), .ZN(n619) );
  XNOR2_X1 U468 ( .A(n605), .B(n724), .ZN(n725) );
  XNOR2_X1 U469 ( .A(n722), .B(G128), .ZN(n452) );
  XNOR2_X1 U470 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U471 ( .A(n359), .B(n398), .ZN(n695) );
  XNOR2_X1 U472 ( .A(n396), .B(n495), .ZN(n359) );
  XNOR2_X1 U473 ( .A(n437), .B(n402), .ZN(n687) );
  XNOR2_X1 U474 ( .A(n427), .B(n475), .ZN(n402) );
  XNOR2_X1 U475 ( .A(n425), .B(n362), .ZN(n427) );
  INV_X1 U476 ( .A(KEYINPUT40), .ZN(n354) );
  NAND2_X1 U477 ( .A1(n390), .A2(n389), .ZN(n642) );
  NOR2_X1 U478 ( .A1(n543), .A2(n394), .ZN(n393) );
  BUF_X1 U479 ( .A(n599), .Z(n617) );
  NOR2_X1 U480 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U481 ( .A(n522), .B(n521), .ZN(n732) );
  AND2_X1 U482 ( .A1(n532), .A2(n511), .ZN(n637) );
  AND2_X1 U483 ( .A1(n369), .A2(n670), .ZN(n627) );
  XNOR2_X1 U484 ( .A(n610), .B(n609), .ZN(n611) );
  NOR2_X1 U485 ( .A1(n532), .A2(n511), .ZN(n346) );
  INV_X1 U486 ( .A(n616), .ZN(n414) );
  XOR2_X1 U487 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n347) );
  NOR2_X1 U488 ( .A1(n695), .A2(G902), .ZN(n348) );
  XNOR2_X1 U489 ( .A(n510), .B(n509), .ZN(n531) );
  XNOR2_X1 U490 ( .A(n363), .B(n604), .ZN(n713) );
  INV_X1 U491 ( .A(n713), .ZN(n372) );
  AND2_X1 U492 ( .A1(n484), .A2(G210), .ZN(n349) );
  INV_X1 U493 ( .A(G237), .ZN(n387) );
  XNOR2_X1 U494 ( .A(KEYINPUT67), .B(KEYINPUT48), .ZN(n350) );
  INV_X1 U495 ( .A(KEYINPUT84), .ZN(n413) );
  NOR2_X2 U496 ( .A1(n662), .A2(n661), .ZN(n665) );
  NAND2_X1 U497 ( .A1(n352), .A2(KEYINPUT2), .ZN(n351) );
  XNOR2_X2 U498 ( .A(n430), .B(n429), .ZN(n384) );
  INV_X1 U499 ( .A(n644), .ZN(n352) );
  NOR2_X1 U500 ( .A1(n616), .A2(KEYINPUT84), .ZN(n381) );
  XNOR2_X2 U501 ( .A(n353), .B(KEYINPUT39), .ZN(n548) );
  XNOR2_X1 U502 ( .A(n555), .B(KEYINPUT33), .ZN(n658) );
  NAND2_X1 U503 ( .A1(n548), .A2(n637), .ZN(n355) );
  XNOR2_X2 U504 ( .A(n499), .B(n421), .ZN(n474) );
  XNOR2_X2 U505 ( .A(n356), .B(G143), .ZN(n499) );
  NAND2_X1 U506 ( .A1(n357), .A2(n603), .ZN(n364) );
  NAND2_X1 U507 ( .A1(n358), .A2(n600), .ZN(n357) );
  INV_X1 U508 ( .A(n602), .ZN(n358) );
  NOR2_X1 U509 ( .A1(n652), .A2(n661), .ZN(n361) );
  NOR2_X1 U510 ( .A1(G902), .A2(n703), .ZN(n457) );
  NOR2_X1 U511 ( .A1(n658), .A2(n580), .ZN(n566) );
  XNOR2_X1 U512 ( .A(n517), .B(n411), .ZN(n410) );
  NOR2_X1 U513 ( .A1(n713), .A2(n605), .ZN(n644) );
  NAND2_X1 U514 ( .A1(n365), .A2(n364), .ZN(n363) );
  XNOR2_X1 U515 ( .A(n588), .B(n587), .ZN(n365) );
  NAND2_X1 U516 ( .A1(n367), .A2(n582), .ZN(n583) );
  NAND2_X1 U517 ( .A1(n370), .A2(n368), .ZN(n367) );
  XNOR2_X1 U518 ( .A(n581), .B(KEYINPUT94), .ZN(n369) );
  INV_X1 U519 ( .A(n639), .ZN(n370) );
  NAND2_X1 U520 ( .A1(n382), .A2(n381), .ZN(n380) );
  INV_X1 U521 ( .A(n382), .ZN(n375) );
  NOR2_X1 U522 ( .A1(n676), .A2(n537), .ZN(n538) );
  NAND2_X1 U523 ( .A1(n385), .A2(n384), .ZN(n383) );
  AND2_X2 U524 ( .A1(n605), .A2(n401), .ZN(n550) );
  NAND2_X1 U525 ( .A1(n543), .A2(n515), .ZN(n389) );
  NOR2_X1 U526 ( .A1(n393), .A2(n391), .ZN(n390) );
  NAND2_X1 U527 ( .A1(n529), .A2(n515), .ZN(n392) );
  INV_X1 U528 ( .A(n515), .ZN(n395) );
  NAND2_X1 U529 ( .A1(n516), .A2(n642), .ZN(n524) );
  XNOR2_X1 U530 ( .A(n489), .B(n492), .ZN(n398) );
  NOR2_X1 U531 ( .A1(n399), .A2(n513), .ZN(n514) );
  NAND2_X1 U532 ( .A1(n541), .A2(n542), .ZN(n400) );
  NAND2_X1 U533 ( .A1(n561), .A2(n560), .ZN(n404) );
  NOR2_X1 U534 ( .A1(n407), .A2(n707), .ZN(n697) );
  XNOR2_X1 U535 ( .A(n408), .B(n696), .ZN(n407) );
  NAND2_X1 U536 ( .A1(n692), .A2(n693), .ZN(n408) );
  NAND2_X1 U537 ( .A1(n412), .A2(n410), .ZN(n409) );
  XOR2_X1 U538 ( .A(n527), .B(KEYINPUT71), .Z(n419) );
  XNOR2_X1 U539 ( .A(n732), .B(KEYINPUT79), .ZN(n523) );
  AND2_X1 U540 ( .A1(n528), .A2(n419), .ZN(n542) );
  INV_X1 U541 ( .A(n573), .ZN(n553) );
  NAND2_X1 U542 ( .A1(n552), .A2(n665), .ZN(n575) );
  INV_X1 U543 ( .A(KEYINPUT111), .ZN(n534) );
  XNOR2_X1 U544 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U545 ( .A(n695), .B(n694), .ZN(n696) );
  INV_X1 U546 ( .A(KEYINPUT109), .ZN(n521) );
  XNOR2_X1 U547 ( .A(n420), .B(KEYINPUT4), .ZN(n421) );
  XNOR2_X1 U548 ( .A(n424), .B(n423), .ZN(n425) );
  NAND2_X1 U549 ( .A1(G227), .A2(n388), .ZN(n426) );
  XNOR2_X1 U550 ( .A(KEYINPUT68), .B(G469), .ZN(n429) );
  XNOR2_X1 U551 ( .A(G137), .B(G116), .ZN(n433) );
  NAND2_X1 U552 ( .A1(G210), .A2(n486), .ZN(n435) );
  XNOR2_X2 U553 ( .A(n439), .B(n438), .ZN(n592) );
  INV_X1 U554 ( .A(n592), .ZN(n670) );
  XNOR2_X2 U555 ( .A(G146), .B(G125), .ZN(n473) );
  XOR2_X1 U556 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n442) );
  XNOR2_X1 U557 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U558 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n444) );
  XNOR2_X1 U559 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U560 ( .A(n446), .B(n445), .Z(n450) );
  NAND2_X1 U561 ( .A1(n388), .A2(G234), .ZN(n448) );
  XNOR2_X1 U562 ( .A(n448), .B(n447), .ZN(n500) );
  NAND2_X1 U563 ( .A1(n500), .A2(G221), .ZN(n449) );
  XNOR2_X1 U564 ( .A(n451), .B(n452), .ZN(n703) );
  NAND2_X1 U565 ( .A1(G234), .A2(n607), .ZN(n453) );
  XNOR2_X1 U566 ( .A(KEYINPUT20), .B(n453), .ZN(n458) );
  NAND2_X1 U567 ( .A1(n458), .A2(G217), .ZN(n455) );
  NAND2_X1 U568 ( .A1(n458), .A2(G221), .ZN(n459) );
  XNOR2_X1 U569 ( .A(n459), .B(KEYINPUT21), .ZN(n460) );
  XOR2_X1 U570 ( .A(KEYINPUT93), .B(n460), .Z(n661) );
  XNOR2_X1 U571 ( .A(n461), .B(KEYINPUT14), .ZN(n463) );
  NAND2_X1 U572 ( .A1(n463), .A2(G952), .ZN(n462) );
  XOR2_X1 U573 ( .A(KEYINPUT87), .B(n462), .Z(n682) );
  NOR2_X1 U574 ( .A1(n682), .A2(G953), .ZN(n556) );
  NAND2_X1 U575 ( .A1(G902), .A2(n463), .ZN(n464) );
  XOR2_X1 U576 ( .A(KEYINPUT88), .B(n464), .Z(n465) );
  NAND2_X1 U577 ( .A1(G953), .A2(n465), .ZN(n557) );
  NOR2_X1 U578 ( .A1(G900), .A2(n557), .ZN(n466) );
  XOR2_X1 U579 ( .A(KEYINPUT107), .B(n466), .Z(n467) );
  NOR2_X1 U580 ( .A1(n556), .A2(n467), .ZN(n518) );
  NOR2_X1 U581 ( .A1(n661), .A2(n518), .ZN(n468) );
  NAND2_X1 U582 ( .A1(n662), .A2(n468), .ZN(n513) );
  NAND2_X1 U583 ( .A1(n388), .A2(G224), .ZN(n470) );
  XNOR2_X1 U584 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U585 ( .A(n473), .B(n472), .ZN(n476) );
  XNOR2_X1 U586 ( .A(n491), .B(n477), .ZN(n479) );
  XNOR2_X1 U587 ( .A(n479), .B(n502), .ZN(n481) );
  XNOR2_X1 U588 ( .A(n481), .B(n480), .ZN(n708) );
  NAND2_X1 U589 ( .A1(n483), .A2(n387), .ZN(n484) );
  NAND2_X1 U590 ( .A1(n484), .A2(G214), .ZN(n649) );
  INV_X1 U591 ( .A(n561), .ZN(n485) );
  NOR2_X2 U592 ( .A1(n537), .A2(n485), .ZN(n635) );
  NAND2_X1 U593 ( .A1(G214), .A2(n486), .ZN(n490) );
  XOR2_X1 U594 ( .A(KEYINPUT100), .B(KEYINPUT11), .Z(n488) );
  XNOR2_X1 U595 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U596 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U597 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n497) );
  INV_X1 U598 ( .A(G475), .ZN(n496) );
  XNOR2_X1 U599 ( .A(n499), .B(KEYINPUT9), .ZN(n508) );
  NAND2_X1 U600 ( .A1(n500), .A2(G217), .ZN(n506) );
  XNOR2_X1 U601 ( .A(KEYINPUT102), .B(KEYINPUT7), .ZN(n504) );
  XNOR2_X1 U602 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U603 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U604 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U605 ( .A(n508), .B(n507), .ZN(n698) );
  NOR2_X1 U606 ( .A1(G902), .A2(n698), .ZN(n510) );
  INV_X1 U607 ( .A(G478), .ZN(n509) );
  INV_X1 U608 ( .A(n531), .ZN(n511) );
  NOR2_X1 U609 ( .A1(n637), .A2(n346), .ZN(n654) );
  INV_X1 U610 ( .A(n654), .ZN(n582) );
  NAND2_X1 U611 ( .A1(n635), .A2(n582), .ZN(n512) );
  NAND2_X1 U612 ( .A1(n512), .A2(KEYINPUT47), .ZN(n516) );
  XOR2_X1 U613 ( .A(KEYINPUT6), .B(n592), .Z(n573) );
  NAND2_X1 U614 ( .A1(n573), .A2(n514), .ZN(n543) );
  XOR2_X1 U615 ( .A(KEYINPUT113), .B(KEYINPUT36), .Z(n515) );
  NAND2_X1 U616 ( .A1(n592), .A2(n649), .ZN(n517) );
  NAND2_X1 U617 ( .A1(n665), .A2(n384), .ZN(n579) );
  AND2_X1 U618 ( .A1(n532), .A2(n531), .ZN(n567) );
  INV_X1 U619 ( .A(n529), .ZN(n546) );
  AND2_X1 U620 ( .A1(n567), .A2(n546), .ZN(n520) );
  NAND2_X1 U621 ( .A1(n530), .A2(n520), .ZN(n522) );
  NOR2_X1 U622 ( .A1(n524), .A2(n523), .ZN(n528) );
  NOR2_X1 U623 ( .A1(n654), .A2(KEYINPUT47), .ZN(n525) );
  XNOR2_X1 U624 ( .A(KEYINPUT72), .B(n525), .ZN(n526) );
  NAND2_X1 U625 ( .A1(n635), .A2(n526), .ZN(n527) );
  XNOR2_X1 U626 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n539) );
  NOR2_X1 U627 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U628 ( .A(n533), .B(KEYINPUT103), .ZN(n652) );
  NAND2_X1 U629 ( .A1(n650), .A2(n649), .ZN(n653) );
  NOR2_X1 U630 ( .A1(n652), .A2(n653), .ZN(n536) );
  XNOR2_X1 U631 ( .A(n536), .B(n535), .ZN(n676) );
  XNOR2_X1 U632 ( .A(n539), .B(n538), .ZN(n731) );
  XNOR2_X1 U633 ( .A(n540), .B(KEYINPUT46), .ZN(n541) );
  NOR2_X1 U634 ( .A1(n666), .A2(n543), .ZN(n545) );
  XNOR2_X1 U635 ( .A(KEYINPUT43), .B(KEYINPUT108), .ZN(n544) );
  XNOR2_X1 U636 ( .A(n545), .B(n544), .ZN(n547) );
  NOR2_X1 U637 ( .A1(n547), .A2(n546), .ZN(n616) );
  NAND2_X1 U638 ( .A1(n548), .A2(n346), .ZN(n643) );
  INV_X1 U639 ( .A(KEYINPUT2), .ZN(n606) );
  NAND2_X1 U640 ( .A1(n606), .A2(KEYINPUT74), .ZN(n549) );
  NOR2_X1 U641 ( .A1(n605), .A2(n549), .ZN(n551) );
  INV_X1 U642 ( .A(n556), .ZN(n559) );
  OR2_X1 U643 ( .A1(n557), .A2(G898), .ZN(n558) );
  NAND2_X1 U644 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U645 ( .A(KEYINPUT64), .B(KEYINPUT0), .ZN(n562) );
  XNOR2_X1 U646 ( .A(KEYINPUT78), .B(KEYINPUT34), .ZN(n564) );
  INV_X1 U647 ( .A(KEYINPUT69), .ZN(n563) );
  XNOR2_X1 U648 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U649 ( .A(n566), .B(n565), .ZN(n568) );
  NAND2_X1 U650 ( .A1(n568), .A2(n567), .ZN(n570) );
  XNOR2_X1 U651 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n569) );
  INV_X1 U652 ( .A(KEYINPUT44), .ZN(n600) );
  NOR2_X1 U653 ( .A1(n599), .A2(n600), .ZN(n586) );
  XNOR2_X1 U654 ( .A(n572), .B(KEYINPUT22), .ZN(n589) );
  NAND2_X1 U655 ( .A1(n589), .A2(n553), .ZN(n597) );
  INV_X1 U656 ( .A(n662), .ZN(n594) );
  INV_X1 U657 ( .A(n666), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n574) );
  NOR2_X1 U659 ( .A1(n597), .A2(n574), .ZN(n624) );
  INV_X1 U660 ( .A(n624), .ZN(n584) );
  NOR2_X1 U661 ( .A1(n670), .A2(n575), .ZN(n576) );
  XOR2_X1 U662 ( .A(KEYINPUT96), .B(n576), .Z(n673) );
  NOR2_X1 U663 ( .A1(n673), .A2(n580), .ZN(n578) );
  XNOR2_X1 U664 ( .A(KEYINPUT31), .B(KEYINPUT97), .ZN(n577) );
  XNOR2_X1 U665 ( .A(n578), .B(n577), .ZN(n639) );
  NOR2_X1 U666 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U667 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U668 ( .A1(n666), .A2(n594), .ZN(n590) );
  NAND2_X1 U669 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U670 ( .A1(n592), .A2(n591), .ZN(n631) );
  NOR2_X1 U671 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U672 ( .A(n595), .B(KEYINPUT105), .ZN(n596) );
  XNOR2_X1 U673 ( .A(KEYINPUT32), .B(n598), .ZN(n733) );
  NOR2_X1 U674 ( .A1(n631), .A2(n733), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n617), .A2(n600), .ZN(n601) );
  NAND2_X1 U676 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U677 ( .A(KEYINPUT82), .B(KEYINPUT45), .Z(n604) );
  INV_X1 U678 ( .A(n607), .ZN(n691) );
  NAND2_X1 U679 ( .A1(n702), .A2(G210), .ZN(n612) );
  XOR2_X1 U680 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n608) );
  XNOR2_X1 U681 ( .A(n608), .B(KEYINPUT55), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n612), .B(n611), .ZN(n614) );
  INV_X1 U683 ( .A(G952), .ZN(n613) );
  NOR2_X1 U684 ( .A1(n614), .A2(n707), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n615), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U686 ( .A(G140), .B(n616), .Z(G42) );
  XNOR2_X1 U687 ( .A(n617), .B(G122), .ZN(G24) );
  NAND2_X1 U688 ( .A1(n702), .A2(G472), .ZN(n620) );
  XNOR2_X1 U689 ( .A(n620), .B(n619), .ZN(n621) );
  NOR2_X1 U690 ( .A1(n621), .A2(n707), .ZN(n623) );
  XOR2_X1 U691 ( .A(KEYINPUT86), .B(KEYINPUT63), .Z(n622) );
  XNOR2_X1 U692 ( .A(n623), .B(n622), .ZN(G57) );
  XOR2_X1 U693 ( .A(G101), .B(n624), .Z(G3) );
  NAND2_X1 U694 ( .A1(n627), .A2(n637), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n625), .B(KEYINPUT114), .ZN(n626) );
  XNOR2_X1 U696 ( .A(G104), .B(n626), .ZN(G6) );
  XOR2_X1 U697 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n629) );
  NAND2_X1 U698 ( .A1(n627), .A2(n346), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U700 ( .A(G107), .B(n630), .ZN(G9) );
  XNOR2_X1 U701 ( .A(G110), .B(n631), .ZN(n632) );
  XNOR2_X1 U702 ( .A(n632), .B(KEYINPUT115), .ZN(G12) );
  XOR2_X1 U703 ( .A(G128), .B(KEYINPUT29), .Z(n634) );
  NAND2_X1 U704 ( .A1(n635), .A2(n346), .ZN(n633) );
  XNOR2_X1 U705 ( .A(n634), .B(n633), .ZN(G30) );
  NAND2_X1 U706 ( .A1(n635), .A2(n637), .ZN(n636) );
  XNOR2_X1 U707 ( .A(n636), .B(G146), .ZN(G48) );
  NAND2_X1 U708 ( .A1(n639), .A2(n637), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n638), .B(G113), .ZN(G15) );
  NAND2_X1 U710 ( .A1(n639), .A2(n346), .ZN(n640) );
  XNOR2_X1 U711 ( .A(n640), .B(G116), .ZN(G18) );
  XOR2_X1 U712 ( .A(G125), .B(KEYINPUT37), .Z(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n641), .ZN(G27) );
  XNOR2_X1 U714 ( .A(G134), .B(n643), .ZN(G36) );
  XNOR2_X1 U715 ( .A(n644), .B(KEYINPUT2), .ZN(n648) );
  OR2_X1 U716 ( .A1(n676), .A2(n658), .ZN(n645) );
  XOR2_X1 U717 ( .A(KEYINPUT120), .B(n645), .Z(n646) );
  NOR2_X1 U718 ( .A1(G953), .A2(n646), .ZN(n647) );
  NAND2_X1 U719 ( .A1(n648), .A2(n647), .ZN(n684) );
  NOR2_X1 U720 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n657) );
  NOR2_X1 U722 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U723 ( .A(KEYINPUT117), .B(n655), .Z(n656) );
  NOR2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n659) );
  NOR2_X1 U725 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U726 ( .A(n660), .B(KEYINPUT118), .ZN(n678) );
  NAND2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U728 ( .A(n663), .B(KEYINPUT49), .ZN(n664) );
  XNOR2_X1 U729 ( .A(KEYINPUT116), .B(n664), .ZN(n669) );
  NOR2_X1 U730 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U731 ( .A(KEYINPUT50), .B(n667), .ZN(n668) );
  NOR2_X1 U732 ( .A1(n669), .A2(n668), .ZN(n671) );
  NAND2_X1 U733 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U734 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U735 ( .A(KEYINPUT51), .B(n674), .ZN(n675) );
  NOR2_X1 U736 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U737 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U738 ( .A(n679), .B(KEYINPUT119), .Z(n680) );
  XNOR2_X1 U739 ( .A(KEYINPUT52), .B(n680), .ZN(n681) );
  NOR2_X1 U740 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U741 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U742 ( .A(n685), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U743 ( .A1(n702), .A2(G469), .ZN(n689) );
  XOR2_X1 U744 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n686) );
  XNOR2_X1 U745 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U746 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U747 ( .A1(n707), .A2(n690), .ZN(G54) );
  AND2_X1 U748 ( .A1(G475), .A2(n691), .ZN(n693) );
  XOR2_X1 U749 ( .A(KEYINPUT59), .B(KEYINPUT122), .Z(n694) );
  XNOR2_X1 U750 ( .A(KEYINPUT60), .B(n697), .ZN(G60) );
  NAND2_X1 U751 ( .A1(n702), .A2(G478), .ZN(n700) );
  XOR2_X1 U752 ( .A(n698), .B(KEYINPUT123), .Z(n699) );
  XNOR2_X1 U753 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U754 ( .A1(n707), .A2(n701), .ZN(G63) );
  NAND2_X1 U755 ( .A1(n702), .A2(G217), .ZN(n705) );
  BUF_X1 U756 ( .A(n703), .Z(n704) );
  XNOR2_X1 U757 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U758 ( .A1(n707), .A2(n706), .ZN(G66) );
  XNOR2_X1 U759 ( .A(G101), .B(G110), .ZN(n709) );
  XOR2_X1 U760 ( .A(n709), .B(n708), .Z(n711) );
  NOR2_X1 U761 ( .A1(G898), .A2(n388), .ZN(n710) );
  NOR2_X1 U762 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U763 ( .A(KEYINPUT126), .B(n712), .ZN(n721) );
  NAND2_X1 U764 ( .A1(n372), .A2(n388), .ZN(n719) );
  XOR2_X1 U765 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n715) );
  NAND2_X1 U766 ( .A1(G224), .A2(G953), .ZN(n714) );
  XNOR2_X1 U767 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U768 ( .A(KEYINPUT124), .B(n716), .ZN(n717) );
  NAND2_X1 U769 ( .A1(n717), .A2(G898), .ZN(n718) );
  NAND2_X1 U770 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U771 ( .A(n721), .B(n720), .ZN(G69) );
  XNOR2_X1 U772 ( .A(n723), .B(n722), .ZN(n726) );
  INV_X1 U773 ( .A(n726), .ZN(n724) );
  NAND2_X1 U774 ( .A1(n725), .A2(n388), .ZN(n730) );
  XOR2_X1 U775 ( .A(G227), .B(n726), .Z(n727) );
  NAND2_X1 U776 ( .A1(n727), .A2(G900), .ZN(n728) );
  NAND2_X1 U777 ( .A1(n728), .A2(G953), .ZN(n729) );
  NAND2_X1 U778 ( .A1(n730), .A2(n729), .ZN(G72) );
  XOR2_X1 U779 ( .A(n731), .B(G137), .Z(G39) );
  XNOR2_X1 U780 ( .A(G143), .B(n732), .ZN(G45) );
  XNOR2_X1 U781 ( .A(G119), .B(KEYINPUT127), .ZN(n734) );
  XNOR2_X1 U782 ( .A(n734), .B(n733), .ZN(G21) );
  XOR2_X1 U783 ( .A(n735), .B(G131), .Z(G33) );
endmodule

