

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U555 ( .A(KEYINPUT32), .B(KEYINPUT100), .ZN(n748) );
  NAND2_X1 U556 ( .A1(n692), .A2(n805), .ZN(n741) );
  XNOR2_X1 U557 ( .A(n749), .B(n748), .ZN(n758) );
  NOR2_X1 U558 ( .A1(G651), .A2(n638), .ZN(n646) );
  XOR2_X1 U559 ( .A(KEYINPUT1), .B(n542), .Z(n653) );
  NOR2_X1 U560 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  XOR2_X2 U561 ( .A(KEYINPUT17), .B(n521), .Z(n895) );
  NAND2_X1 U562 ( .A1(n895), .A2(G137), .ZN(n523) );
  AND2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n901) );
  NAND2_X1 U564 ( .A1(n901), .A2(G113), .ZN(n522) );
  NAND2_X1 U565 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U566 ( .A(n524), .B(KEYINPUT65), .ZN(n526) );
  INV_X1 U567 ( .A(G2105), .ZN(n527) );
  NOR2_X1 U568 ( .A1(G2104), .A2(n527), .ZN(n902) );
  NAND2_X1 U569 ( .A1(G125), .A2(n902), .ZN(n525) );
  NAND2_X1 U570 ( .A1(n526), .A2(n525), .ZN(n531) );
  AND2_X1 U571 ( .A1(G2104), .A2(n527), .ZN(n528) );
  XNOR2_X1 U572 ( .A(n528), .B(KEYINPUT64), .ZN(n897) );
  NAND2_X1 U573 ( .A1(G101), .A2(n897), .ZN(n529) );
  XNOR2_X1 U574 ( .A(KEYINPUT23), .B(n529), .ZN(n530) );
  NOR2_X2 U575 ( .A1(n531), .A2(n530), .ZN(G160) );
  XOR2_X1 U576 ( .A(G2443), .B(G2446), .Z(n533) );
  XNOR2_X1 U577 ( .A(G2427), .B(G2451), .ZN(n532) );
  XNOR2_X1 U578 ( .A(n533), .B(n532), .ZN(n539) );
  XOR2_X1 U579 ( .A(G2430), .B(G2454), .Z(n535) );
  XNOR2_X1 U580 ( .A(G1341), .B(G1348), .ZN(n534) );
  XNOR2_X1 U581 ( .A(n535), .B(n534), .ZN(n537) );
  XOR2_X1 U582 ( .A(G2435), .B(G2438), .Z(n536) );
  XNOR2_X1 U583 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U584 ( .A(n539), .B(n538), .Z(n540) );
  AND2_X1 U585 ( .A1(G14), .A2(n540), .ZN(G401) );
  AND2_X1 U586 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U587 ( .A(G57), .ZN(G237) );
  INV_X1 U588 ( .A(G108), .ZN(G238) );
  INV_X1 U589 ( .A(G132), .ZN(G219) );
  INV_X1 U590 ( .A(G82), .ZN(G220) );
  XNOR2_X1 U591 ( .A(G543), .B(KEYINPUT0), .ZN(n541) );
  XNOR2_X1 U592 ( .A(n541), .B(KEYINPUT67), .ZN(n638) );
  NAND2_X1 U593 ( .A1(G52), .A2(n646), .ZN(n544) );
  INV_X1 U594 ( .A(G651), .ZN(n545) );
  NOR2_X1 U595 ( .A1(G543), .A2(n545), .ZN(n542) );
  NAND2_X1 U596 ( .A1(G64), .A2(n653), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n550) );
  NOR2_X1 U598 ( .A1(G543), .A2(G651), .ZN(n649) );
  NAND2_X1 U599 ( .A1(G90), .A2(n649), .ZN(n547) );
  NOR2_X1 U600 ( .A1(n638), .A2(n545), .ZN(n645) );
  NAND2_X1 U601 ( .A1(G77), .A2(n645), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U603 ( .A(KEYINPUT9), .B(n548), .Z(n549) );
  NOR2_X1 U604 ( .A1(n550), .A2(n549), .ZN(G171) );
  NAND2_X1 U605 ( .A1(n649), .A2(G89), .ZN(n551) );
  XNOR2_X1 U606 ( .A(n551), .B(KEYINPUT4), .ZN(n553) );
  NAND2_X1 U607 ( .A1(G76), .A2(n645), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U609 ( .A(KEYINPUT5), .B(n554), .ZN(n561) );
  XNOR2_X1 U610 ( .A(KEYINPUT6), .B(KEYINPUT72), .ZN(n559) );
  NAND2_X1 U611 ( .A1(n653), .A2(G63), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n646), .A2(G51), .ZN(n555) );
  XOR2_X1 U613 ( .A(KEYINPUT71), .B(n555), .Z(n556) );
  NAND2_X1 U614 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U615 ( .A(n559), .B(n558), .Z(n560) );
  NAND2_X1 U616 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U617 ( .A(KEYINPUT7), .B(n562), .ZN(G168) );
  XNOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .ZN(n563) );
  XNOR2_X1 U619 ( .A(n563), .B(KEYINPUT73), .ZN(G286) );
  NAND2_X1 U620 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U621 ( .A(n564), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U622 ( .A(G567), .ZN(n681) );
  NOR2_X1 U623 ( .A1(n681), .A2(G223), .ZN(n565) );
  XNOR2_X1 U624 ( .A(n565), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U625 ( .A1(n649), .A2(G81), .ZN(n566) );
  XNOR2_X1 U626 ( .A(n566), .B(KEYINPUT12), .ZN(n568) );
  NAND2_X1 U627 ( .A1(G68), .A2(n645), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U629 ( .A(n569), .B(KEYINPUT13), .ZN(n571) );
  NAND2_X1 U630 ( .A1(G43), .A2(n646), .ZN(n570) );
  NAND2_X1 U631 ( .A1(n571), .A2(n570), .ZN(n574) );
  NAND2_X1 U632 ( .A1(n653), .A2(G56), .ZN(n572) );
  XOR2_X1 U633 ( .A(KEYINPUT14), .B(n572), .Z(n573) );
  NOR2_X1 U634 ( .A1(n574), .A2(n573), .ZN(n1004) );
  NAND2_X1 U635 ( .A1(n1004), .A2(G860), .ZN(G153) );
  INV_X1 U636 ( .A(G171), .ZN(G301) );
  NAND2_X1 U637 ( .A1(G868), .A2(G301), .ZN(n585) );
  NAND2_X1 U638 ( .A1(G54), .A2(n646), .ZN(n575) );
  XNOR2_X1 U639 ( .A(n575), .B(KEYINPUT70), .ZN(n582) );
  NAND2_X1 U640 ( .A1(G92), .A2(n649), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G66), .A2(n653), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n580) );
  NAND2_X1 U643 ( .A1(G79), .A2(n645), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT69), .B(n578), .ZN(n579) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(KEYINPUT15), .B(n583), .ZN(n910) );
  INV_X1 U648 ( .A(n910), .ZN(n998) );
  INV_X1 U649 ( .A(G868), .ZN(n665) );
  NAND2_X1 U650 ( .A1(n998), .A2(n665), .ZN(n584) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(G284) );
  NAND2_X1 U652 ( .A1(G78), .A2(n645), .ZN(n587) );
  NAND2_X1 U653 ( .A1(G53), .A2(n646), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U655 ( .A1(n649), .A2(G91), .ZN(n588) );
  XOR2_X1 U656 ( .A(KEYINPUT68), .B(n588), .Z(n589) );
  NOR2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U658 ( .A1(n653), .A2(G65), .ZN(n591) );
  NAND2_X1 U659 ( .A1(n592), .A2(n591), .ZN(G299) );
  NOR2_X1 U660 ( .A1(G868), .A2(G299), .ZN(n593) );
  XNOR2_X1 U661 ( .A(n593), .B(KEYINPUT74), .ZN(n595) );
  NOR2_X1 U662 ( .A1(n665), .A2(G286), .ZN(n594) );
  NOR2_X1 U663 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U664 ( .A(KEYINPUT75), .B(n596), .Z(G297) );
  INV_X1 U665 ( .A(G860), .ZN(n620) );
  NAND2_X1 U666 ( .A1(n620), .A2(G559), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n597), .A2(n910), .ZN(n598) );
  XNOR2_X1 U668 ( .A(n598), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U669 ( .A1(n910), .A2(G868), .ZN(n599) );
  NOR2_X1 U670 ( .A1(G559), .A2(n599), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(KEYINPUT76), .ZN(n602) );
  AND2_X1 U672 ( .A1(n1004), .A2(n665), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U674 ( .A1(G111), .A2(n901), .ZN(n604) );
  NAND2_X1 U675 ( .A1(G99), .A2(n897), .ZN(n603) );
  NAND2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n605), .B(KEYINPUT77), .ZN(n607) );
  NAND2_X1 U678 ( .A1(G135), .A2(n895), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U680 ( .A1(n902), .A2(G123), .ZN(n608) );
  XOR2_X1 U681 ( .A(KEYINPUT18), .B(n608), .Z(n609) );
  NOR2_X1 U682 ( .A1(n610), .A2(n609), .ZN(n925) );
  XNOR2_X1 U683 ( .A(n925), .B(G2096), .ZN(n612) );
  INV_X1 U684 ( .A(G2100), .ZN(n611) );
  NAND2_X1 U685 ( .A1(n612), .A2(n611), .ZN(G156) );
  NAND2_X1 U686 ( .A1(G93), .A2(n649), .ZN(n614) );
  NAND2_X1 U687 ( .A1(G80), .A2(n645), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U689 ( .A1(G55), .A2(n646), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G67), .A2(n653), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  OR2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n666) );
  XNOR2_X1 U693 ( .A(n666), .B(KEYINPUT78), .ZN(n622) );
  NAND2_X1 U694 ( .A1(G559), .A2(n910), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n619), .B(n1004), .ZN(n662) );
  NAND2_X1 U696 ( .A1(n662), .A2(n620), .ZN(n621) );
  XNOR2_X1 U697 ( .A(n622), .B(n621), .ZN(G145) );
  NAND2_X1 U698 ( .A1(G50), .A2(n646), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n623), .B(KEYINPUT80), .ZN(n626) );
  NAND2_X1 U700 ( .A1(G75), .A2(n645), .ZN(n624) );
  XOR2_X1 U701 ( .A(KEYINPUT81), .B(n624), .Z(n625) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U703 ( .A1(G88), .A2(n649), .ZN(n628) );
  NAND2_X1 U704 ( .A1(G62), .A2(n653), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U706 ( .A1(n630), .A2(n629), .ZN(G166) );
  NAND2_X1 U707 ( .A1(G86), .A2(n649), .ZN(n632) );
  NAND2_X1 U708 ( .A1(G48), .A2(n646), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n645), .A2(G73), .ZN(n633) );
  XOR2_X1 U711 ( .A(KEYINPUT2), .B(n633), .Z(n634) );
  NOR2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n653), .A2(G61), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(G305) );
  NAND2_X1 U715 ( .A1(G87), .A2(n638), .ZN(n640) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U718 ( .A1(n653), .A2(n641), .ZN(n644) );
  NAND2_X1 U719 ( .A1(G49), .A2(n646), .ZN(n642) );
  XOR2_X1 U720 ( .A(KEYINPUT79), .B(n642), .Z(n643) );
  NAND2_X1 U721 ( .A1(n644), .A2(n643), .ZN(G288) );
  NAND2_X1 U722 ( .A1(G72), .A2(n645), .ZN(n648) );
  NAND2_X1 U723 ( .A1(G47), .A2(n646), .ZN(n647) );
  NAND2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U725 ( .A1(G85), .A2(n649), .ZN(n650) );
  XOR2_X1 U726 ( .A(KEYINPUT66), .B(n650), .Z(n651) );
  NOR2_X1 U727 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n653), .A2(G60), .ZN(n654) );
  NAND2_X1 U729 ( .A1(n655), .A2(n654), .ZN(G290) );
  XNOR2_X1 U730 ( .A(G166), .B(G305), .ZN(n656) );
  XNOR2_X1 U731 ( .A(n656), .B(G288), .ZN(n657) );
  XNOR2_X1 U732 ( .A(KEYINPUT19), .B(n657), .ZN(n659) );
  XNOR2_X1 U733 ( .A(G299), .B(KEYINPUT82), .ZN(n658) );
  XNOR2_X1 U734 ( .A(n659), .B(n658), .ZN(n660) );
  XOR2_X1 U735 ( .A(n666), .B(n660), .Z(n661) );
  XNOR2_X1 U736 ( .A(n661), .B(G290), .ZN(n913) );
  XNOR2_X1 U737 ( .A(n662), .B(n913), .ZN(n663) );
  NAND2_X1 U738 ( .A1(n663), .A2(G868), .ZN(n664) );
  XOR2_X1 U739 ( .A(KEYINPUT83), .B(n664), .Z(n668) );
  NAND2_X1 U740 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U741 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U744 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U745 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U746 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U748 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U749 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U750 ( .A1(G218), .A2(n674), .ZN(n675) );
  XNOR2_X1 U751 ( .A(KEYINPUT84), .B(n675), .ZN(n676) );
  NAND2_X1 U752 ( .A1(n676), .A2(G96), .ZN(n844) );
  NAND2_X1 U753 ( .A1(G2106), .A2(n844), .ZN(n677) );
  XNOR2_X1 U754 ( .A(n677), .B(KEYINPUT85), .ZN(n683) );
  NAND2_X1 U755 ( .A1(G120), .A2(G69), .ZN(n678) );
  NOR2_X1 U756 ( .A1(G237), .A2(n678), .ZN(n679) );
  XOR2_X1 U757 ( .A(KEYINPUT86), .B(n679), .Z(n680) );
  NOR2_X1 U758 ( .A1(G238), .A2(n680), .ZN(n843) );
  NOR2_X1 U759 ( .A1(n681), .A2(n843), .ZN(n682) );
  NOR2_X1 U760 ( .A1(n683), .A2(n682), .ZN(G319) );
  INV_X1 U761 ( .A(G319), .ZN(n685) );
  NAND2_X1 U762 ( .A1(G483), .A2(G661), .ZN(n684) );
  NOR2_X1 U763 ( .A1(n685), .A2(n684), .ZN(n842) );
  NAND2_X1 U764 ( .A1(n842), .A2(G36), .ZN(G176) );
  NAND2_X1 U765 ( .A1(G138), .A2(n895), .ZN(n687) );
  NAND2_X1 U766 ( .A1(G102), .A2(n897), .ZN(n686) );
  NAND2_X1 U767 ( .A1(n687), .A2(n686), .ZN(n691) );
  NAND2_X1 U768 ( .A1(G114), .A2(n901), .ZN(n689) );
  NAND2_X1 U769 ( .A1(G126), .A2(n902), .ZN(n688) );
  NAND2_X1 U770 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U771 ( .A1(n691), .A2(n690), .ZN(G164) );
  XNOR2_X1 U772 ( .A(KEYINPUT87), .B(G166), .ZN(G303) );
  NAND2_X1 U773 ( .A1(G160), .A2(G40), .ZN(n804) );
  INV_X1 U774 ( .A(n804), .ZN(n692) );
  NOR2_X1 U775 ( .A1(G164), .A2(G1384), .ZN(n805) );
  NAND2_X1 U776 ( .A1(n741), .A2(G8), .ZN(n693) );
  XNOR2_X1 U777 ( .A(n693), .B(KEYINPUT90), .ZN(n781) );
  OR2_X1 U778 ( .A1(n781), .A2(G1966), .ZN(n696) );
  NOR2_X1 U779 ( .A1(G2084), .A2(n741), .ZN(n750) );
  INV_X1 U780 ( .A(G8), .ZN(n694) );
  NOR2_X1 U781 ( .A1(n750), .A2(n694), .ZN(n695) );
  NAND2_X1 U782 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U783 ( .A(n697), .B(KEYINPUT30), .ZN(n698) );
  NOR2_X1 U784 ( .A1(G168), .A2(n698), .ZN(n699) );
  XNOR2_X1 U785 ( .A(n699), .B(KEYINPUT99), .ZN(n703) );
  XOR2_X1 U786 ( .A(G2078), .B(KEYINPUT25), .Z(n951) );
  NOR2_X1 U787 ( .A1(n951), .A2(n741), .ZN(n701) );
  INV_X1 U788 ( .A(n741), .ZN(n717) );
  NOR2_X1 U789 ( .A1(n717), .A2(G1961), .ZN(n700) );
  NOR2_X1 U790 ( .A1(n701), .A2(n700), .ZN(n735) );
  NAND2_X1 U791 ( .A1(n735), .A2(G301), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U793 ( .A(n704), .B(KEYINPUT31), .ZN(n739) );
  INV_X1 U794 ( .A(G2072), .ZN(n942) );
  NOR2_X1 U795 ( .A1(n741), .A2(n942), .ZN(n706) );
  XNOR2_X1 U796 ( .A(KEYINPUT92), .B(KEYINPUT27), .ZN(n705) );
  XNOR2_X1 U797 ( .A(n706), .B(n705), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n741), .A2(G1956), .ZN(n707) );
  AND2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U800 ( .A(KEYINPUT93), .B(n709), .ZN(n728) );
  NOR2_X1 U801 ( .A1(n728), .A2(G299), .ZN(n710) );
  XNOR2_X1 U802 ( .A(n710), .B(KEYINPUT97), .ZN(n727) );
  NAND2_X1 U803 ( .A1(G1996), .A2(n717), .ZN(n711) );
  XNOR2_X1 U804 ( .A(KEYINPUT26), .B(n711), .ZN(n716) );
  NAND2_X1 U805 ( .A1(G1341), .A2(n741), .ZN(n712) );
  XNOR2_X1 U806 ( .A(KEYINPUT95), .B(n712), .ZN(n714) );
  INV_X1 U807 ( .A(n1004), .ZN(n713) );
  NOR2_X1 U808 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U809 ( .A1(n716), .A2(n715), .ZN(n723) );
  NAND2_X1 U810 ( .A1(n723), .A2(n910), .ZN(n721) );
  NOR2_X1 U811 ( .A1(n717), .A2(G1348), .ZN(n719) );
  NOR2_X1 U812 ( .A1(G2067), .A2(n741), .ZN(n718) );
  NOR2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U815 ( .A(n722), .B(KEYINPUT96), .ZN(n725) );
  OR2_X1 U816 ( .A1(n723), .A2(n910), .ZN(n724) );
  NAND2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U818 ( .A1(n727), .A2(n726), .ZN(n732) );
  NAND2_X1 U819 ( .A1(n728), .A2(G299), .ZN(n730) );
  XNOR2_X1 U820 ( .A(KEYINPUT94), .B(KEYINPUT28), .ZN(n729) );
  XNOR2_X1 U821 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U822 ( .A1(n732), .A2(n731), .ZN(n734) );
  XOR2_X1 U823 ( .A(KEYINPUT98), .B(KEYINPUT29), .Z(n733) );
  XNOR2_X1 U824 ( .A(n734), .B(n733), .ZN(n737) );
  OR2_X1 U825 ( .A1(n735), .A2(G301), .ZN(n736) );
  NAND2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U827 ( .A1(n739), .A2(n738), .ZN(n752) );
  AND2_X1 U828 ( .A1(G286), .A2(G8), .ZN(n740) );
  NAND2_X1 U829 ( .A1(n752), .A2(n740), .ZN(n747) );
  NOR2_X1 U830 ( .A1(n781), .A2(G1971), .ZN(n743) );
  NOR2_X1 U831 ( .A1(G2090), .A2(n741), .ZN(n742) );
  NOR2_X1 U832 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U833 ( .A1(n744), .A2(G303), .ZN(n745) );
  OR2_X1 U834 ( .A1(n694), .A2(n745), .ZN(n746) );
  AND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n749) );
  NAND2_X1 U836 ( .A1(G8), .A2(n750), .ZN(n751) );
  XOR2_X1 U837 ( .A(KEYINPUT91), .B(n751), .Z(n756) );
  INV_X1 U838 ( .A(n752), .ZN(n754) );
  NOR2_X1 U839 ( .A1(n781), .A2(G1966), .ZN(n753) );
  NOR2_X1 U840 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U841 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U842 ( .A1(n758), .A2(n757), .ZN(n780) );
  NOR2_X1 U843 ( .A1(G1971), .A2(G303), .ZN(n759) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n1011) );
  NOR2_X1 U845 ( .A1(n759), .A2(n1011), .ZN(n764) );
  INV_X1 U846 ( .A(KEYINPUT33), .ZN(n762) );
  INV_X1 U847 ( .A(n781), .ZN(n776) );
  NAND2_X1 U848 ( .A1(n1011), .A2(n776), .ZN(n760) );
  NOR2_X1 U849 ( .A1(n762), .A2(n760), .ZN(n761) );
  XNOR2_X1 U850 ( .A(n761), .B(KEYINPUT101), .ZN(n767) );
  INV_X1 U851 ( .A(n767), .ZN(n763) );
  OR2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n766) );
  AND2_X1 U853 ( .A1(n764), .A2(n766), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n780), .A2(n765), .ZN(n773) );
  INV_X1 U855 ( .A(n766), .ZN(n770) );
  NAND2_X1 U856 ( .A1(G1976), .A2(G288), .ZN(n1012) );
  AND2_X1 U857 ( .A1(n1012), .A2(n767), .ZN(n768) );
  AND2_X1 U858 ( .A1(n776), .A2(n768), .ZN(n769) );
  NOR2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U860 ( .A(G1981), .B(G305), .ZN(n1000) );
  NOR2_X1 U861 ( .A1(n771), .A2(n1000), .ZN(n772) );
  AND2_X1 U862 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U863 ( .A(n774), .B(KEYINPUT102), .ZN(n786) );
  NOR2_X1 U864 ( .A1(G1981), .A2(G305), .ZN(n775) );
  XNOR2_X1 U865 ( .A(KEYINPUT24), .B(n775), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n784) );
  NOR2_X1 U867 ( .A1(G2090), .A2(G303), .ZN(n778) );
  NAND2_X1 U868 ( .A1(G8), .A2(n778), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n818) );
  XOR2_X1 U873 ( .A(G1986), .B(G290), .Z(n1008) );
  NAND2_X1 U874 ( .A1(n897), .A2(G105), .ZN(n787) );
  XNOR2_X1 U875 ( .A(n787), .B(KEYINPUT38), .ZN(n794) );
  NAND2_X1 U876 ( .A1(G117), .A2(n901), .ZN(n789) );
  NAND2_X1 U877 ( .A1(G141), .A2(n895), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U879 ( .A1(G129), .A2(n902), .ZN(n790) );
  XNOR2_X1 U880 ( .A(KEYINPUT89), .B(n790), .ZN(n791) );
  NOR2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n892) );
  NAND2_X1 U883 ( .A1(G1996), .A2(n892), .ZN(n803) );
  NAND2_X1 U884 ( .A1(G131), .A2(n895), .ZN(n796) );
  NAND2_X1 U885 ( .A1(G95), .A2(n897), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U887 ( .A(KEYINPUT88), .B(n797), .Z(n801) );
  NAND2_X1 U888 ( .A1(n901), .A2(G107), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G119), .A2(n902), .ZN(n798) );
  AND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n888) );
  NAND2_X1 U892 ( .A1(G1991), .A2(n888), .ZN(n802) );
  NAND2_X1 U893 ( .A1(n803), .A2(n802), .ZN(n822) );
  INV_X1 U894 ( .A(n822), .ZN(n924) );
  NAND2_X1 U895 ( .A1(n1008), .A2(n924), .ZN(n806) );
  NOR2_X1 U896 ( .A1(n805), .A2(n804), .ZN(n832) );
  NAND2_X1 U897 ( .A1(n806), .A2(n832), .ZN(n816) );
  XNOR2_X1 U898 ( .A(G2067), .B(KEYINPUT37), .ZN(n830) );
  NAND2_X1 U899 ( .A1(G140), .A2(n895), .ZN(n808) );
  NAND2_X1 U900 ( .A1(G104), .A2(n897), .ZN(n807) );
  NAND2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U902 ( .A(KEYINPUT34), .B(n809), .ZN(n814) );
  NAND2_X1 U903 ( .A1(G116), .A2(n901), .ZN(n811) );
  NAND2_X1 U904 ( .A1(G128), .A2(n902), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U906 ( .A(KEYINPUT35), .B(n812), .Z(n813) );
  NOR2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U908 ( .A(KEYINPUT36), .B(n815), .ZN(n882) );
  NOR2_X1 U909 ( .A1(n830), .A2(n882), .ZN(n937) );
  NAND2_X1 U910 ( .A1(n832), .A2(n937), .ZN(n828) );
  NAND2_X1 U911 ( .A1(n816), .A2(n828), .ZN(n817) );
  NOR2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U913 ( .A(n819), .B(KEYINPUT103), .ZN(n835) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n892), .ZN(n932) );
  NOR2_X1 U915 ( .A1(G1991), .A2(n888), .ZN(n926) );
  NOR2_X1 U916 ( .A1(G1986), .A2(G290), .ZN(n820) );
  XNOR2_X1 U917 ( .A(KEYINPUT104), .B(n820), .ZN(n821) );
  NOR2_X1 U918 ( .A1(n926), .A2(n821), .ZN(n823) );
  NOR2_X1 U919 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U920 ( .A1(n932), .A2(n824), .ZN(n825) );
  XOR2_X1 U921 ( .A(n825), .B(KEYINPUT105), .Z(n826) );
  XNOR2_X1 U922 ( .A(KEYINPUT39), .B(n826), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U924 ( .A(n829), .B(KEYINPUT106), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n830), .A2(n882), .ZN(n939) );
  NAND2_X1 U926 ( .A1(n831), .A2(n939), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U929 ( .A(n836), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U930 ( .A(G223), .ZN(n837) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n837), .ZN(G217) );
  NAND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n839) );
  INV_X1 U933 ( .A(G661), .ZN(n838) );
  NOR2_X1 U934 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U935 ( .A(n840), .B(KEYINPUT107), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U937 ( .A1(n842), .A2(n841), .ZN(G188) );
  INV_X1 U939 ( .A(G120), .ZN(G236) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  INV_X1 U941 ( .A(G69), .ZN(G235) );
  INV_X1 U942 ( .A(n843), .ZN(n845) );
  NOR2_X1 U943 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U944 ( .A(KEYINPUT108), .B(n846), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  XOR2_X1 U946 ( .A(G2100), .B(G2096), .Z(n848) );
  XNOR2_X1 U947 ( .A(KEYINPUT42), .B(G2678), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U949 ( .A(KEYINPUT43), .B(G2072), .Z(n850) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2090), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U952 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(G227) );
  XOR2_X1 U955 ( .A(G1976), .B(G1966), .Z(n856) );
  XNOR2_X1 U956 ( .A(G1981), .B(G1956), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U958 ( .A(G1971), .B(G1986), .Z(n858) );
  XNOR2_X1 U959 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U961 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U962 ( .A(G2474), .B(KEYINPUT41), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n864) );
  XOR2_X1 U964 ( .A(G1961), .B(KEYINPUT109), .Z(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(G229) );
  NAND2_X1 U966 ( .A1(G124), .A2(n902), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n865), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G112), .A2(n901), .ZN(n866) );
  XNOR2_X1 U969 ( .A(n866), .B(KEYINPUT110), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G136), .A2(n895), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G100), .A2(n897), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U974 ( .A1(n872), .A2(n871), .ZN(G162) );
  NAND2_X1 U975 ( .A1(G118), .A2(n901), .ZN(n881) );
  NAND2_X1 U976 ( .A1(n902), .A2(G130), .ZN(n873) );
  XNOR2_X1 U977 ( .A(KEYINPUT111), .B(n873), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G142), .A2(n895), .ZN(n875) );
  NAND2_X1 U979 ( .A1(G106), .A2(n897), .ZN(n874) );
  NAND2_X1 U980 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U981 ( .A(KEYINPUT112), .B(n876), .Z(n877) );
  XNOR2_X1 U982 ( .A(KEYINPUT45), .B(n877), .ZN(n878) );
  NOR2_X1 U983 ( .A1(n879), .A2(n878), .ZN(n880) );
  NAND2_X1 U984 ( .A1(n881), .A2(n880), .ZN(n886) );
  XNOR2_X1 U985 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n882), .B(KEYINPUT46), .ZN(n883) );
  XNOR2_X1 U987 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U988 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U989 ( .A(G162), .B(n887), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n888), .B(n925), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(n894) );
  XNOR2_X1 U993 ( .A(G160), .B(G164), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n908) );
  NAND2_X1 U995 ( .A1(n895), .A2(G139), .ZN(n896) );
  XOR2_X1 U996 ( .A(KEYINPUT113), .B(n896), .Z(n899) );
  NAND2_X1 U997 ( .A1(G103), .A2(n897), .ZN(n898) );
  NAND2_X1 U998 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U999 ( .A(KEYINPUT114), .B(n900), .ZN(n907) );
  NAND2_X1 U1000 ( .A1(G115), .A2(n901), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(G127), .A2(n902), .ZN(n903) );
  NAND2_X1 U1002 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1003 ( .A(KEYINPUT47), .B(n905), .Z(n906) );
  NOR2_X1 U1004 ( .A1(n907), .A2(n906), .ZN(n941) );
  XNOR2_X1 U1005 ( .A(n908), .B(n941), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n909), .ZN(G395) );
  XOR2_X1 U1007 ( .A(n1004), .B(n910), .Z(n912) );
  XNOR2_X1 U1008 ( .A(G286), .B(G171), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n915), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(KEYINPUT116), .B(n916), .ZN(G397) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(G401), .A2(n918), .ZN(n919) );
  AND2_X1 U1016 ( .A1(G319), .A2(n919), .ZN(n921) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1020 ( .A(G160), .B(G2084), .Z(n922) );
  XNOR2_X1 U1021 ( .A(KEYINPUT117), .B(n922), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n929) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1024 ( .A(KEYINPUT118), .B(n927), .Z(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n935) );
  XNOR2_X1 U1026 ( .A(G2090), .B(G162), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(n930), .B(KEYINPUT119), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1029 ( .A(KEYINPUT51), .B(n933), .Z(n934) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(n938), .B(KEYINPUT120), .ZN(n940) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n947) );
  XOR2_X1 U1034 ( .A(G164), .B(G2078), .Z(n944) );
  XNOR2_X1 U1035 ( .A(n942), .B(n941), .ZN(n943) );
  NOR2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1037 ( .A(KEYINPUT50), .B(n945), .Z(n946) );
  NOR2_X1 U1038 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1039 ( .A(KEYINPUT52), .B(n948), .ZN(n949) );
  INV_X1 U1040 ( .A(KEYINPUT55), .ZN(n970) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n970), .ZN(n950) );
  NAND2_X1 U1042 ( .A1(n950), .A2(G29), .ZN(n1029) );
  XOR2_X1 U1043 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n963) );
  XNOR2_X1 U1044 ( .A(G1996), .B(G32), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(G27), .B(n951), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n961) );
  XOR2_X1 U1047 ( .A(G1991), .B(G25), .Z(n954) );
  NAND2_X1 U1048 ( .A1(n954), .A2(G28), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(G2067), .B(G26), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(G33), .B(G2072), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(n957), .B(KEYINPUT121), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(n963), .B(n962), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(G35), .B(G2090), .ZN(n964) );
  NOR2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n968) );
  XOR2_X1 U1058 ( .A(G2084), .B(G34), .Z(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT54), .B(n966), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(n970), .B(n969), .ZN(n972) );
  INV_X1 U1062 ( .A(G29), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1064 ( .A1(G11), .A2(n973), .ZN(n1027) );
  XOR2_X1 U1065 ( .A(G1986), .B(G24), .Z(n976) );
  XOR2_X1 U1066 ( .A(G22), .B(KEYINPUT126), .Z(n974) );
  XNOR2_X1 U1067 ( .A(n974), .B(G1971), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(G23), .B(G1976), .ZN(n977) );
  NOR2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1071 ( .A(KEYINPUT58), .B(n979), .Z(n994) );
  XOR2_X1 U1072 ( .A(G1961), .B(G5), .Z(n989) );
  XNOR2_X1 U1073 ( .A(G1348), .B(KEYINPUT59), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(n980), .B(G4), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(G1981), .B(G6), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(G19), .B(G1341), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(G20), .B(G1956), .ZN(n985) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(KEYINPUT60), .B(n987), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(G21), .B(G1966), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(KEYINPUT125), .B(n992), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1087 ( .A(KEYINPUT61), .B(n995), .Z(n996) );
  NOR2_X1 U1088 ( .A1(G16), .A2(n996), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(KEYINPUT127), .B(n997), .ZN(n1025) );
  XNOR2_X1 U1090 ( .A(KEYINPUT56), .B(G16), .ZN(n1023) );
  XNOR2_X1 U1091 ( .A(n998), .B(G1348), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(G168), .B(G1966), .Z(n999) );
  NOR2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1094 ( .A(KEYINPUT57), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1021) );
  XOR2_X1 U1096 ( .A(n1004), .B(G1341), .Z(n1006) );
  XOR2_X1 U1097 ( .A(G171), .B(G1961), .Z(n1005) );
  NOR2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1019) );
  XNOR2_X1 U1100 ( .A(G303), .B(G1971), .ZN(n1010) );
  XNOR2_X1 U1101 ( .A(G299), .B(G1956), .ZN(n1009) );
  NOR2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1016) );
  INV_X1 U1103 ( .A(n1011), .ZN(n1013) );
  NAND2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1105 ( .A(n1014), .B(KEYINPUT123), .ZN(n1015) );
  NAND2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(KEYINPUT124), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

