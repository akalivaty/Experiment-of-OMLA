//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT88), .Z(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT99), .B(G952), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(G234), .A2(G237), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT21), .B(G898), .Z(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(G902), .A3(G953), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT89), .ZN(new_n197));
  XOR2_X1   g011(.A(G116), .B(G119), .Z(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT2), .B(G113), .ZN(new_n199));
  XOR2_X1   g013(.A(new_n198), .B(new_n199), .Z(new_n200));
  INV_X1    g014(.A(KEYINPUT78), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .A4(G104), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n205), .A2(G107), .B1(KEYINPUT78), .B2(KEYINPUT3), .ZN(new_n206));
  OAI22_X1  g020(.A1(new_n205), .A2(G107), .B1(KEYINPUT78), .B2(KEYINPUT3), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(G101), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT82), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT82), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n208), .A2(new_n212), .A3(G101), .A4(new_n209), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n204), .A2(new_n206), .A3(new_n207), .A4(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT79), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n208), .A2(G101), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n208), .A2(new_n217), .A3(G101), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT4), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT80), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n221), .A2(KEYINPUT4), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT80), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n218), .A2(new_n219), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  AOI211_X1 g041(.A(new_n200), .B(new_n214), .C1(new_n223), .C2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT5), .ZN(new_n229));
  INV_X1    g043(.A(G119), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(G116), .ZN(new_n231));
  OAI211_X1 g045(.A(G113), .B(new_n231), .C1(new_n198), .C2(new_n229), .ZN(new_n232));
  OR2_X1    g046(.A1(new_n198), .A2(new_n199), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n203), .A2(G104), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n205), .A2(G107), .ZN(new_n236));
  OAI21_X1  g050(.A(G101), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n216), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n197), .B1(new_n228), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G110), .B(G122), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n200), .ZN(new_n243));
  INV_X1    g057(.A(new_n214), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n220), .A2(KEYINPUT80), .A3(new_n222), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n225), .B1(new_n224), .B2(new_n226), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n243), .B(new_n244), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n239), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(KEYINPUT89), .A3(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n240), .A2(KEYINPUT6), .A3(new_n242), .A4(new_n249), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n247), .A2(KEYINPUT89), .A3(new_n248), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT89), .B1(new_n247), .B2(new_n248), .ZN(new_n252));
  NOR3_X1   g066(.A1(new_n251), .A2(new_n252), .A3(new_n241), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT6), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n214), .B1(new_n223), .B2(new_n227), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n239), .B1(new_n255), .B2(new_n243), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n254), .B1(new_n256), .B2(new_n241), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n250), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G143), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(G146), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT65), .B(G143), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(G146), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n263));
  INV_X1    g077(.A(G128), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(KEYINPUT1), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(KEYINPUT65), .A2(G143), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT65), .A2(G143), .ZN(new_n268));
  OAI21_X1  g082(.A(G146), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n260), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(new_n265), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT67), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  OR2_X1    g087(.A1(KEYINPUT65), .A2(G143), .ZN(new_n274));
  INV_X1    g088(.A(G146), .ZN(new_n275));
  NAND2_X1  g089(.A1(KEYINPUT65), .A2(G143), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n275), .A2(G143), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT1), .ZN(new_n281));
  OAI21_X1  g095(.A(G128), .B1(new_n260), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(G125), .B1(new_n273), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G125), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT64), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT0), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n264), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n280), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n287), .A2(new_n264), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n267), .A2(new_n268), .A3(G146), .ZN(new_n293));
  OAI211_X1 g107(.A(KEYINPUT64), .B(new_n288), .C1(new_n293), .C2(new_n278), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n291), .B1(new_n269), .B2(new_n270), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n285), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n284), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT90), .B(G224), .ZN(new_n299));
  INV_X1    g113(.A(G953), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n301), .B1(new_n284), .B2(new_n297), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n258), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G210), .B1(G237), .B2(G902), .ZN(new_n308));
  INV_X1    g122(.A(new_n284), .ZN(new_n309));
  INV_X1    g123(.A(new_n297), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT7), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  OAI211_X1 g126(.A(KEYINPUT7), .B(new_n301), .C1(new_n284), .C2(new_n297), .ZN(new_n313));
  INV_X1    g127(.A(new_n238), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n234), .A2(KEYINPUT91), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n241), .B(KEYINPUT8), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT91), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n233), .B(new_n232), .C1(new_n238), .C2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n303), .A2(new_n312), .A3(new_n313), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT92), .ZN(new_n321));
  INV_X1    g135(.A(new_n319), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(new_n298), .B2(new_n302), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT92), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n323), .A2(new_n324), .A3(new_n313), .A4(new_n312), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n256), .A2(new_n241), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n321), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G902), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n307), .A2(new_n308), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n308), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n240), .A2(new_n242), .A3(new_n249), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n326), .A2(KEYINPUT6), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n305), .B1(new_n335), .B2(new_n250), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n332), .B1(new_n336), .B2(new_n329), .ZN(new_n337));
  AOI211_X1 g151(.A(new_n188), .B(new_n196), .C1(new_n331), .C2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G237), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n300), .A3(G214), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n340), .A2(G143), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n274), .A3(new_n276), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(KEYINPUT18), .A2(G131), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n285), .A2(KEYINPUT74), .A3(G140), .ZN(new_n346));
  INV_X1    g160(.A(G140), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G125), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(new_n347), .B2(G125), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n346), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT93), .B1(new_n351), .B2(new_n275), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n348), .ZN(new_n353));
  INV_X1    g167(.A(new_n346), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT93), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n356), .A3(G146), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n285), .A2(G140), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n348), .A2(new_n358), .A3(new_n275), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n352), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n345), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT19), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n348), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n351), .B2(new_n362), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT95), .B1(new_n364), .B2(G146), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT16), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n348), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(new_n351), .B2(new_n366), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G146), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n355), .A2(KEYINPUT19), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT95), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n370), .A2(new_n371), .A3(new_n275), .A4(new_n363), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n365), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n341), .A2(new_n342), .A3(G131), .ZN(new_n374));
  AOI21_X1  g188(.A(G131), .B1(new_n341), .B2(new_n342), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT94), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G131), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n343), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT94), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n341), .A2(new_n342), .A3(G131), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n361), .B1(new_n373), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G113), .B(G122), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(new_n205), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT17), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n378), .A2(new_n388), .A3(new_n380), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n275), .B(new_n367), .C1(new_n351), .C2(new_n366), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n374), .A2(KEYINPUT17), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n389), .A2(new_n369), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n361), .A3(new_n385), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n387), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(KEYINPUT97), .A3(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(G475), .A2(G902), .ZN(new_n397));
  XOR2_X1   g211(.A(new_n397), .B(KEYINPUT96), .Z(new_n398));
  AOI21_X1  g212(.A(KEYINPUT20), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n398), .ZN(new_n400));
  AOI211_X1 g214(.A(new_n395), .B(new_n400), .C1(new_n387), .C2(new_n393), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n396), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G475), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n392), .A2(new_n361), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n386), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n393), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n403), .B1(new_n406), .B2(new_n328), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT97), .ZN(new_n408));
  AOI211_X1 g222(.A(new_n408), .B(KEYINPUT20), .C1(new_n387), .C2(new_n393), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n407), .B1(new_n409), .B2(new_n398), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n402), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT98), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n259), .A2(G128), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n261), .B2(G128), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT13), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT13), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n261), .A2(new_n416), .A3(G128), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n415), .A2(G134), .A3(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G116), .B(G122), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(new_n203), .ZN(new_n420));
  INV_X1    g234(.A(G134), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n414), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n419), .A2(new_n203), .ZN(new_n424));
  INV_X1    g238(.A(G116), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(KEYINPUT14), .A3(G122), .ZN(new_n426));
  INV_X1    g240(.A(new_n419), .ZN(new_n427));
  OAI211_X1 g241(.A(G107), .B(new_n426), .C1(new_n427), .C2(KEYINPUT14), .ZN(new_n428));
  INV_X1    g242(.A(new_n422), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n414), .A2(new_n421), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n424), .B(new_n428), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT9), .B(G234), .ZN(new_n432));
  INV_X1    g246(.A(G217), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n432), .A2(new_n433), .A3(G953), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n423), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n434), .B1(new_n423), .B2(new_n431), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n412), .B(new_n328), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G478), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(KEYINPUT15), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n437), .B(new_n439), .Z(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n411), .A2(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n338), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT30), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT11), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n421), .B2(G137), .ZN(new_n446));
  INV_X1    g260(.A(G137), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(KEYINPUT11), .A3(G134), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n421), .A2(G137), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n450), .A2(new_n377), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n447), .A2(G134), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n452), .A2(new_n449), .A3(G131), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(new_n273), .B2(new_n283), .ZN(new_n455));
  NAND2_X1  g269(.A1(KEYINPUT66), .A2(G131), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n450), .B(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n292), .B2(new_n296), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n444), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n263), .B1(new_n262), .B2(new_n265), .ZN(new_n460));
  AND4_X1   g274(.A1(new_n263), .A2(new_n269), .A3(new_n270), .A4(new_n265), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n283), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n454), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n457), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n275), .B1(new_n274), .B2(new_n276), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n290), .B1(new_n466), .B2(new_n260), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n277), .A2(new_n279), .B1(new_n287), .B2(new_n264), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n467), .B1(KEYINPUT64), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n290), .B1(new_n468), .B2(new_n286), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n464), .A2(new_n471), .A3(KEYINPUT30), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n459), .A2(new_n472), .A3(new_n243), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n455), .A2(new_n458), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n200), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n339), .A2(new_n300), .A3(G210), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n476), .B(new_n215), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n477), .B(new_n478), .Z(new_n479));
  NAND3_X1  g293(.A1(new_n473), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT31), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n473), .A2(KEYINPUT31), .A3(new_n475), .A4(new_n479), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n479), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT68), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n243), .B1(new_n474), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n464), .A2(new_n471), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT68), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT28), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT28), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n243), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n491), .B1(new_n475), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n485), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n484), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT69), .ZN(new_n496));
  NOR2_X1   g310(.A1(G472), .A2(G902), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT69), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n484), .A2(new_n498), .A3(new_n494), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT32), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n496), .A2(KEYINPUT32), .A3(new_n497), .A4(new_n499), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n493), .A2(new_n485), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT70), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n490), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n490), .A2(new_n505), .ZN(new_n507));
  OAI211_X1 g321(.A(KEYINPUT29), .B(new_n504), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n473), .A2(new_n475), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT29), .B1(new_n509), .B2(new_n485), .ZN(new_n510));
  INV_X1    g324(.A(new_n504), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n510), .B1(new_n511), .B2(new_n490), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(new_n512), .A3(new_n328), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G472), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n502), .A2(new_n503), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n433), .B1(G234), .B2(new_n328), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n264), .A2(KEYINPUT71), .A3(G119), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT71), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n230), .B2(G128), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n264), .A2(G119), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(KEYINPUT72), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT24), .B(G110), .Z(new_n523));
  OAI21_X1  g337(.A(KEYINPUT23), .B1(new_n264), .B2(G119), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT73), .B1(new_n230), .B2(G128), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n524), .B(new_n525), .Z(new_n526));
  OAI22_X1  g340(.A1(new_n522), .A2(new_n523), .B1(new_n526), .B2(G110), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(new_n369), .A3(new_n359), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n369), .A2(new_n390), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(G110), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n522), .A2(new_n523), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT75), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n528), .A2(KEYINPUT75), .A3(new_n532), .ZN(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT22), .B(G137), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n300), .A2(G221), .A3(G234), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n539), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n533), .A2(new_n534), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT25), .B1(new_n543), .B2(new_n328), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT25), .ZN(new_n545));
  AOI211_X1 g359(.A(new_n545), .B(G902), .C1(new_n540), .C2(new_n542), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n516), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n516), .A2(G902), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n515), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G221), .ZN(new_n552));
  INV_X1    g366(.A(new_n432), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n552), .B1(new_n553), .B2(new_n328), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT76), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n300), .A2(G227), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT77), .ZN(new_n558));
  XNOR2_X1  g372(.A(G110), .B(G140), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G128), .B1(new_n293), .B2(new_n281), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n260), .B2(new_n466), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n273), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n314), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n273), .B2(new_n283), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n565), .A2(new_n567), .B1(new_n569), .B2(new_n314), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n292), .A2(new_n296), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n571), .B(new_n244), .C1(new_n245), .C2(new_n246), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n457), .B(KEYINPUT84), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n570), .A2(new_n572), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT86), .B1(new_n575), .B2(new_n465), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT86), .ZN(new_n577));
  AOI211_X1 g391(.A(new_n577), .B(new_n457), .C1(new_n570), .C2(new_n572), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n561), .B(new_n574), .C1(new_n576), .C2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT87), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n462), .A2(new_n314), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n238), .B1(new_n273), .B2(new_n563), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n465), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT12), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g399(.A(KEYINPUT12), .B(new_n465), .C1(new_n581), .C2(new_n582), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(KEYINPUT85), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT85), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n583), .A2(new_n588), .A3(new_n584), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n574), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n560), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n579), .A2(new_n580), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n580), .B1(new_n579), .B2(new_n591), .ZN(new_n593));
  OAI21_X1  g407(.A(G469), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n560), .B(new_n574), .C1(new_n576), .C2(new_n578), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n590), .A2(new_n561), .ZN(new_n596));
  INV_X1    g410(.A(G469), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .A4(new_n328), .ZN(new_n598));
  NAND2_X1  g412(.A1(G469), .A2(G902), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n556), .B1(new_n594), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n443), .A2(new_n551), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  AND2_X1   g417(.A1(new_n496), .A2(new_n499), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n496), .A2(new_n328), .A3(new_n499), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n604), .A2(new_n497), .B1(new_n605), .B2(G472), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n606), .A2(new_n601), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(new_n550), .A3(new_n338), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  OAI22_X1  g423(.A1(new_n435), .A2(new_n436), .B1(KEYINPUT100), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n423), .A2(new_n431), .ZN(new_n611));
  INV_X1    g425(.A(new_n434), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n423), .A2(new_n431), .A3(new_n434), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT100), .B(KEYINPUT33), .Z(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n610), .A2(new_n616), .A3(G478), .A4(new_n328), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n328), .B1(new_n435), .B2(new_n436), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n438), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n411), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n622), .B(KEYINPUT101), .Z(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n608), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT34), .B(G104), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  NOR2_X1   g441(.A1(new_n399), .A2(new_n401), .ZN(new_n628));
  INV_X1    g442(.A(new_n407), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n441), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n608), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT102), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT35), .B(G107), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NOR2_X1   g448(.A1(new_n539), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n533), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n548), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n547), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n443), .A2(new_n607), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT37), .B(G110), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G12));
  AND3_X1   g457(.A1(new_n515), .A2(new_n601), .A3(new_n640), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n188), .B1(new_n331), .B2(new_n337), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n192), .B1(G900), .B2(new_n194), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n630), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n645), .A2(KEYINPUT104), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(KEYINPUT104), .B1(new_n645), .B2(new_n648), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n644), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  AOI21_X1  g467(.A(new_n440), .B1(new_n402), .B2(new_n410), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT106), .B(KEYINPUT39), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n646), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n601), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT40), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n331), .A2(new_n337), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT38), .ZN(new_n663));
  INV_X1    g477(.A(new_n640), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n475), .A2(new_n492), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n485), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n667), .A2(KEYINPUT105), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n480), .B1(new_n667), .B2(KEYINPUT105), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n328), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(G472), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n502), .A2(new_n503), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n188), .B1(new_n658), .B2(KEYINPUT40), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n661), .A2(new_n665), .A3(new_n672), .A4(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n674), .B(new_n261), .Z(G45));
  AOI211_X1 g489(.A(new_n647), .B(new_n620), .C1(new_n402), .C2(new_n410), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n644), .A2(new_n645), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  NAND3_X1  g492(.A1(new_n595), .A2(new_n328), .A3(new_n596), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G469), .ZN(new_n680));
  INV_X1    g494(.A(new_n554), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n680), .A2(new_n598), .A3(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n551), .A2(new_n623), .A3(new_n338), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT41), .B(G113), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G15));
  INV_X1    g499(.A(new_n630), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n551), .A2(new_n338), .A3(new_n686), .A4(new_n682), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G116), .ZN(G18));
  AND2_X1   g502(.A1(new_n515), .A2(new_n195), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n640), .A2(new_n442), .ZN(new_n690));
  AOI21_X1  g504(.A(KEYINPUT107), .B1(new_n645), .B2(new_n682), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n645), .A2(new_n682), .A3(KEYINPUT107), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n689), .B(new_n690), .C1(new_n691), .C2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G119), .ZN(G21));
  INV_X1    g509(.A(new_n188), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n308), .B1(new_n307), .B2(new_n330), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n336), .A2(new_n332), .A3(new_n329), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n696), .B(new_n654), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT108), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n645), .A2(new_n701), .A3(new_n654), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n506), .A2(new_n507), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n485), .B1(new_n704), .B2(new_n493), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n484), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n497), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n605), .A2(G472), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n707), .A2(new_n708), .A3(new_n550), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n682), .A2(new_n195), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n703), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  NAND3_X1  g527(.A1(new_n707), .A2(new_n708), .A3(new_n676), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n715), .B(new_n640), .C1(new_n693), .C2(new_n691), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G125), .ZN(G27));
  AND4_X1   g531(.A1(new_n696), .A2(new_n676), .A3(new_n331), .A4(new_n337), .ZN(new_n718));
  INV_X1    g532(.A(new_n576), .ZN(new_n719));
  INV_X1    g533(.A(new_n578), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n721), .A2(KEYINPUT109), .A3(new_n561), .A4(new_n574), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n579), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n722), .A2(G469), .A3(new_n591), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n554), .B1(new_n600), .B2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n515), .A2(new_n718), .A3(new_n550), .A4(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n728), .A3(KEYINPUT111), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT111), .B1(new_n727), .B2(new_n728), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT42), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n727), .A2(new_n728), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n727), .A2(KEYINPUT42), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n729), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  NAND3_X1  g553(.A1(new_n551), .A2(new_n648), .A3(new_n726), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n331), .A2(new_n337), .A3(new_n696), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n421), .ZN(G36));
  NAND3_X1  g557(.A1(new_n621), .A2(new_n402), .A3(new_n410), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT43), .ZN(new_n745));
  OR3_X1    g559(.A1(new_n606), .A2(new_n745), .A3(new_n664), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(KEYINPUT112), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n606), .A2(new_n745), .A3(new_n664), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n749), .B1(new_n750), .B2(KEYINPUT44), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n741), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n579), .A2(new_n591), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT87), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n579), .A2(new_n580), .A3(new_n591), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n722), .A2(KEYINPUT45), .A3(new_n591), .A4(new_n724), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(G469), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(KEYINPUT46), .A3(new_n599), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n598), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT46), .B1(new_n759), .B2(new_n599), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n681), .B(new_n657), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n746), .A2(new_n747), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n752), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  OAI21_X1  g581(.A(new_n681), .B1(new_n761), .B2(new_n762), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT113), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n515), .A2(new_n550), .ZN(new_n772));
  XOR2_X1   g586(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n773));
  OAI211_X1 g587(.A(new_n681), .B(new_n773), .C1(new_n761), .C2(new_n762), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n771), .A2(new_n718), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  INV_X1    g590(.A(new_n192), .ZN(new_n777));
  INV_X1    g591(.A(new_n745), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n709), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n645), .A2(new_n682), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT107), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n779), .B1(new_n782), .B2(new_n692), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n771), .A2(new_n774), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n680), .A2(new_n598), .A3(new_n556), .ZN(new_n786));
  AOI211_X1 g600(.A(new_n741), .B(new_n779), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n779), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n663), .A2(new_n696), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n789), .A3(new_n682), .ZN(new_n790));
  NOR2_X1   g604(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n790), .A2(new_n794), .A3(new_n792), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n680), .A2(new_n598), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n741), .A2(new_n796), .A3(new_n554), .A4(new_n192), .ZN(new_n797));
  AND4_X1   g611(.A1(new_n502), .A2(new_n503), .A3(new_n550), .A4(new_n671), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n411), .A2(new_n621), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n797), .A2(new_n778), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(new_n708), .A3(new_n640), .A4(new_n707), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n793), .A2(new_n795), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n784), .B1(new_n787), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n190), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n801), .A2(new_n551), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT48), .Z(new_n807));
  NOR3_X1   g621(.A1(new_n787), .A2(new_n803), .A3(new_n784), .ZN(new_n808));
  OR4_X1    g622(.A1(new_n783), .A2(new_n805), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n715), .A2(new_n726), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n440), .A2(new_n628), .A3(new_n629), .A4(new_n646), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n515), .A2(new_n601), .A3(new_n811), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n664), .B(new_n741), .C1(new_n810), .C2(new_n812), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n742), .B(new_n813), .C1(new_n732), .C2(new_n737), .ZN(new_n814));
  INV_X1    g628(.A(new_n338), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n441), .A2(new_n410), .A3(new_n402), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT115), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n818));
  INV_X1    g632(.A(new_n816), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n338), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n817), .A2(new_n607), .A3(new_n820), .A4(new_n550), .ZN(new_n821));
  INV_X1    g635(.A(new_n622), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n607), .A2(new_n550), .A3(new_n338), .A4(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n821), .A2(new_n602), .A3(new_n641), .A4(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n694), .A2(new_n683), .A3(new_n687), .A4(new_n712), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n515), .A2(new_n338), .A3(new_n550), .A4(new_n682), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n710), .B1(new_n700), .B2(new_n702), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n686), .A2(new_n828), .B1(new_n829), .B2(new_n709), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(KEYINPUT114), .A3(new_n683), .A4(new_n694), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n824), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n664), .B(new_n714), .C1(new_n782), .C2(new_n692), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n515), .A2(new_n601), .A3(new_n640), .ZN(new_n834));
  INV_X1    g648(.A(new_n649), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n834), .A2(new_n835), .A3(new_n650), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT117), .B1(new_n640), .B2(new_n647), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n547), .A2(new_n639), .A3(new_n839), .A4(new_n646), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n703), .A2(new_n672), .A3(new_n726), .A4(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n837), .A2(KEYINPUT52), .A3(new_n677), .A4(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n652), .A3(new_n677), .A4(new_n716), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n814), .A2(new_n832), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT53), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n833), .B2(new_n836), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n652), .A2(new_n716), .A3(KEYINPUT116), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n677), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n842), .A2(KEYINPUT52), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n846), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n814), .A3(new_n832), .A4(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n849), .A2(KEYINPUT54), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n848), .A2(new_n856), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n742), .B1(new_n732), .B2(new_n737), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n824), .A2(new_n825), .A3(new_n813), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n855), .A2(KEYINPUT53), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n859), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n797), .A2(new_n623), .A3(new_n798), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n858), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI22_X1  g680(.A1(new_n809), .A2(new_n866), .B1(G952), .B2(G953), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n796), .A2(KEYINPUT49), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n796), .A2(KEYINPUT49), .ZN(new_n869));
  NOR4_X1   g683(.A1(new_n663), .A2(new_n744), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n555), .A3(new_n696), .A4(new_n798), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n867), .A2(new_n871), .ZN(G75));
  INV_X1    g686(.A(G210), .ZN(new_n873));
  AOI211_X1 g687(.A(new_n873), .B(new_n328), .C1(new_n859), .C2(new_n863), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n258), .B(KEYINPUT119), .Z(new_n875));
  XNOR2_X1  g689(.A(new_n305), .B(KEYINPUT55), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n875), .B(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT56), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n878), .B1(KEYINPUT120), .B2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n874), .A2(KEYINPUT56), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n880), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n859), .A2(new_n863), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n883), .A2(G210), .A3(G902), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n882), .B1(new_n884), .B2(new_n879), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n300), .A2(G952), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n881), .A2(new_n885), .A3(new_n886), .ZN(G51));
  NAND2_X1  g701(.A1(new_n599), .A2(KEYINPUT57), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n599), .A2(KEYINPUT57), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n859), .A2(new_n860), .A3(new_n863), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n860), .B1(new_n859), .B2(new_n863), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n888), .B(new_n889), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n595), .A2(new_n596), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n759), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n883), .A2(G902), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n886), .B1(new_n894), .B2(new_n896), .ZN(G54));
  INV_X1    g711(.A(new_n886), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n883), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n899));
  INV_X1    g713(.A(new_n394), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n899), .A2(KEYINPUT121), .A3(new_n900), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(G60));
  NAND2_X1  g720(.A1(G478), .A2(G902), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT59), .Z(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n858), .B2(new_n864), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n610), .A2(new_n616), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT122), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n898), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n908), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n913), .B(new_n911), .C1(new_n890), .C2(new_n891), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n912), .A2(new_n915), .ZN(G63));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT60), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n883), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n543), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n886), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n918), .B1(new_n859), .B2(new_n863), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n636), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n922), .B(new_n924), .C1(KEYINPUT123), .C2(KEYINPUT61), .ZN(new_n925));
  OAI211_X1 g739(.A(KEYINPUT123), .B(new_n898), .C1(new_n923), .C2(new_n543), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n898), .B1(new_n923), .B2(new_n543), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n883), .A2(new_n636), .A3(new_n919), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n926), .B(new_n927), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n930), .ZN(G66));
  AOI21_X1  g745(.A(new_n300), .B1(new_n193), .B2(new_n299), .ZN(new_n932));
  INV_X1    g746(.A(new_n832), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(new_n300), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n875), .B1(G898), .B2(new_n300), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n934), .B(new_n935), .Z(G69));
  NAND2_X1  g750(.A1(new_n459), .A2(new_n472), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(new_n364), .Z(new_n938));
  NOR2_X1   g752(.A1(new_n658), .A2(new_n741), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n622), .A2(new_n816), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n939), .A2(new_n551), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT124), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n766), .A2(new_n775), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n652), .A2(new_n716), .A3(KEYINPUT116), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT116), .B1(new_n652), .B2(new_n716), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n948), .A2(KEYINPUT62), .A3(new_n674), .A4(new_n677), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n851), .A2(new_n674), .A3(new_n677), .A4(new_n852), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n945), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n938), .B1(new_n953), .B2(G953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT125), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT125), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n956), .B(new_n938), .C1(new_n953), .C2(G953), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n300), .B1(G227), .B2(G900), .ZN(new_n958));
  INV_X1    g772(.A(new_n763), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n551), .A3(new_n703), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n861), .A2(new_n960), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n948), .A2(new_n677), .A3(new_n775), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n961), .A2(new_n962), .A3(new_n300), .A4(new_n766), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n938), .B1(G900), .B2(G953), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n958), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n955), .A2(new_n957), .A3(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n955), .A2(KEYINPUT126), .A3(new_n957), .A4(new_n965), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n963), .A2(KEYINPUT127), .A3(new_n964), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n955), .A2(new_n957), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT127), .B1(new_n963), .B2(new_n964), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n958), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n970), .A2(new_n974), .ZN(G72));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  NAND3_X1  g791(.A1(new_n961), .A2(new_n962), .A3(new_n766), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n978), .B2(new_n933), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n509), .A2(new_n479), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n485), .B1(new_n473), .B2(new_n475), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n953), .A2(new_n832), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n984), .B2(new_n977), .ZN(new_n985));
  INV_X1    g799(.A(new_n980), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n986), .A2(new_n977), .A3(new_n983), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n849), .A2(new_n857), .A3(new_n987), .ZN(new_n988));
  NOR4_X1   g802(.A1(new_n981), .A2(new_n985), .A3(new_n988), .A4(new_n886), .ZN(G57));
endmodule


