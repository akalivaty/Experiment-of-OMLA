//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT22), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(G137), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G125), .B(G140), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT77), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G125), .ZN(new_n196));
  AOI22_X1  g010(.A1(new_n192), .A2(KEYINPUT16), .B1(new_n193), .B2(new_n196), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n194), .A2(new_n195), .A3(KEYINPUT77), .A4(G125), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n195), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT16), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n196), .A2(new_n193), .ZN(new_n206));
  AND4_X1   g020(.A1(G146), .A2(new_n205), .A3(new_n206), .A4(new_n198), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n201), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n211));
  INV_X1    g025(.A(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G128), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT23), .B1(new_n210), .B2(G119), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G110), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT76), .B1(new_n212), .B2(G128), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT76), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n210), .A3(G119), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n221), .A3(new_n213), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT24), .B(G110), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n209), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n222), .A2(new_n223), .ZN(new_n228));
  OR2_X1    g042(.A1(new_n228), .A2(KEYINPUT78), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n228), .A2(KEYINPUT78), .B1(new_n216), .B2(new_n217), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n192), .A2(new_n200), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n208), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n191), .B1(new_n227), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G902), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n226), .B(new_n190), .C1(new_n231), .C2(new_n233), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT74), .B(G217), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(G234), .B2(new_n236), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(KEYINPUT75), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n235), .A2(new_n237), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n242), .A2(G902), .ZN(new_n247));
  XOR2_X1   g061(.A(new_n247), .B(KEYINPUT80), .Z(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT73), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(G101), .ZN(new_n252));
  NOR2_X1   g066(.A1(G237), .A2(G953), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G210), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n252), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n200), .A2(G143), .ZN(new_n260));
  INV_X1    g074(.A(G143), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G146), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n261), .A2(G146), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT65), .B1(new_n200), .B2(G143), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n261), .A3(G146), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n264), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n210), .B1(new_n260), .B2(KEYINPUT1), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n263), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT69), .ZN(new_n271));
  INV_X1    g085(.A(G137), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n272), .A2(KEYINPUT11), .A3(G134), .ZN(new_n273));
  AND2_X1   g087(.A1(KEYINPUT66), .A2(G134), .ZN(new_n274));
  NOR2_X1   g088(.A1(KEYINPUT66), .A2(G134), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n273), .B1(new_n276), .B2(G137), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n272), .B1(new_n274), .B2(new_n275), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT11), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G131), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n277), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n278), .B1(G134), .B2(new_n272), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G131), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n285), .B(new_n263), .C1(new_n268), .C2(new_n269), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n271), .A2(new_n282), .A3(new_n284), .A4(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(G143), .B(G146), .ZN(new_n288));
  AND2_X1   g102(.A1(KEYINPUT0), .A2(G128), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT0), .B(G128), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n290), .B1(new_n268), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n277), .A2(new_n281), .A3(new_n280), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n281), .B1(new_n277), .B2(new_n280), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(KEYINPUT2), .A2(G113), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT67), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT67), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(KEYINPUT2), .A3(G113), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT2), .ZN(new_n302));
  INV_X1    g116(.A(G113), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G116), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n212), .ZN(new_n306));
  NAND2_X1  g120(.A1(G116), .A2(G119), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n301), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT68), .ZN(new_n310));
  AND2_X1   g124(.A1(G116), .A2(G119), .ZN(new_n311));
  NOR2_X1   g125(.A1(G116), .A2(G119), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n306), .A2(KEYINPUT68), .A3(new_n307), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n298), .A2(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n309), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OR2_X1    g131(.A1(new_n317), .A2(KEYINPUT70), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(KEYINPUT70), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n287), .A2(new_n296), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT28), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n282), .A2(new_n284), .A3(new_n270), .ZN(new_n324));
  OR2_X1    g138(.A1(KEYINPUT66), .A2(G134), .ZN(new_n325));
  NAND2_X1  g139(.A1(KEYINPUT66), .A2(G134), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT11), .B1(new_n327), .B2(new_n272), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(G137), .A3(new_n326), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n272), .A2(KEYINPUT11), .A3(G134), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(G131), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n292), .B1(new_n332), .B2(new_n282), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n317), .B1(new_n324), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n321), .B1(new_n320), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n258), .B1(new_n323), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(new_n324), .B2(new_n333), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n287), .A2(new_n296), .A3(KEYINPUT30), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n338), .A2(new_n339), .A3(new_n317), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n320), .A2(new_n257), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT31), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n338), .A2(new_n339), .A3(new_n317), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT31), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n343), .A2(new_n344), .A3(new_n320), .A4(new_n257), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n336), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(G472), .A2(G902), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT32), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n346), .A2(KEYINPUT32), .A3(new_n347), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G472), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n354));
  INV_X1    g168(.A(new_n335), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT72), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n355), .A2(new_n356), .A3(new_n322), .A4(new_n257), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n343), .A2(new_n320), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT72), .B1(new_n358), .B2(new_n258), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n323), .A2(new_n335), .A3(new_n258), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n354), .B(new_n357), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n287), .A2(new_n296), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n318), .A2(new_n319), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n320), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n323), .B1(new_n365), .B2(KEYINPUT28), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n258), .A2(new_n354), .ZN(new_n367));
  AOI21_X1  g181(.A(G902), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n353), .B1(new_n361), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n251), .B1(new_n352), .B2(new_n369), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n346), .A2(KEYINPUT32), .A3(new_n347), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT32), .B1(new_n346), .B2(new_n347), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n361), .A2(new_n368), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G472), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n375), .A3(KEYINPUT73), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n250), .B1(new_n370), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT96), .B1(new_n210), .B2(G143), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT96), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n261), .A3(G128), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n380), .A3(KEYINPUT13), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n210), .A2(G143), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT13), .B1(new_n378), .B2(new_n380), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n381), .B(new_n382), .C1(new_n383), .C2(KEYINPUT97), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n383), .A2(KEYINPUT97), .ZN(new_n385));
  OAI21_X1  g199(.A(G134), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n378), .A2(new_n380), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n387), .A2(new_n276), .A3(new_n382), .ZN(new_n388));
  INV_X1    g202(.A(G122), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G116), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n305), .A2(G122), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT95), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT95), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(G107), .ZN(new_n395));
  INV_X1    g209(.A(G107), .ZN(new_n396));
  INV_X1    g210(.A(new_n394), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n396), .B1(new_n397), .B2(new_n392), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n388), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n386), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n305), .A2(KEYINPUT14), .A3(G122), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n390), .A2(new_n391), .ZN(new_n402));
  OAI211_X1 g216(.A(G107), .B(new_n401), .C1(new_n402), .C2(KEYINPUT14), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n276), .B1(new_n387), .B2(new_n382), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n398), .B(new_n403), .C1(new_n388), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT9), .B(G234), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n241), .A2(new_n407), .A3(G953), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n400), .A2(new_n405), .A3(new_n408), .ZN(new_n411));
  AOI21_X1  g225(.A(G902), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G478), .ZN(new_n413));
  OAI22_X1  g227(.A1(new_n412), .A2(KEYINPUT98), .B1(KEYINPUT15), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n411), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n408), .B1(new_n400), .B2(new_n405), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n236), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT98), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n413), .A2(KEYINPUT15), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n412), .A2(KEYINPUT98), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n414), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT99), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n414), .A2(new_n420), .A3(KEYINPUT99), .A4(new_n421), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(G146), .B1(new_n197), .B2(new_n198), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(new_n207), .ZN(new_n428));
  INV_X1    g242(.A(G237), .ZN(new_n429));
  AND4_X1   g243(.A1(G143), .A2(new_n429), .A3(new_n187), .A4(G214), .ZN(new_n430));
  AOI21_X1  g244(.A(G143), .B1(new_n253), .B2(G214), .ZN(new_n431));
  OAI21_X1  g245(.A(G131), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT17), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n429), .A2(new_n187), .A3(G214), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n261), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n253), .A2(G143), .A3(G214), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n281), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n432), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT92), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n432), .A2(new_n437), .A3(KEYINPUT92), .A4(new_n433), .ZN(new_n441));
  OR2_X1    g255(.A1(new_n432), .A2(new_n433), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n428), .A2(new_n440), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G113), .B(G122), .ZN(new_n444));
  INV_X1    g258(.A(G104), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n444), .B(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(KEYINPUT18), .B(G131), .C1(new_n430), .C2(new_n431), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n202), .A2(new_n204), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G146), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n232), .ZN(new_n450));
  NAND2_X1  g264(.A1(KEYINPUT18), .A2(G131), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n435), .A2(new_n436), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n447), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT91), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT91), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n447), .A2(new_n450), .A3(new_n452), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n443), .A2(new_n446), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT93), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n443), .A2(KEYINPUT93), .A3(new_n457), .A4(new_n446), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n443), .A2(new_n457), .ZN(new_n463));
  INV_X1    g277(.A(new_n446), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT94), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT94), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n463), .A2(new_n467), .A3(new_n464), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n462), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n236), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G475), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n432), .A2(new_n437), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n448), .B(KEYINPUT19), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n208), .B(new_n472), .C1(new_n473), .C2(G146), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n446), .B1(new_n457), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n462), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT20), .ZN(new_n478));
  NOR2_X1   g292(.A1(G475), .A2(G902), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n475), .B1(new_n460), .B2(new_n461), .ZN(new_n481));
  INV_X1    g295(.A(new_n479), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT20), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n471), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n187), .A2(G952), .ZN(new_n486));
  INV_X1    g300(.A(G234), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n486), .B1(new_n487), .B2(new_n429), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI211_X1 g303(.A(new_n236), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT21), .B(G898), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n426), .A2(new_n485), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G221), .B1(new_n407), .B2(G902), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  XOR2_X1   g309(.A(KEYINPUT86), .B(G469), .Z(new_n496));
  OAI21_X1  g310(.A(KEYINPUT3), .B1(new_n445), .B2(G107), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT3), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n396), .A3(G104), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n445), .A2(G107), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G101), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT81), .ZN(new_n503));
  INV_X1    g317(.A(G101), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n497), .A2(new_n499), .A3(new_n504), .A4(new_n500), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT81), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n501), .A2(new_n507), .A3(G101), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n503), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT4), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n501), .A2(new_n510), .A3(G101), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(new_n292), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n263), .B1(new_n269), .B2(new_n288), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT82), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n396), .A2(G104), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n500), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n514), .B1(new_n516), .B2(G101), .ZN(new_n517));
  AOI211_X1 g331(.A(KEYINPUT82), .B(new_n504), .C1(new_n515), .C2(new_n500), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n513), .B(new_n505), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT10), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n509), .A2(new_n512), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n294), .A2(new_n295), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT83), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n523), .B(new_n505), .C1(new_n517), .C2(new_n518), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(G104), .B(G107), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT82), .B1(new_n526), .B2(new_n504), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n516), .A2(new_n514), .A3(G101), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n523), .B1(new_n529), .B2(new_n505), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n271), .A2(KEYINPUT10), .A3(new_n286), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n521), .B(new_n522), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(G110), .B(G140), .ZN(new_n534));
  INV_X1    g348(.A(G227), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(G953), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n534), .B(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n533), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n505), .B1(new_n517), .B2(new_n518), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT83), .ZN(new_n541));
  INV_X1    g355(.A(new_n270), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n524), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n519), .ZN(new_n544));
  INV_X1    g358(.A(new_n522), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT12), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT84), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n547), .B1(new_n522), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n544), .A2(new_n545), .A3(new_n549), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n539), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n531), .A2(new_n532), .ZN(new_n554));
  INV_X1    g368(.A(new_n521), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n545), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n538), .B1(new_n556), .B2(new_n533), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n236), .B(new_n496), .C1(new_n553), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT87), .ZN(new_n559));
  AOI221_X4 g373(.A(new_n522), .B1(new_n548), .B2(new_n547), .C1(new_n543), .C2(new_n519), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n549), .B1(new_n544), .B2(new_n545), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n533), .B(new_n538), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n533), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n541), .A2(new_n524), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n271), .A2(new_n286), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT10), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n522), .B1(new_n566), .B2(new_n521), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n537), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(G902), .B1(new_n562), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT87), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n570), .A3(new_n496), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n559), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n533), .A2(KEYINPUT85), .A3(new_n538), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n573), .A2(new_n556), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT85), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n539), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n533), .B1(new_n560), .B2(new_n561), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n574), .A2(new_n576), .B1(new_n577), .B2(new_n537), .ZN(new_n578));
  OAI21_X1  g392(.A(G469), .B1(new_n578), .B2(G902), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n495), .B1(new_n572), .B2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(G110), .B(G122), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT5), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n313), .B2(new_n314), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n212), .A3(G116), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G113), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n309), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n587), .B1(new_n541), .B2(new_n524), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n501), .A2(new_n507), .A3(G101), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n507), .B1(new_n501), .B2(G101), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n501), .A2(new_n510), .A3(G101), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n317), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n582), .B1(new_n588), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n587), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n525), .B2(new_n530), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n317), .A2(new_n593), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n509), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n600), .A3(new_n581), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n596), .A2(new_n601), .A3(KEYINPUT6), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n292), .A2(G125), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n203), .B(new_n263), .C1(new_n268), .C2(new_n269), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(G224), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(G953), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n605), .B(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT6), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n609), .B(new_n582), .C1(new_n588), .C2(new_n595), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n602), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT7), .B1(new_n606), .B2(G953), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n603), .A2(new_n604), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n612), .B1(new_n603), .B2(new_n604), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n564), .A2(new_n597), .B1(new_n509), .B2(new_n599), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n616), .B2(new_n581), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n581), .B(KEYINPUT8), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n583), .B1(new_n306), .B2(new_n307), .ZN(new_n619));
  OAI211_X1 g433(.A(G113), .B(new_n585), .C1(new_n619), .C2(KEYINPUT88), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n308), .A2(KEYINPUT88), .A3(KEYINPUT5), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n309), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n541), .B2(new_n524), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n587), .A2(new_n540), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n618), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT89), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n619), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT88), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n586), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n632), .A2(new_n621), .B1(new_n316), .B2(new_n308), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n633), .B1(new_n525), .B2(new_n530), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n625), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(KEYINPUT89), .A3(new_n618), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n617), .A2(new_n629), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n611), .A2(new_n637), .A3(new_n236), .ZN(new_n638));
  OAI21_X1  g452(.A(G210), .B1(G237), .B2(G902), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n611), .A2(new_n637), .A3(new_n236), .A4(new_n639), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(KEYINPUT90), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT90), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n638), .A2(new_n644), .A3(new_n640), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(G214), .B1(G237), .B2(G902), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n377), .A2(new_n493), .A3(new_n580), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G101), .ZN(G3));
  NAND2_X1  g465(.A1(new_n346), .A2(new_n236), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n653), .A3(G472), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n346), .B(new_n236), .C1(KEYINPUT100), .C2(new_n353), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n250), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n580), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT33), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n411), .B2(KEYINPUT101), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n660), .B1(new_n415), .B2(new_n416), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n410), .B(new_n411), .C1(KEYINPUT101), .C2(new_n659), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(G478), .A3(new_n236), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n664), .B1(G478), .B2(new_n412), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n485), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n648), .B1(new_n641), .B2(new_n642), .ZN(new_n667));
  INV_X1    g481(.A(new_n492), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n658), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT34), .B(G104), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G6));
  NAND3_X1  g486(.A1(new_n480), .A2(KEYINPUT102), .A3(new_n483), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT102), .B1(new_n480), .B2(new_n483), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n467), .B1(new_n463), .B2(new_n464), .ZN(new_n677));
  AOI211_X1 g491(.A(KEYINPUT94), .B(new_n446), .C1(new_n443), .C2(new_n457), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(G902), .B1(new_n679), .B2(new_n462), .ZN(new_n680));
  INV_X1    g494(.A(G475), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT103), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n470), .A2(new_n683), .A3(G475), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n424), .A2(new_n682), .A3(new_n684), .A4(new_n425), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n676), .A2(new_n669), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n580), .A3(new_n657), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT35), .B(G107), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G9));
  NOR2_X1   g503(.A1(new_n227), .A2(new_n234), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n240), .A2(new_n243), .B1(new_n248), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n656), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n493), .A2(new_n580), .A3(new_n694), .A4(new_n649), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT37), .B(G110), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G12));
  NOR2_X1   g511(.A1(new_n558), .A2(KEYINPUT87), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n570), .B1(new_n569), .B2(new_n496), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n579), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n692), .A2(new_n248), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n244), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n700), .A2(new_n494), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(new_n370), .B2(new_n376), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n682), .A2(new_n684), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n478), .B1(new_n477), .B2(new_n479), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n481), .A2(KEYINPUT20), .A3(new_n482), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n673), .ZN(new_n710));
  INV_X1    g524(.A(new_n490), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n488), .B1(new_n711), .B2(G900), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n426), .A2(new_n705), .A3(new_n710), .A4(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n685), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(KEYINPUT104), .A3(new_n710), .A4(new_n712), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n704), .A2(new_n667), .A3(new_n715), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G128), .ZN(G30));
  XNOR2_X1  g533(.A(new_n712), .B(KEYINPUT39), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n580), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT40), .ZN(new_n722));
  INV_X1    g536(.A(new_n485), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n424), .A2(new_n425), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n358), .A2(new_n257), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n236), .B1(new_n365), .B2(new_n257), .ZN(new_n728));
  OAI21_X1  g542(.A(G472), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n373), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n725), .A2(new_n730), .A3(new_n647), .A4(new_n693), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n646), .B(KEYINPUT38), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n722), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G143), .ZN(G45));
  NAND2_X1  g549(.A1(new_n370), .A2(new_n376), .ZN(new_n736));
  AOI211_X1 g550(.A(new_n495), .B(new_n693), .C1(new_n572), .C2(new_n579), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n485), .A2(new_n665), .A3(new_n712), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n736), .A2(new_n737), .A3(new_n667), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G146), .ZN(G48));
  INV_X1    g554(.A(G469), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n569), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n572), .A2(new_n494), .A3(new_n743), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n744), .A2(new_n666), .A3(new_n669), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n377), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT41), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G113), .ZN(G15));
  INV_X1    g562(.A(new_n744), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n377), .A2(new_n686), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G116), .ZN(G18));
  NAND4_X1  g565(.A1(new_n723), .A2(new_n724), .A3(new_n702), .A4(new_n668), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n752), .B1(new_n370), .B2(new_n376), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n572), .A2(new_n494), .A3(new_n667), .A4(new_n743), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n742), .B1(new_n559), .B2(new_n571), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n757), .A2(KEYINPUT105), .A3(new_n494), .A4(new_n667), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n753), .A2(new_n759), .A3(KEYINPUT106), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT106), .B1(new_n753), .B2(new_n759), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n212), .ZN(G21));
  NAND3_X1  g577(.A1(new_n426), .A2(new_n485), .A3(new_n667), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n764), .A2(new_n744), .A3(new_n492), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n366), .A2(new_n257), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n342), .A2(new_n345), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n347), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n353), .B1(new_n346), .B2(new_n236), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AOI211_X1 g585(.A(KEYINPUT107), .B(new_n353), .C1(new_n346), .C2(new_n236), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n771), .A2(new_n250), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n765), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G122), .ZN(G24));
  NAND3_X1  g589(.A1(new_n485), .A2(new_n665), .A3(new_n712), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n776), .A2(new_n771), .A3(new_n693), .A4(new_n772), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT108), .B1(new_n759), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n759), .A2(KEYINPUT108), .A3(new_n777), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G125), .ZN(G27));
  XOR2_X1   g596(.A(KEYINPUT110), .B(KEYINPUT42), .Z(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n572), .A2(new_n785), .A3(new_n579), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n785), .B1(new_n572), .B2(new_n579), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n495), .A2(new_n648), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n643), .B2(new_n645), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n377), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n784), .B1(new_n792), .B2(new_n776), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n700), .A2(KEYINPUT109), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n572), .A2(new_n785), .A3(new_n579), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n795), .A3(new_n791), .ZN(new_n796));
  INV_X1    g610(.A(new_n250), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n352), .B2(new_n369), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n738), .A2(KEYINPUT42), .ZN(new_n799));
  OR3_X1    g613(.A1(new_n796), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n793), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT111), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n793), .A2(new_n803), .A3(new_n800), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(new_n281), .ZN(G33));
  AND3_X1   g620(.A1(new_n794), .A2(new_n795), .A3(new_n791), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n807), .A2(new_n377), .A3(new_n715), .A4(new_n717), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G134), .ZN(G36));
  NAND2_X1  g623(.A1(new_n577), .A2(new_n537), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n576), .A2(new_n556), .A3(new_n573), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n741), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n578), .A2(KEYINPUT45), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n814), .A2(KEYINPUT112), .A3(new_n815), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(G469), .A2(G902), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(KEYINPUT46), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n818), .A2(new_n819), .B1(G469), .B2(G902), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(KEYINPUT113), .A3(KEYINPUT46), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n572), .B1(new_n825), .B2(KEYINPUT46), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n494), .A3(new_n720), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n723), .A2(new_n665), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT43), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n693), .B1(new_n655), .B2(new_n654), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n836), .A2(KEYINPUT44), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(KEYINPUT44), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT89), .B1(new_n635), .B2(new_n618), .ZN(new_n839));
  INV_X1    g653(.A(new_n614), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n603), .A2(new_n604), .A3(new_n612), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n601), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(G902), .B1(new_n844), .B2(new_n636), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n639), .B1(new_n845), .B2(new_n611), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n642), .A2(KEYINPUT90), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n645), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n647), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OR4_X1    g664(.A1(new_n831), .A2(new_n837), .A3(new_n838), .A4(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(G137), .ZN(G39));
  INV_X1    g666(.A(KEYINPUT47), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n830), .B2(new_n494), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n828), .B1(new_n824), .B2(new_n826), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n856), .A2(KEYINPUT114), .A3(new_n495), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n853), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n830), .A2(new_n854), .A3(new_n494), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT114), .B1(new_n856), .B2(new_n495), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n860), .A3(KEYINPUT47), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NOR4_X1   g676(.A1(new_n736), .A2(new_n797), .A3(new_n776), .A4(new_n850), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n862), .A2(KEYINPUT115), .A3(new_n863), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(G140), .ZN(G42));
  NOR4_X1   g683(.A1(new_n832), .A2(new_n730), .A3(new_n250), .A4(new_n790), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n757), .B(KEYINPUT49), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n871), .A3(new_n732), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT116), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n649), .A2(new_n580), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n377), .A2(new_n876), .A3(new_n493), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n646), .A2(new_n492), .A3(new_n648), .ZN(new_n878));
  INV_X1    g692(.A(new_n422), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n666), .B1(new_n485), .B2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n878), .A2(new_n880), .A3(new_n580), .A4(new_n657), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n695), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n875), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n650), .A2(KEYINPUT117), .A3(new_n695), .A4(new_n881), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n750), .A2(new_n774), .A3(new_n746), .ZN(new_n886));
  INV_X1    g700(.A(new_n761), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n753), .A2(new_n759), .A3(KEYINPUT106), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n771), .A2(new_n772), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n738), .A3(new_n702), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n796), .A2(new_n891), .ZN(new_n892));
  AND4_X1   g706(.A1(new_n420), .A2(new_n414), .A3(new_n421), .A4(new_n712), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(new_n682), .A3(new_n684), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n676), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n648), .B1(new_n643), .B2(new_n645), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT118), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n893), .A2(new_n682), .A3(new_n684), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n896), .A2(new_n898), .A3(KEYINPUT118), .A4(new_n710), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n892), .B1(new_n901), .B2(new_n704), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT119), .B1(new_n902), .B2(new_n808), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n788), .A2(new_n777), .A3(new_n791), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT118), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n705), .A2(new_n710), .A3(new_n893), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n905), .B1(new_n906), .B2(new_n850), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n907), .A2(new_n736), .A3(new_n737), .A4(new_n899), .ZN(new_n908));
  AND4_X1   g722(.A1(KEYINPUT119), .A2(new_n808), .A3(new_n904), .A4(new_n908), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n885), .B(new_n889), .C1(new_n903), .C2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n805), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT52), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n759), .A2(KEYINPUT108), .A3(new_n777), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n718), .B1(new_n913), .B2(new_n778), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n693), .A2(new_n494), .A3(new_n712), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n373), .B2(new_n729), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n788), .A2(new_n916), .A3(new_n667), .A4(new_n725), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n739), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n912), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n918), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n781), .A2(KEYINPUT52), .A3(new_n718), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n911), .A2(KEYINPUT53), .A3(new_n922), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n793), .A2(new_n803), .A3(new_n800), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n803), .B1(new_n793), .B2(new_n800), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI22_X1  g740(.A1(new_n773), .A2(new_n765), .B1(new_n377), .B2(new_n745), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n750), .B(new_n927), .C1(new_n760), .C2(new_n761), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n883), .B2(new_n884), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n715), .A2(new_n717), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n908), .B(new_n904), .C1(new_n792), .C2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT119), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n808), .A2(KEYINPUT119), .A3(new_n904), .A4(new_n908), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n922), .A2(new_n926), .A3(new_n929), .A4(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT53), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n874), .B1(new_n923), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n937), .B1(new_n793), .B2(new_n800), .ZN(new_n941));
  AND4_X1   g755(.A1(new_n885), .A2(new_n935), .A3(new_n889), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n922), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n938), .A2(new_n943), .ZN(new_n944));
  OAI22_X1  g758(.A1(new_n939), .A2(new_n940), .B1(new_n944), .B2(KEYINPUT54), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n834), .A2(new_n489), .A3(new_n773), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n946), .A2(new_n648), .A3(new_n732), .A4(new_n749), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT50), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n757), .A2(new_n495), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n858), .A2(new_n861), .A3(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n946), .A2(new_n896), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n730), .A2(new_n250), .A3(new_n488), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n850), .A2(new_n744), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n485), .A2(new_n665), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n834), .A2(new_n489), .A3(new_n954), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n890), .A2(new_n702), .ZN(new_n959));
  OAI22_X1  g773(.A1(new_n956), .A2(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n960), .A2(KEYINPUT121), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(KEYINPUT121), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n961), .A2(KEYINPUT51), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n952), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n486), .B1(new_n956), .B2(new_n666), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n958), .A2(new_n798), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT48), .ZN(new_n967));
  AOI211_X1 g781(.A(new_n965), .B(new_n967), .C1(new_n759), .C2(new_n946), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n960), .B(new_n948), .C1(new_n950), .C2(new_n951), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n964), .B(new_n968), .C1(new_n969), .C2(KEYINPUT51), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n939), .A2(new_n940), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n945), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(G952), .A2(G953), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n873), .B1(new_n972), .B2(new_n973), .ZN(G75));
  NOR2_X1   g788(.A1(new_n187), .A2(G952), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(G210), .A2(G902), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n944), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n602), .A2(new_n610), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(new_n608), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT55), .Z(new_n982));
  NOR2_X1   g796(.A1(new_n982), .A2(KEYINPUT56), .ZN(new_n983));
  AOI21_X1  g797(.A(KEYINPUT124), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT124), .ZN(new_n985));
  INV_X1    g799(.A(new_n983), .ZN(new_n986));
  AOI211_X1 g800(.A(new_n985), .B(new_n986), .C1(new_n944), .C2(new_n978), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n976), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  AOI22_X1  g802(.A1(new_n936), .A2(new_n937), .B1(new_n942), .B2(new_n922), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT122), .B1(new_n989), .B2(new_n977), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT122), .ZN(new_n991));
  AOI21_X1  g805(.A(KEYINPUT53), .B1(new_n911), .B2(new_n922), .ZN(new_n992));
  AND4_X1   g806(.A1(new_n922), .A2(new_n929), .A3(new_n935), .A4(new_n941), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n991), .B(new_n978), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT56), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n990), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n982), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(KEYINPUT123), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT123), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n996), .A2(new_n999), .A3(new_n982), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n988), .B1(new_n998), .B2(new_n1000), .ZN(G51));
  XNOR2_X1  g815(.A(new_n989), .B(KEYINPUT54), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n821), .B(KEYINPUT57), .ZN(new_n1003));
  OAI22_X1  g817(.A1(new_n1002), .A2(new_n1003), .B1(new_n553), .B2(new_n557), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n989), .A2(new_n236), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1005), .A2(new_n818), .A3(new_n819), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n975), .B1(new_n1004), .B2(new_n1006), .ZN(G54));
  NAND3_X1  g821(.A1(new_n1005), .A2(KEYINPUT58), .A3(G475), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n1008), .A2(new_n481), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1008), .A2(new_n481), .ZN(new_n1010));
  NOR3_X1   g824(.A1(new_n1009), .A2(new_n1010), .A3(new_n975), .ZN(G60));
  NAND2_X1  g825(.A1(G478), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT59), .Z(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n663), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n976), .B1(new_n1002), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1014), .B1(new_n945), .B2(new_n971), .ZN(new_n1017));
  INV_X1    g831(.A(new_n663), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(G63));
  NAND2_X1  g833(.A1(G217), .A2(G902), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT60), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n989), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g836(.A(KEYINPUT125), .B(new_n976), .C1(new_n1022), .C2(new_n246), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT61), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n976), .B1(new_n1022), .B2(new_n246), .ZN(new_n1026));
  INV_X1    g840(.A(new_n692), .ZN(new_n1027));
  NOR3_X1   g841(.A1(new_n989), .A2(new_n1027), .A3(new_n1021), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g844(.A(new_n1023), .B(new_n1024), .C1(new_n1026), .C2(new_n1028), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(new_n1031), .ZN(G66));
  NOR3_X1   g846(.A1(new_n491), .A2(new_n606), .A3(new_n187), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1033), .B1(new_n929), .B2(new_n187), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1034), .B(KEYINPUT126), .Z(new_n1035));
  OAI21_X1  g849(.A(new_n980), .B1(G898), .B2(new_n187), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1035), .B(new_n1036), .ZN(G69));
  NAND2_X1  g851(.A1(new_n338), .A2(new_n339), .ZN(new_n1038));
  XOR2_X1   g852(.A(new_n1038), .B(new_n473), .Z(new_n1039));
  NAND2_X1  g853(.A1(new_n1039), .A2(new_n535), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n187), .B1(new_n1040), .B2(G900), .ZN(new_n1041));
  NAND4_X1  g855(.A1(new_n377), .A2(new_n721), .A3(new_n896), .A4(new_n880), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n851), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(KEYINPUT127), .ZN(new_n1044));
  INV_X1    g858(.A(KEYINPUT127), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n851), .A2(new_n1045), .A3(new_n1042), .ZN(new_n1046));
  INV_X1    g860(.A(new_n914), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1047), .A2(new_n739), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1048), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1049), .A2(KEYINPUT62), .A3(new_n734), .ZN(new_n1050));
  INV_X1    g864(.A(KEYINPUT62), .ZN(new_n1051));
  INV_X1    g865(.A(new_n734), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1051), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g867(.A1(new_n1044), .A2(new_n1046), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1054), .A2(new_n868), .ZN(new_n1055));
  AND2_X1   g869(.A1(new_n1039), .A2(new_n187), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n1041), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OR3_X1    g871(.A1(new_n831), .A2(new_n764), .A3(new_n798), .ZN(new_n1058));
  AND3_X1   g872(.A1(new_n851), .A2(new_n1058), .A3(new_n1049), .ZN(new_n1059));
  AND2_X1   g873(.A1(new_n868), .A2(new_n1059), .ZN(new_n1060));
  AND3_X1   g874(.A1(new_n926), .A2(new_n187), .A3(new_n808), .ZN(new_n1061));
  AOI22_X1  g875(.A1(new_n1060), .A2(new_n1061), .B1(G227), .B2(G953), .ZN(new_n1062));
  OAI21_X1  g876(.A(new_n1057), .B1(new_n1062), .B2(new_n1039), .ZN(G72));
  NAND3_X1  g877(.A1(new_n1054), .A2(new_n868), .A3(new_n929), .ZN(new_n1064));
  NAND2_X1  g878(.A1(G472), .A2(G902), .ZN(new_n1065));
  XOR2_X1   g879(.A(new_n1065), .B(KEYINPUT63), .Z(new_n1066));
  AOI21_X1  g880(.A(new_n726), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g881(.A1(new_n343), .A2(new_n320), .A3(new_n258), .ZN(new_n1068));
  AND3_X1   g882(.A1(new_n926), .A2(new_n929), .A3(new_n808), .ZN(new_n1069));
  NAND3_X1  g883(.A1(new_n868), .A2(new_n1059), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n1068), .B1(new_n1070), .B2(new_n1066), .ZN(new_n1071));
  AND2_X1   g885(.A1(new_n923), .A2(new_n938), .ZN(new_n1072));
  NAND3_X1  g886(.A1(new_n726), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1073));
  OAI21_X1  g887(.A(new_n976), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NOR3_X1   g888(.A1(new_n1067), .A2(new_n1071), .A3(new_n1074), .ZN(G57));
endmodule


