//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024;
  XOR2_X1   g000(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G169gat), .B(G197gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT86), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G113gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n206), .B(G113gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(new_n211), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n203), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n211), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n208), .A2(new_n212), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(new_n218), .A3(new_n202), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n222));
  NAND2_X1  g021(.A1(G229gat), .A2(G233gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n226), .A2(G1gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n226), .B1(new_n228), .B2(G1gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT91), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(new_n226), .B2(G1gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(G8gat), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G8gat), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n227), .B(new_n229), .C1(new_n231), .C2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G29gat), .A2(G36gat), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n238));
  NOR3_X1   g037(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT88), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n242));
  INV_X1    g041(.A(G36gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n237), .B1(new_n241), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G50gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G43gat), .ZN(new_n248));
  INV_X1    g047(.A(G43gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G50gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n250), .A3(KEYINPUT15), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT89), .ZN(new_n254));
  NOR4_X1   g053(.A1(new_n254), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT89), .B1(new_n242), .B2(new_n243), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n238), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT15), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n249), .A2(G50gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n247), .A2(G43gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n257), .A2(new_n251), .A3(new_n237), .A4(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n253), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n236), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n233), .A2(new_n235), .B1(new_n253), .B2(new_n262), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n225), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n223), .ZN(new_n267));
  NAND2_X1  g066(.A1(KEYINPUT90), .A2(KEYINPUT17), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT90), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT17), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n261), .A2(new_n251), .A3(new_n237), .ZN(new_n272));
  INV_X1    g071(.A(new_n238), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT14), .ZN(new_n274));
  INV_X1    g073(.A(G29gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n275), .A3(new_n243), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(new_n254), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n242), .A2(KEYINPUT89), .A3(new_n243), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(KEYINPUT88), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(new_n244), .A3(new_n238), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n251), .B1(new_n282), .B2(new_n237), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n268), .B(new_n271), .C1(new_n280), .C2(new_n283), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n253), .A2(new_n262), .A3(new_n269), .A4(new_n270), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n236), .ZN(new_n287));
  AOI211_X1 g086(.A(new_n267), .B(new_n265), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n266), .B1(new_n288), .B2(KEYINPUT18), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n265), .B1(new_n286), .B2(new_n287), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(KEYINPUT18), .A3(new_n223), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n221), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n286), .A2(new_n287), .ZN(new_n294));
  INV_X1    g093(.A(new_n265), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n223), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT18), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n298), .A2(new_n220), .A3(new_n291), .A4(new_n266), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT93), .B1(G71gat), .B2(G78gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(G71gat), .A2(G78gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT94), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT9), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G57gat), .A2(G64gat), .ZN(new_n307));
  OR2_X1    g106(.A1(G57gat), .A2(G64gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n304), .B1(new_n303), .B2(new_n305), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n302), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(G71gat), .B(G78gat), .Z(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n312), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n314), .B(new_n302), .C1(new_n309), .C2(new_n310), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT95), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n313), .A2(KEYINPUT95), .A3(new_n315), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT21), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n287), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n322), .B(KEYINPUT96), .Z(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n324));
  INV_X1    g123(.A(G155gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n316), .A2(KEYINPUT21), .ZN(new_n329));
  AND2_X1   g128(.A1(G231gat), .A2(G233gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G127gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G183gat), .B(G211gat), .Z(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n331), .B(G127gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n334), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n322), .B(KEYINPUT96), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n326), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n328), .A2(new_n335), .A3(new_n338), .A4(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n328), .A2(new_n340), .B1(new_n335), .B2(new_n338), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(G232gat), .A2(G233gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n345), .A2(KEYINPUT41), .ZN(new_n346));
  XNOR2_X1  g145(.A(G134gat), .B(G162gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G85gat), .A2(G92gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT7), .ZN(new_n351));
  NAND2_X1  g150(.A1(G99gat), .A2(G106gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT8), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT97), .ZN(new_n354));
  OR2_X1    g153(.A1(G85gat), .A2(G92gat), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n354), .B1(new_n353), .B2(new_n355), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n351), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(G99gat), .B(G106gat), .Z(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n359), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n361), .B(new_n351), .C1(new_n356), .C2(new_n357), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n286), .A2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(G190gat), .B(G218gat), .Z(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n360), .A2(new_n362), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n367), .A2(new_n263), .B1(KEYINPUT41), .B2(new_n345), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n366), .B1(new_n364), .B2(new_n368), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n349), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n371), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(new_n369), .A3(new_n348), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT98), .B1(new_n344), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n343), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n341), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT98), .ZN(new_n379));
  INV_X1    g178(.A(new_n375), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G230gat), .ZN(new_n382));
  INV_X1    g181(.A(G233gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT99), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n362), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n316), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n367), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n313), .A2(new_n315), .B1(new_n362), .B2(new_n386), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n363), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT10), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n360), .A2(KEYINPUT10), .A3(new_n362), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n393), .B1(new_n318), .B2(new_n319), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n385), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n389), .A2(new_n384), .A3(new_n391), .ZN(new_n396));
  XNOR2_X1  g195(.A(G120gat), .B(G148gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(G176gat), .B(G204gat), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n397), .B(new_n398), .Z(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n395), .B2(new_n396), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n376), .A2(new_n381), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT76), .ZN(new_n406));
  INV_X1    g205(.A(G120gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n207), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT1), .ZN(new_n409));
  NAND2_X1  g208(.A1(G113gat), .A2(G120gat), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n332), .A2(KEYINPUT68), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT68), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(G127gat), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n412), .A2(new_n414), .A3(G134gat), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT67), .B1(new_n332), .B2(G134gat), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT67), .ZN(new_n417));
  INV_X1    g216(.A(G134gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n418), .A3(G127gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n411), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  XOR2_X1   g220(.A(G141gat), .B(G148gat), .Z(new_n422));
  XNOR2_X1  g221(.A(G155gat), .B(G162gat), .ZN(new_n423));
  INV_X1    g222(.A(G162gat), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n325), .A2(KEYINPUT75), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT75), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(G155gat), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n424), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT2), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n422), .B(new_n423), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n423), .ZN(new_n431));
  OR2_X1    g230(.A1(G141gat), .A2(G148gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(G141gat), .A2(G148gat), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n410), .ZN(new_n436));
  NOR2_X1   g235(.A1(G113gat), .A2(G120gat), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT69), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT69), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n408), .A2(new_n439), .A3(new_n410), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n332), .A2(G134gat), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT1), .B1(new_n418), .B2(G127gat), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n438), .A2(new_n440), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n421), .A2(new_n430), .A3(new_n435), .A4(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n421), .A2(new_n443), .B1(new_n430), .B2(new_n435), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n406), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT78), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT5), .ZN(new_n449));
  INV_X1    g248(.A(new_n406), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n421), .A2(new_n443), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n425), .A2(new_n427), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n429), .B1(new_n452), .B2(G162gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n422), .A2(new_n423), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n435), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n450), .B1(new_n456), .B2(new_n444), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT5), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT78), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n451), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n423), .A2(new_n432), .A3(new_n433), .ZN(new_n461));
  XNOR2_X1  g260(.A(KEYINPUT75), .B(G155gat), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT2), .B1(new_n462), .B2(new_n424), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n461), .A2(new_n463), .B1(new_n434), .B2(new_n431), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n460), .A2(KEYINPUT4), .A3(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n444), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n455), .A2(KEYINPUT3), .B1(new_n421), .B2(new_n443), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n406), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n449), .A2(new_n459), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G1gat), .B(G29gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT0), .ZN(new_n475));
  XNOR2_X1  g274(.A(G57gat), .B(G85gat), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n475), .B(new_n476), .Z(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n444), .A2(new_n466), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n479), .B(new_n458), .C1(KEYINPUT4), .C2(new_n445), .ZN(new_n480));
  INV_X1    g279(.A(new_n472), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n473), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT79), .B1(new_n483), .B2(KEYINPUT6), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n478), .B1(new_n473), .B2(new_n482), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n449), .A2(new_n459), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n472), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n482), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n489), .A3(new_n477), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT79), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n484), .A2(new_n485), .A3(new_n493), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n485), .A2(new_n492), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G8gat), .B(G36gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(G64gat), .B(G92gat), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n497), .B(new_n498), .Z(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G197gat), .B(G204gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT22), .ZN(new_n502));
  INV_X1    g301(.A(G211gat), .ZN(new_n503));
  INV_X1    g302(.A(G218gat), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G211gat), .B(G218gat), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n501), .A3(new_n505), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G226gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(new_n383), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT25), .ZN(new_n515));
  NAND2_X1  g314(.A1(G183gat), .A2(G190gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT24), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT24), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(G183gat), .A3(G190gat), .ZN(new_n519));
  INV_X1    g318(.A(G183gat), .ZN(new_n520));
  INV_X1    g319(.A(G190gat), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n517), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(G169gat), .A2(G176gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT23), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT23), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(G169gat), .B2(G176gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(G169gat), .A2(G176gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n515), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n526), .A2(KEYINPUT25), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n517), .A2(new_n519), .ZN(new_n531));
  NAND2_X1  g330(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n533), .A2(new_n534), .A3(G190gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n530), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT64), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n525), .A2(G169gat), .A3(G176gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n527), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n524), .A2(KEYINPUT64), .A3(new_n527), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n529), .B1(new_n536), .B2(new_n542), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n539), .A2(new_n523), .A3(KEYINPUT26), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n523), .A2(KEYINPUT26), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n516), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  OR2_X1    g346(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n548), .A2(KEYINPUT27), .A3(new_n532), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT27), .ZN(new_n550));
  AOI211_X1 g349(.A(KEYINPUT28), .B(G190gat), .C1(new_n550), .C2(G183gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(G183gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n520), .A2(KEYINPUT27), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n553), .A3(new_n521), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n549), .A2(new_n551), .B1(new_n554), .B2(KEYINPUT28), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n547), .B1(new_n555), .B2(KEYINPUT66), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n549), .A2(new_n551), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT28), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT27), .B(G183gat), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(new_n559), .B2(new_n521), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT66), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n557), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n543), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT29), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n514), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n514), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n561), .B1(new_n557), .B2(new_n560), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n555), .A2(KEYINPUT66), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n547), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n566), .B1(new_n569), .B2(new_n543), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n512), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n563), .A2(new_n514), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT29), .B1(new_n569), .B2(new_n543), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n572), .B(new_n511), .C1(new_n573), .C2(new_n514), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n571), .A2(KEYINPUT72), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT72), .B1(new_n571), .B2(new_n574), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n500), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n571), .A2(new_n499), .A3(new_n574), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT30), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT74), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT73), .B(KEYINPUT30), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n578), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n581), .B1(new_n578), .B2(new_n582), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n577), .B(new_n580), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n496), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT29), .B1(new_n509), .B2(new_n510), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT81), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n470), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI211_X1 g389(.A(KEYINPUT81), .B(KEYINPUT29), .C1(new_n509), .C2(new_n510), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n455), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n471), .A2(new_n564), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(new_n512), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G228gat), .A2(G233gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n596), .B(KEYINPUT80), .Z(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G22gat), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n596), .B1(new_n455), .B2(KEYINPUT3), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n511), .A2(new_n564), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n600), .B1(new_n464), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n511), .B1(new_n471), .B2(new_n564), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n598), .A2(new_n599), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n597), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n607), .B1(new_n592), .B2(new_n594), .ZN(new_n608));
  OAI21_X1  g407(.A(G22gat), .B1(new_n608), .B2(new_n604), .ZN(new_n609));
  INV_X1    g408(.A(G78gat), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n606), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n610), .B1(new_n606), .B2(new_n609), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT31), .B(G50gat), .ZN(new_n613));
  INV_X1    g412(.A(G106gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n611), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n599), .B1(new_n598), .B2(new_n605), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n608), .A2(new_n604), .A3(G22gat), .ZN(new_n619));
  OAI21_X1  g418(.A(G78gat), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n606), .A2(new_n609), .A3(new_n610), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n615), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n587), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n563), .A2(new_n460), .ZN(new_n626));
  AND2_X1   g425(.A1(G227gat), .A2(G233gat), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n569), .A2(new_n451), .A3(new_n543), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT32), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G15gat), .B(G43gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(G71gat), .B(G99gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n634), .B1(new_n639), .B2(new_n635), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT70), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n639), .A2(new_n641), .A3(KEYINPUT32), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n641), .B1(new_n639), .B2(KEYINPUT32), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT71), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI211_X1 g445(.A(KEYINPUT71), .B(new_n640), .C1(new_n642), .C2(new_n643), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n638), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n626), .A2(new_n628), .ZN(new_n649));
  OR3_X1    g448(.A1(new_n649), .A2(KEYINPUT34), .A3(new_n627), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT34), .B1(new_n649), .B2(new_n627), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  AOI211_X1 g453(.A(new_n652), .B(new_n638), .C1(new_n646), .C2(new_n647), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT36), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT70), .B1(new_n629), .B2(new_n630), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n639), .A2(new_n641), .A3(KEYINPUT32), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT71), .B1(new_n660), .B2(new_n640), .ZN(new_n661));
  INV_X1    g460(.A(new_n647), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n637), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n652), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n653), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT36), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n625), .B1(new_n657), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT82), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n625), .B(KEYINPUT82), .C1(new_n657), .C2(new_n666), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT83), .B(KEYINPUT37), .Z(new_n671));
  NAND3_X1  g470(.A1(new_n571), .A2(new_n574), .A3(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n672), .A2(new_n500), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n571), .A2(new_n574), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT38), .B1(new_n674), .B2(KEYINPUT37), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n579), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n490), .A2(new_n485), .A3(new_n492), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(new_n495), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT38), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT37), .B1(new_n575), .B2(new_n576), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n680), .B2(new_n673), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n623), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n469), .A2(new_n471), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n683), .B(new_n479), .C1(KEYINPUT4), .C2(new_n445), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n406), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n456), .A2(new_n450), .A3(new_n444), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n685), .A2(KEYINPUT39), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n477), .B1(new_n685), .B2(KEYINPUT39), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT40), .ZN(new_n689));
  OR3_X1    g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n687), .B2(new_n688), .ZN(new_n691));
  AND4_X1   g490(.A1(new_n485), .A2(new_n585), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n682), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n669), .A2(new_n670), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n664), .A2(new_n623), .A3(new_n665), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT35), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n495), .A2(new_n677), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n586), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n585), .B1(new_n494), .B2(new_n495), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n701), .A2(new_n664), .A3(new_n665), .A4(new_n623), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n702), .A2(KEYINPUT84), .A3(KEYINPUT35), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT84), .B1(new_n702), .B2(KEYINPUT35), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n700), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI211_X1 g504(.A(new_n301), .B(new_n404), .C1(new_n694), .C2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n496), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g508(.A1(new_n706), .A2(new_n585), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n228), .A2(new_n234), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n234), .B2(new_n711), .ZN(new_n715));
  MUX2_X1   g514(.A(new_n714), .B(new_n715), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g515(.A(new_n656), .B1(new_n654), .B2(new_n655), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n664), .A2(KEYINPUT36), .A3(new_n665), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT101), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n717), .B2(new_n718), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n706), .A2(G15gat), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n654), .A2(new_n655), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n706), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(G15gat), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n726), .A2(KEYINPUT100), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT100), .B1(new_n726), .B2(new_n727), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n724), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT102), .ZN(G1326gat));
  NAND2_X1  g530(.A1(new_n706), .A2(new_n624), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT43), .B(G22gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1327gat));
  OAI21_X1  g533(.A(KEYINPUT101), .B1(new_n657), .B2(new_n666), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n735), .A2(new_n693), .A3(new_n625), .A4(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n380), .B1(new_n705), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n380), .B1(new_n694), .B2(new_n705), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n403), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n378), .A2(new_n301), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G29gat), .B1(new_n745), .B2(new_n496), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n741), .A2(new_n744), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n747), .A2(G29gat), .A3(new_n496), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT103), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n749), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n751), .B1(new_n750), .B2(new_n752), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n746), .B1(new_n753), .B2(new_n754), .ZN(G1328gat));
  INV_X1    g554(.A(new_n747), .ZN(new_n756));
  AOI21_X1  g555(.A(G36gat), .B1(KEYINPUT104), .B2(KEYINPUT46), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n756), .A2(new_n585), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G36gat), .B1(new_n745), .B2(new_n586), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(G1329gat));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(KEYINPUT47), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n741), .A2(new_n249), .A3(new_n725), .A4(new_n744), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n765), .A2(KEYINPUT105), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(KEYINPUT105), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n745), .A2(new_n722), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n769), .B2(new_n249), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n763), .A2(KEYINPUT47), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT107), .Z(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n768), .B(new_n772), .C1(new_n769), .C2(new_n249), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(G1330gat));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n623), .B1(new_n756), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n747), .A2(KEYINPUT108), .ZN(new_n779));
  AOI21_X1  g578(.A(G50gat), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n624), .A2(G50gat), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n745), .A2(new_n781), .ZN(new_n782));
  OR3_X1    g581(.A1(new_n780), .A2(new_n782), .A3(KEYINPUT48), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT48), .B1(new_n780), .B2(new_n782), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1331gat));
  NAND4_X1  g584(.A1(new_n376), .A2(new_n301), .A3(new_n381), .A4(new_n743), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n705), .B2(new_n737), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n707), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n585), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n791));
  XOR2_X1   g590(.A(KEYINPUT49), .B(G64gat), .Z(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n790), .B2(new_n792), .ZN(G1333gat));
  NAND2_X1  g592(.A1(new_n787), .A2(new_n723), .ZN(new_n794));
  INV_X1    g593(.A(new_n725), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(G71gat), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n794), .A2(G71gat), .B1(new_n787), .B2(new_n796), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g597(.A1(new_n787), .A2(new_n624), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g599(.A1(new_n378), .A2(new_n300), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(new_n403), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n694), .A2(new_n705), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n739), .B1(new_n804), .B2(new_n375), .ZN(new_n805));
  AOI211_X1 g604(.A(KEYINPUT44), .B(new_n380), .C1(new_n705), .C2(new_n737), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n707), .B(new_n803), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT109), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT109), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n742), .A2(new_n809), .A3(new_n707), .A4(new_n803), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(new_n810), .A3(G85gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT35), .B1(new_n695), .B2(new_n587), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT84), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n702), .A2(KEYINPUT84), .A3(KEYINPUT35), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n699), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n682), .A2(new_n692), .B1(new_n701), .B2(new_n623), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n720), .A2(new_n721), .A3(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(KEYINPUT110), .B(new_n375), .C1(new_n820), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n801), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n705), .A2(new_n737), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT110), .B1(new_n825), .B2(new_n375), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n812), .B(new_n815), .C1(new_n824), .C2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n802), .B1(new_n738), .B2(KEYINPUT110), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n375), .B1(new_n820), .B2(new_n822), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT110), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n828), .A2(new_n813), .A3(new_n814), .A4(new_n831), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n496), .A2(G85gat), .A3(new_n403), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n827), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n811), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT112), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n811), .A2(new_n837), .A3(new_n834), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(G1336gat));
  AND2_X1   g638(.A1(new_n827), .A2(new_n832), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n586), .A2(G92gat), .A3(new_n403), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n742), .A2(new_n803), .ZN(new_n844));
  OAI21_X1  g643(.A(G92gat), .B1(new_n844), .B2(new_n586), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n842), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT113), .B1(new_n824), .B2(new_n826), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n814), .ZN(new_n848));
  OAI211_X1 g647(.A(KEYINPUT113), .B(KEYINPUT51), .C1(new_n824), .C2(new_n826), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n849), .A3(new_n841), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n850), .A2(new_n845), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n846), .B1(new_n851), .B2(new_n843), .ZN(G1337gat));
  NOR2_X1   g651(.A1(new_n795), .A2(G99gat), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n840), .A2(new_n743), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(G99gat), .B1(new_n844), .B2(new_n722), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1338gat));
  NOR2_X1   g655(.A1(new_n623), .A2(G106gat), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n840), .A2(KEYINPUT114), .A3(new_n743), .A4(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n827), .A2(new_n832), .A3(new_n743), .A4(new_n857), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n742), .A2(new_n624), .A3(new_n803), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT53), .B1(new_n862), .B2(G106gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n858), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n623), .A2(G106gat), .A3(new_n403), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n848), .A2(new_n849), .A3(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n862), .A2(G106gat), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT53), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n864), .A2(new_n868), .ZN(G1339gat));
  NAND4_X1  g668(.A1(new_n376), .A2(new_n301), .A3(new_n381), .A4(new_n403), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n290), .A2(new_n223), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n264), .A2(new_n265), .A3(new_n225), .ZN(new_n872));
  OAI22_X1  g671(.A1(new_n871), .A2(new_n872), .B1(new_n213), .B2(new_n215), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n299), .B(new_n873), .C1(new_n401), .C2(new_n402), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT55), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT10), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n363), .A2(new_n316), .A3(new_n387), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n390), .A2(new_n363), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n394), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n384), .A3(new_n880), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n395), .A2(new_n881), .A3(KEYINPUT54), .ZN(new_n882));
  XNOR2_X1  g681(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n385), .B(new_n883), .C1(new_n392), .C2(new_n394), .ZN(new_n884));
  INV_X1    g683(.A(new_n399), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n875), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n300), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n395), .A2(new_n881), .A3(KEYINPUT54), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n889), .A2(KEYINPUT55), .A3(new_n885), .A4(new_n884), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n400), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n874), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n380), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n887), .A2(new_n375), .A3(new_n400), .A4(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n299), .A2(new_n873), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT116), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT116), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n299), .A2(new_n897), .A3(new_n873), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n893), .B1(new_n894), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n344), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n870), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(new_n695), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n707), .A3(new_n586), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(new_n207), .A3(new_n301), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n707), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n906), .A2(KEYINPUT117), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(KEYINPUT117), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n586), .A3(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n300), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n905), .B1(new_n911), .B2(new_n207), .ZN(G1340gat));
  OAI21_X1  g711(.A(G120gat), .B1(new_n904), .B2(new_n403), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n743), .A2(new_n407), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT118), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT118), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n913), .B(new_n917), .C1(new_n909), .C2(new_n914), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1341gat));
  NAND2_X1  g718(.A1(new_n412), .A2(new_n414), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n904), .B2(new_n344), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n378), .A2(new_n412), .A3(new_n414), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n909), .B2(new_n922), .ZN(G1342gat));
  NOR2_X1   g722(.A1(new_n380), .A2(G134gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n910), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT56), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT56), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n910), .A2(new_n927), .A3(new_n924), .ZN(new_n928));
  OAI21_X1  g727(.A(G134gat), .B1(new_n904), .B2(new_n380), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(G1343gat));
  NOR2_X1   g729(.A1(new_n496), .A2(new_n585), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n722), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n902), .A2(new_n623), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT57), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n902), .A2(new_n935), .A3(new_n623), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n932), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n210), .B1(new_n939), .B2(new_n300), .ZN(new_n940));
  INV_X1    g739(.A(new_n932), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n933), .A2(new_n941), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n942), .A2(G141gat), .A3(new_n301), .ZN(new_n943));
  XNOR2_X1  g742(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  OR3_X1    g744(.A1(new_n940), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n940), .B2(new_n943), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1344gat));
  NAND2_X1  g747(.A1(new_n939), .A2(new_n743), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT59), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n949), .A2(new_n950), .A3(G148gat), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n932), .A2(new_n403), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n899), .B1(new_n894), .B2(KEYINPUT120), .ZN(new_n953));
  INV_X1    g752(.A(new_n891), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n954), .A2(new_n955), .A3(new_n375), .A4(new_n887), .ZN(new_n956));
  AOI22_X1  g755(.A1(new_n953), .A2(new_n956), .B1(new_n892), .B2(new_n380), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT121), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n344), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n953), .A2(new_n956), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n960), .A2(new_n958), .A3(new_n893), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n870), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n623), .B1(new_n962), .B2(KEYINPUT122), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n870), .B(new_n964), .C1(new_n959), .C2(new_n961), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT57), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n952), .B1(new_n966), .B2(new_n937), .ZN(new_n967));
  AOI211_X1 g766(.A(KEYINPUT123), .B(new_n950), .C1(new_n967), .C2(G148gat), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n962), .A2(KEYINPUT122), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n970), .A2(new_n624), .A3(new_n965), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n937), .B1(new_n971), .B2(new_n935), .ZN(new_n972));
  INV_X1    g771(.A(new_n952), .ZN(new_n973));
  OAI21_X1  g772(.A(G148gat), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n969), .B1(new_n974), .B2(KEYINPUT59), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n951), .B1(new_n968), .B2(new_n975), .ZN(new_n976));
  OR3_X1    g775(.A1(new_n934), .A2(new_n973), .A3(G148gat), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1345gat));
  INV_X1    g777(.A(new_n942), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n452), .B1(new_n979), .B2(new_n378), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n344), .A2(new_n462), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n980), .B1(new_n939), .B2(new_n981), .ZN(G1346gat));
  NAND3_X1  g781(.A1(new_n979), .A2(new_n424), .A3(new_n375), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n939), .A2(new_n375), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n983), .B1(new_n984), .B2(new_n424), .ZN(G1347gat));
  INV_X1    g784(.A(G169gat), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n707), .A2(new_n586), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n903), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n986), .B1(new_n988), .B2(new_n300), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n989), .B(KEYINPUT124), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n988), .A2(new_n986), .A3(new_n300), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1348gat));
  NAND2_X1  g791(.A1(new_n988), .A2(new_n743), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n993), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g793(.A1(new_n988), .A2(new_n378), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n995), .A2(new_n548), .A3(new_n532), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n996), .B1(new_n559), .B2(new_n995), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT60), .ZN(new_n998));
  XNOR2_X1  g797(.A(new_n997), .B(new_n998), .ZN(G1350gat));
  NOR2_X1   g798(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n1000));
  AOI21_X1  g799(.A(new_n1000), .B1(new_n988), .B2(new_n375), .ZN(new_n1001));
  NAND2_X1  g800(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n1002));
  XOR2_X1   g801(.A(new_n1001), .B(new_n1002), .Z(G1351gat));
  NAND3_X1  g802(.A1(new_n933), .A2(new_n722), .A3(new_n987), .ZN(new_n1004));
  INV_X1    g803(.A(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g804(.A(KEYINPUT125), .B(G197gat), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n1005), .A2(new_n300), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n722), .A2(new_n987), .ZN(new_n1008));
  NOR3_X1   g807(.A1(new_n972), .A2(new_n301), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1007), .B1(new_n1009), .B2(new_n1006), .ZN(G1352gat));
  XNOR2_X1  g809(.A(KEYINPUT126), .B(G204gat), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1005), .A2(new_n743), .A3(new_n1011), .ZN(new_n1012));
  XOR2_X1   g811(.A(new_n1012), .B(KEYINPUT62), .Z(new_n1013));
  NOR3_X1   g812(.A1(new_n972), .A2(new_n403), .A3(new_n1008), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1013), .B1(new_n1014), .B2(new_n1011), .ZN(G1353gat));
  NAND3_X1  g814(.A1(new_n1005), .A2(new_n503), .A3(new_n378), .ZN(new_n1016));
  NOR2_X1   g815(.A1(new_n972), .A2(new_n1008), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1017), .A2(new_n378), .ZN(new_n1018));
  AND3_X1   g817(.A1(new_n1018), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1019));
  AOI21_X1  g818(.A(KEYINPUT63), .B1(new_n1018), .B2(G211gat), .ZN(new_n1020));
  OAI21_X1  g819(.A(new_n1016), .B1(new_n1019), .B2(new_n1020), .ZN(G1354gat));
  AOI21_X1  g820(.A(G218gat), .B1(new_n1005), .B2(new_n375), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n375), .A2(G218gat), .ZN(new_n1023));
  XNOR2_X1  g822(.A(new_n1023), .B(KEYINPUT127), .ZN(new_n1024));
  AOI21_X1  g823(.A(new_n1022), .B1(new_n1017), .B2(new_n1024), .ZN(G1355gat));
endmodule


