//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT70), .B(KEYINPUT32), .Z(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT68), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G953), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G237), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(G210), .A3(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n195), .B(KEYINPUT27), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT26), .B(G101), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  OR2_X1    g013(.A1(new_n195), .A2(KEYINPUT27), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(KEYINPUT27), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(new_n197), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT0), .A4(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n206), .A2(G146), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n204), .A2(G143), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT0), .B(G128), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n208), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  INV_X1    g028(.A(G134), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n214), .A2(new_n215), .A3(G137), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(KEYINPUT64), .A2(G134), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT64), .A2(G134), .ZN(new_n219));
  INV_X1    g033(.A(G137), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n217), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n215), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT64), .A2(G134), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n225), .A2(new_n222), .A3(G137), .A4(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(G137), .B1(new_n225), .B2(new_n226), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(KEYINPUT11), .ZN(new_n229));
  OAI21_X1  g043(.A(G131), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n225), .A2(G137), .A3(new_n226), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n216), .B1(new_n231), .B2(KEYINPUT65), .ZN(new_n232));
  INV_X1    g046(.A(G131), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n220), .B1(new_n218), .B2(new_n219), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n214), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n232), .A2(new_n233), .A3(new_n227), .A4(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n213), .B1(new_n230), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT1), .B1(new_n206), .B2(G146), .ZN(new_n238));
  OAI211_X1 g052(.A(G128), .B(new_n238), .C1(new_n209), .C2(new_n210), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n205), .B(new_n207), .C1(KEYINPUT1), .C2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n215), .A2(G137), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n233), .B1(new_n234), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n245), .A2(new_n236), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n237), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G119), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G116), .ZN(new_n249));
  INV_X1    g063(.A(G116), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G119), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT2), .B(G113), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n253), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n257), .B(KEYINPUT67), .Z(new_n258));
  AOI21_X1  g072(.A(new_n203), .B1(new_n247), .B2(new_n258), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n245), .A2(new_n236), .A3(KEYINPUT66), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n237), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n245), .A2(new_n236), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT30), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n213), .ZN(new_n266));
  INV_X1    g080(.A(new_n236), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n221), .A2(new_n222), .B1(new_n234), .B2(new_n214), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n233), .B1(new_n268), .B2(new_n232), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n266), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT30), .A3(new_n262), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n257), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n259), .B1(new_n265), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT31), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n259), .B(KEYINPUT31), .C1(new_n265), .C2(new_n272), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n247), .A2(new_n258), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n245), .A2(new_n236), .A3(KEYINPUT66), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n270), .A2(new_n264), .A3(new_n280), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n281), .A2(new_n257), .B1(new_n247), .B2(new_n258), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n283));
  OAI21_X1  g097(.A(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n275), .A2(new_n276), .B1(new_n203), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(G472), .A2(G902), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n188), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n284), .A2(new_n203), .ZN(new_n289));
  INV_X1    g103(.A(new_n276), .ZN(new_n290));
  INV_X1    g104(.A(new_n257), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n291), .B1(new_n247), .B2(KEYINPUT30), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT30), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n281), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT31), .B1(new_n295), .B2(new_n259), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n289), .B1(new_n290), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(KEYINPUT32), .A3(new_n286), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n288), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G472), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT71), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n292), .A2(new_n294), .B1(new_n247), .B2(new_n258), .ZN(new_n302));
  INV_X1    g116(.A(new_n203), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n277), .B1(new_n265), .B2(new_n272), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(KEYINPUT71), .A3(new_n203), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n303), .B(new_n279), .C1(new_n282), .C2(new_n283), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n304), .A2(new_n306), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n279), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n257), .B(KEYINPUT67), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n311), .B1(new_n237), .B2(new_n246), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n278), .B1(new_n277), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n203), .A2(new_n307), .ZN(new_n315));
  AOI21_X1  g129(.A(G902), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n300), .B1(new_n309), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n187), .B1(new_n299), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n309), .A2(new_n316), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G472), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n320), .A2(KEYINPUT72), .A3(new_n298), .A4(new_n288), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n213), .A2(G125), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n239), .A2(new_n241), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(G125), .ZN(new_n325));
  INV_X1    g139(.A(G224), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT7), .B1(new_n326), .B2(G953), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G101), .ZN(new_n329));
  INV_X1    g143(.A(G104), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G107), .ZN(new_n331));
  INV_X1    g145(.A(G107), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G104), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n329), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(KEYINPUT80), .A3(G104), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n332), .A2(KEYINPUT80), .A3(KEYINPUT3), .A4(G104), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n332), .A2(G104), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(G101), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n334), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n249), .A2(new_n251), .A3(KEYINPUT5), .ZN(new_n343));
  OAI21_X1  g157(.A(G113), .B1(new_n249), .B2(KEYINPUT5), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n342), .B1(new_n254), .B2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G110), .B(G122), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(KEYINPUT8), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT84), .B1(new_n343), .B2(new_n344), .ZN(new_n349));
  INV_X1    g163(.A(G113), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n250), .A2(G119), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT5), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n353), .B(new_n354), .C1(new_n352), .C2(new_n252), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n349), .A2(new_n355), .A3(new_n255), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n346), .B(new_n348), .C1(new_n356), .C2(new_n342), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n325), .A2(new_n327), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n328), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n360), .B1(new_n339), .B2(new_n341), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n340), .B1(new_n337), .B2(new_n338), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n361), .B1(new_n329), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n362), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n360), .A2(G101), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n363), .A2(new_n367), .A3(new_n257), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n342), .A2(new_n255), .A3(new_n349), .A4(new_n355), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(new_n347), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n359), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G902), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n347), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n252), .A2(new_n253), .ZN(new_n375));
  OAI22_X1  g189(.A1(new_n362), .A2(new_n365), .B1(new_n375), .B2(new_n254), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n364), .A2(G101), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n376), .B1(new_n377), .B2(new_n361), .ZN(new_n378));
  INV_X1    g192(.A(new_n369), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n374), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(KEYINPUT6), .A3(new_n370), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n326), .A2(G953), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n325), .B(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n384), .B(new_n374), .C1(new_n378), .C2(new_n379), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n381), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT85), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n381), .A2(KEYINPUT85), .A3(new_n383), .A4(new_n385), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n373), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(G210), .B1(G237), .B2(G902), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n391), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(new_n390), .B2(KEYINPUT86), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT86), .ZN(new_n395));
  AOI211_X1 g209(.A(new_n395), .B(new_n373), .C1(new_n388), .C2(new_n389), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n392), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G214), .B1(G237), .B2(G902), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT20), .ZN(new_n400));
  XNOR2_X1  g214(.A(G113), .B(G122), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(new_n330), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n193), .A2(G143), .A3(G214), .A4(new_n194), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n190), .A2(new_n192), .A3(G214), .A4(new_n194), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n206), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n407), .A2(KEYINPUT87), .A3(KEYINPUT18), .A4(G131), .ZN(new_n408));
  NAND3_X1  g222(.A1(KEYINPUT87), .A2(KEYINPUT18), .A3(G131), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n404), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G140), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G125), .ZN(new_n412));
  INV_X1    g226(.A(G125), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G140), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G146), .ZN(new_n416));
  XNOR2_X1  g230(.A(G125), .B(G140), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n204), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT88), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n416), .A2(new_n418), .A3(KEYINPUT88), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n408), .A2(new_n410), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n412), .A2(new_n414), .A3(KEYINPUT16), .ZN(new_n425));
  OR3_X1    g239(.A1(new_n413), .A2(KEYINPUT16), .A3(G140), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n425), .A2(G146), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n415), .B(KEYINPUT19), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n428), .B1(new_n429), .B2(G146), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n407), .A2(G131), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n404), .A2(new_n233), .A3(new_n406), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n403), .B1(new_n424), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n408), .A2(new_n410), .A3(new_n423), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT17), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n431), .A2(new_n436), .A3(new_n432), .ZN(new_n437));
  AOI21_X1  g251(.A(G146), .B1(new_n425), .B2(new_n426), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n427), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n439), .B1(new_n431), .B2(new_n436), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n402), .B(new_n435), .C1(new_n437), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(G475), .A2(G902), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n443), .B(KEYINPUT89), .Z(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n400), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  AOI211_X1 g260(.A(KEYINPUT20), .B(new_n444), .C1(new_n434), .C2(new_n441), .ZN(new_n447));
  INV_X1    g261(.A(G475), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n435), .B1(new_n437), .B2(new_n440), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n403), .ZN(new_n450));
  AOI21_X1  g264(.A(G902), .B1(new_n450), .B2(new_n441), .ZN(new_n451));
  OAI22_X1  g265(.A1(new_n446), .A2(new_n447), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n206), .A2(G128), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n240), .A2(G143), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n225), .A2(new_n226), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n455), .B(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G116), .B(G122), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n332), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n250), .A2(KEYINPUT14), .A3(G122), .ZN(new_n460));
  INV_X1    g274(.A(new_n458), .ZN(new_n461));
  OAI211_X1 g275(.A(G107), .B(new_n460), .C1(new_n461), .C2(KEYINPUT14), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n457), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n458), .B(new_n332), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT13), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n453), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n454), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n453), .A2(new_n465), .ZN(new_n468));
  OAI21_X1  g282(.A(G134), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OR2_X1    g283(.A1(new_n456), .A2(new_n455), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n464), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n463), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT9), .B(G234), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(G217), .A3(new_n189), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n475), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n463), .A2(new_n471), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(G902), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT90), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G478), .ZN(new_n485));
  NOR2_X1   g299(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT92), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n490), .B1(new_n479), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n479), .A2(KEYINPUT92), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n484), .A2(new_n492), .B1(new_n493), .B2(new_n490), .ZN(new_n494));
  INV_X1    g308(.A(G952), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(G953), .ZN(new_n496));
  INV_X1    g310(.A(G234), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n496), .B1(new_n497), .B2(new_n194), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n372), .B(new_n193), .C1(G234), .C2(G237), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT21), .B(G898), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n452), .A2(new_n494), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G221), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(new_n474), .B2(new_n372), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G469), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n193), .A2(G227), .ZN(new_n508));
  XOR2_X1   g322(.A(G110), .B(G140), .Z(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n363), .A2(new_n367), .A3(new_n266), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n324), .A2(new_n342), .A3(KEYINPUT10), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n330), .A2(G107), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT3), .B1(new_n514), .B2(KEYINPUT80), .ZN(new_n515));
  INV_X1    g329(.A(new_n338), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n341), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n334), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n517), .A2(new_n241), .A3(new_n239), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT81), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT81), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n324), .A2(new_n342), .A3(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT82), .B(KEYINPUT10), .Z(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT83), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT83), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n520), .A2(new_n526), .A3(new_n522), .A4(new_n523), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n513), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n230), .A2(new_n236), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n510), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n513), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n324), .A2(new_n342), .A3(new_n521), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n521), .B1(new_n324), .B2(new_n342), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n526), .B1(new_n535), .B2(new_n523), .ZN(new_n536));
  INV_X1    g350(.A(new_n527), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n529), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n531), .A2(new_n539), .ZN(new_n540));
  AOI211_X1 g354(.A(new_n529), .B(new_n513), .C1(new_n525), .C2(new_n527), .ZN(new_n541));
  INV_X1    g355(.A(new_n342), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n242), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n520), .A2(new_n543), .A3(new_n522), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n544), .A2(KEYINPUT12), .A3(new_n529), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT12), .B1(new_n544), .B2(new_n529), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n510), .B1(new_n541), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n507), .B1(new_n549), .B2(new_n372), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n525), .A2(new_n527), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n530), .B1(new_n551), .B2(new_n532), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n510), .B1(new_n552), .B2(new_n541), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n530), .A3(new_n532), .ZN(new_n554));
  INV_X1    g368(.A(new_n546), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n544), .A2(KEYINPUT12), .A3(new_n529), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n510), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI211_X1 g373(.A(G469), .B(G902), .C1(new_n553), .C2(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n503), .B(new_n506), .C1(new_n550), .C2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n399), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT78), .ZN(new_n563));
  INV_X1    g377(.A(new_n193), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n564), .A2(new_n504), .A3(new_n497), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT22), .B(G137), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT77), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n565), .B(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n415), .A2(G146), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n413), .A2(KEYINPUT16), .A3(G140), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n417), .B2(KEYINPUT16), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n569), .B1(new_n571), .B2(G146), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT74), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n248), .B2(G128), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n248), .A2(G128), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n240), .A2(KEYINPUT74), .A3(G119), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT24), .B(G110), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(KEYINPUT75), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT23), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(new_n248), .B2(G128), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n240), .A2(KEYINPUT23), .A3(G119), .ZN(new_n582));
  INV_X1    g396(.A(G110), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(new_n575), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT75), .B1(new_n577), .B2(new_n578), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n572), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g401(.A1(new_n577), .A2(new_n578), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n581), .A2(new_n575), .A3(new_n582), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G110), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n588), .B(new_n590), .C1(new_n427), .C2(new_n438), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n568), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(KEYINPUT76), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT76), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n587), .A2(new_n591), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n568), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n593), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n563), .B1(new_n599), .B2(G902), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT25), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(G217), .B1(new_n497), .B2(G902), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT73), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n587), .A2(new_n591), .A3(new_n595), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n595), .B1(new_n587), .B2(new_n591), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n598), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n568), .A2(new_n592), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT78), .B1(new_n609), .B2(new_n372), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n604), .B1(new_n610), .B2(KEYINPUT25), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n599), .B(KEYINPUT79), .ZN(new_n612));
  AOI21_X1  g426(.A(G902), .B1(new_n497), .B2(G217), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n602), .A2(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n322), .A2(new_n562), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT93), .B(G101), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G3));
  INV_X1    g431(.A(new_n398), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n388), .A2(new_n389), .ZN(new_n619));
  INV_X1    g433(.A(new_n373), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n393), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n618), .B1(new_n622), .B2(new_n392), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n485), .A2(G902), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n476), .A2(new_n478), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(KEYINPUT33), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n476), .B2(new_n478), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n624), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT94), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n481), .A2(new_n485), .A3(new_n483), .ZN(new_n632));
  OAI211_X1 g446(.A(KEYINPUT94), .B(new_n624), .C1(new_n626), .C2(new_n628), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n452), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n502), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n623), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n297), .A2(new_n286), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n285), .A2(G902), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n639), .B(new_n614), .C1(new_n640), .C2(new_n300), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n506), .B1(new_n550), .B2(new_n560), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n390), .A2(new_n391), .ZN(new_n648));
  AOI211_X1 g462(.A(new_n393), .B(new_n373), .C1(new_n388), .C2(new_n389), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n398), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n446), .ZN(new_n651));
  INV_X1    g465(.A(new_n447), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT95), .ZN(new_n653));
  INV_X1    g467(.A(new_n451), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT95), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n654), .A2(G475), .B1(new_n447), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n502), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n653), .A2(new_n656), .A3(new_n657), .A4(new_n494), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n647), .B1(new_n650), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n658), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n623), .A2(new_n660), .A3(KEYINPUT96), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n643), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT35), .B(G107), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  OAI21_X1  g479(.A(new_n639), .B1(new_n640), .B2(new_n300), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n611), .A2(new_n602), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n598), .A2(KEYINPUT36), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(new_n597), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n613), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n562), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  NOR2_X1   g490(.A1(new_n507), .A2(new_n372), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n554), .A2(new_n557), .ZN(new_n678));
  AOI22_X1  g492(.A1(new_n678), .A2(new_n510), .B1(new_n531), .B2(new_n539), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n677), .B1(new_n679), .B2(G469), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n553), .A2(new_n559), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n507), .A3(new_n372), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n505), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n499), .B1(new_n500), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  AND4_X1   g500(.A1(new_n494), .A2(new_n653), .A3(new_n656), .A4(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n683), .A2(new_n623), .A3(new_n671), .A4(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n318), .B2(new_n321), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n240), .ZN(G30));
  NAND3_X1  g504(.A1(new_n452), .A2(new_n494), .A3(new_n398), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n685), .B(KEYINPUT39), .Z(new_n692));
  NAND2_X1  g506(.A1(new_n683), .A2(new_n692), .ZN(new_n693));
  AOI211_X1 g507(.A(new_n671), .B(new_n691), .C1(new_n693), .C2(KEYINPUT40), .ZN(new_n694));
  INV_X1    g508(.A(new_n273), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n277), .A2(new_n312), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n696), .A2(KEYINPUT97), .A3(new_n203), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT97), .B1(new_n696), .B2(new_n203), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(G472), .B1(new_n699), .B2(G902), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n288), .A3(new_n298), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT98), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n397), .B(KEYINPUT38), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n694), .A2(new_n702), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT99), .B(G143), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G45));
  AND3_X1   g521(.A1(new_n634), .A2(new_n452), .A3(new_n686), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n683), .A2(new_n623), .A3(new_n671), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n322), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT100), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT100), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n322), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  AOI21_X1  g529(.A(new_n507), .B1(new_n681), .B2(new_n372), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n716), .A2(new_n560), .A3(new_n505), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n322), .A2(new_n614), .A3(new_n638), .A4(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT41), .B(G113), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT101), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n718), .B(new_n720), .ZN(G15));
  NAND4_X1  g535(.A1(new_n322), .A2(new_n662), .A3(new_n614), .A4(new_n717), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  INV_X1    g537(.A(new_n503), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n558), .B1(new_n539), .B2(new_n554), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n541), .A2(new_n547), .A3(new_n510), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n372), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(G469), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n506), .A3(new_n682), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT102), .B1(new_n729), .B2(new_n650), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n716), .A2(new_n560), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT102), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n623), .A2(new_n731), .A3(new_n732), .A4(new_n506), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n724), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n672), .B1(new_n318), .B2(new_n321), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT103), .B(G119), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G21));
  XNOR2_X1  g552(.A(KEYINPUT104), .B(G472), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n285), .B2(G902), .ZN(new_n740));
  OAI22_X1  g554(.A1(new_n290), .A2(new_n296), .B1(new_n314), .B2(new_n303), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n286), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n740), .A2(new_n614), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n691), .B1(new_n392), .B2(new_n622), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n743), .A2(new_n717), .A3(new_n657), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT105), .ZN(new_n746));
  INV_X1    g560(.A(new_n691), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n747), .B(new_n657), .C1(new_n649), .C2(new_n648), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n749), .A2(new_n743), .A3(new_n750), .A4(new_n717), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  NAND4_X1  g567(.A1(new_n708), .A2(new_n740), .A3(new_n671), .A4(new_n742), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n754), .B1(new_n730), .B2(new_n733), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n413), .ZN(G27));
  INV_X1    g570(.A(KEYINPUT106), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n391), .B1(new_n621), .B2(new_n395), .ZN(new_n758));
  INV_X1    g572(.A(new_n396), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n618), .B1(new_n390), .B2(new_n391), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n683), .A2(new_n760), .A3(new_n614), .A4(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n318), .B2(new_n321), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT42), .B1(new_n763), .B2(new_n708), .ZN(new_n764));
  INV_X1    g578(.A(new_n762), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT32), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n639), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n320), .A2(new_n298), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT42), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n635), .A2(new_n769), .A3(new_n685), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n765), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n757), .B1(new_n764), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n322), .A2(new_n765), .A3(new_n708), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n769), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(KEYINPUT106), .A3(new_n771), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(KEYINPUT107), .B(G131), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(G33));
  NAND3_X1  g593(.A1(new_n322), .A2(new_n765), .A3(new_n687), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  OAI21_X1  g595(.A(G469), .B1(new_n679), .B2(KEYINPUT45), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n540), .A2(KEYINPUT45), .A3(new_n548), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n677), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n785), .A2(KEYINPUT46), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n682), .B1(new_n785), .B2(KEYINPUT46), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n506), .B(new_n692), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n452), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n789), .A2(new_n634), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT43), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n666), .A3(new_n671), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n761), .B1(new_n394), .B2(new_n396), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n788), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  XOR2_X1   g611(.A(KEYINPUT108), .B(G137), .Z(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(G39));
  OAI21_X1  g613(.A(new_n506), .B1(new_n786), .B2(new_n787), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n800), .B(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n322), .ZN(new_n803));
  INV_X1    g617(.A(new_n614), .ZN(new_n804));
  INV_X1    g618(.A(new_n796), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n803), .A2(new_n804), .A3(new_n708), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT109), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n802), .A2(KEYINPUT109), .A3(new_n806), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  NAND3_X1  g626(.A1(new_n790), .A2(new_n398), .A3(new_n506), .ZN(new_n813));
  INV_X1    g627(.A(new_n731), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n804), .B(new_n813), .C1(KEYINPUT49), .C2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT110), .ZN(new_n816));
  INV_X1    g630(.A(new_n702), .ZN(new_n817));
  INV_X1    g631(.A(new_n704), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n814), .A2(KEYINPUT49), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n322), .A2(new_n712), .A3(new_n709), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n712), .B1(new_n322), .B2(new_n709), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n730), .A2(new_n733), .ZN(new_n824));
  INV_X1    g638(.A(new_n754), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n642), .A2(new_n650), .A3(new_n672), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n322), .A2(new_n687), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n671), .A2(new_n685), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n701), .A2(new_n744), .A3(new_n683), .A4(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n826), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n823), .A2(new_n831), .A3(KEYINPUT52), .ZN(new_n832));
  OR3_X1    g646(.A1(new_n689), .A2(new_n755), .A3(KEYINPUT113), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT113), .B1(new_n689), .B2(new_n755), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n714), .A3(new_n830), .A4(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n832), .B1(new_n835), .B2(KEYINPUT52), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n683), .A2(new_n760), .A3(new_n761), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT112), .B1(new_n837), .B2(new_n754), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT112), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n825), .A2(new_n839), .A3(new_n683), .A4(new_n805), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n494), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n653), .A3(new_n656), .A4(new_n686), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n642), .A2(new_n796), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n322), .A2(new_n671), .A3(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n841), .A2(new_n780), .A3(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n397), .A2(new_n398), .A3(new_n636), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n562), .A2(new_n673), .B1(new_n847), .B2(new_n643), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n842), .A2(new_n452), .A3(new_n502), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n397), .A2(new_n398), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT111), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT111), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n397), .A2(new_n852), .A3(new_n398), .A4(new_n849), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(new_n643), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n848), .A2(new_n615), .A3(new_n854), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n804), .B(new_n729), .C1(new_n318), .C2(new_n321), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n856), .A2(new_n638), .B1(new_n746), .B2(new_n751), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n856), .A2(new_n662), .B1(new_n735), .B2(new_n734), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n846), .A2(new_n855), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n777), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n836), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT52), .B1(new_n823), .B2(new_n831), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT114), .ZN(new_n864));
  INV_X1    g678(.A(new_n830), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n689), .A2(new_n755), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n714), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n863), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n864), .B1(new_n863), .B2(new_n868), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n841), .A2(new_n780), .A3(new_n845), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n848), .A2(new_n615), .A3(new_n854), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n718), .A2(new_n752), .A3(new_n736), .A4(new_n722), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n873), .A2(new_n874), .A3(new_n773), .A4(new_n776), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n869), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n862), .B1(new_n876), .B2(new_n861), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n729), .A2(new_n796), .A3(new_n498), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n817), .A2(new_n614), .A3(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n881), .A2(new_n452), .A3(new_n634), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT116), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n791), .A2(new_n880), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n740), .A2(new_n671), .A3(new_n742), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n791), .A2(new_n499), .A3(new_n743), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n888), .A2(new_n618), .A3(new_n818), .A4(new_n717), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT50), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n886), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n883), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n731), .A2(new_n505), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT115), .Z(new_n896));
  OAI211_X1 g710(.A(new_n805), .B(new_n888), .C1(new_n802), .C2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT51), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n888), .A2(new_n824), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n899), .B(new_n496), .C1(new_n881), .C2(new_n635), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n900), .A2(KEYINPUT117), .ZN(new_n901));
  INV_X1    g715(.A(new_n768), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n884), .A2(new_n804), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT48), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n900), .B2(KEYINPUT117), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n883), .A2(new_n893), .A3(KEYINPUT51), .ZN(new_n906));
  INV_X1    g720(.A(new_n802), .ZN(new_n907));
  AOI211_X1 g721(.A(new_n796), .B(new_n887), .C1(new_n907), .C2(new_n895), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n901), .B(new_n905), .C1(new_n906), .C2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n898), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n867), .B1(new_n714), .B2(new_n866), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT114), .B1(new_n832), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n863), .A2(new_n864), .A3(new_n868), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n860), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n861), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT53), .B1(new_n764), .B2(new_n772), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n859), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n836), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n915), .A2(new_n878), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n879), .A2(new_n910), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT118), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n495), .A2(new_n189), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n923), .B1(new_n920), .B2(new_n921), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n820), .B1(new_n922), .B2(new_n924), .ZN(G75));
  NAND2_X1  g739(.A1(new_n915), .A2(new_n918), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(G210), .A3(G902), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n381), .A2(new_n385), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(new_n383), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT55), .ZN(new_n930));
  XOR2_X1   g744(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n931));
  AND3_X1   g745(.A1(new_n927), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT56), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n930), .B1(new_n927), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n193), .A2(G952), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT120), .Z(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n932), .A2(new_n934), .A3(new_n937), .ZN(G51));
  INV_X1    g752(.A(KEYINPUT121), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n926), .A2(G902), .A3(new_n784), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n677), .B(KEYINPUT57), .ZN(new_n941));
  AOI221_X4 g755(.A(KEYINPUT54), .B1(new_n836), .B2(new_n917), .C1(new_n914), .C2(new_n861), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n878), .B1(new_n915), .B2(new_n918), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n940), .B1(new_n944), .B2(new_n681), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n939), .B1(new_n945), .B2(new_n935), .ZN(new_n946));
  INV_X1    g760(.A(new_n935), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n870), .A2(new_n875), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT53), .B1(new_n948), .B2(new_n913), .ZN(new_n949));
  INV_X1    g763(.A(new_n918), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT54), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n919), .ZN(new_n952));
  AOI22_X1  g766(.A1(new_n952), .A2(new_n941), .B1(new_n553), .B2(new_n559), .ZN(new_n953));
  OAI211_X1 g767(.A(KEYINPUT121), .B(new_n947), .C1(new_n953), .C2(new_n940), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n946), .A2(new_n954), .ZN(G54));
  NAND4_X1  g769(.A1(new_n926), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT122), .ZN(new_n957));
  INV_X1    g771(.A(new_n442), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n947), .B1(new_n956), .B2(new_n958), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n957), .B1(new_n956), .B2(new_n958), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(G60));
  NOR2_X1   g776(.A1(new_n626), .A2(new_n628), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT123), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n879), .A2(new_n919), .ZN(new_n965));
  NAND2_X1  g779(.A1(G478), .A2(G902), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT59), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n964), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n952), .A2(new_n964), .A3(new_n967), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n968), .A2(new_n937), .A3(new_n969), .ZN(G63));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT60), .Z(new_n972));
  NAND3_X1  g786(.A1(new_n926), .A2(new_n669), .A3(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n926), .A2(new_n972), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n936), .B(new_n973), .C1(new_n974), .C2(new_n612), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G66));
  OAI21_X1  g791(.A(G953), .B1(new_n501), .B2(new_n326), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n874), .A2(new_n855), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(new_n564), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n928), .B1(G898), .B2(new_n193), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G69));
  AOI21_X1  g796(.A(new_n193), .B1(G227), .B2(G900), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n833), .A2(new_n714), .A3(new_n834), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n768), .A2(new_n614), .A3(new_n744), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n788), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n797), .A2(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n811), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n773), .A2(new_n776), .A3(new_n780), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT126), .Z(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n193), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n294), .A2(new_n271), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(new_n429), .Z(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n193), .A2(G900), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT125), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n993), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n996), .A2(new_n564), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n985), .A2(new_n705), .ZN(new_n1003));
  OR2_X1    g817(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n803), .A2(new_n804), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n789), .A2(new_n494), .ZN(new_n1007));
  AOI211_X1 g821(.A(new_n796), .B(new_n693), .C1(new_n635), .C2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n797), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1004), .A2(new_n811), .A3(new_n1005), .A4(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT124), .ZN(new_n1011));
  OR2_X1    g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1002), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n984), .B1(new_n1000), .B2(new_n1014), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n999), .B(new_n983), .C1(new_n1016), .C2(new_n1002), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1015), .A2(new_n1017), .ZN(G72));
  XNOR2_X1  g832(.A(new_n305), .B(KEYINPUT127), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n303), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1012), .A2(new_n979), .A3(new_n1013), .ZN(new_n1021));
  NAND2_X1  g835(.A1(G472), .A2(G902), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT63), .Z(new_n1023));
  AOI21_X1  g837(.A(new_n1020), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n989), .A2(new_n979), .A3(new_n991), .ZN(new_n1025));
  AOI211_X1 g839(.A(new_n303), .B(new_n1019), .C1(new_n1025), .C2(new_n1023), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n304), .A2(new_n306), .A3(new_n273), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(new_n1023), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n947), .B1(new_n877), .B2(new_n1028), .ZN(new_n1029));
  NOR3_X1   g843(.A1(new_n1024), .A2(new_n1026), .A3(new_n1029), .ZN(G57));
endmodule


