//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202));
  OR2_X1    g001(.A1(G57gat), .A2(G64gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G57gat), .A2(G64gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G71gat), .A2(G78gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n203), .B(new_n204), .C1(new_n206), .C2(KEYINPUT9), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(KEYINPUT96), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G71gat), .A2(G78gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n211), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n213), .B1(new_n207), .B2(new_n208), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n202), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(new_n211), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n208), .A3(new_n207), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(KEYINPUT97), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT21), .ZN(new_n221));
  NAND2_X1  g020(.A1(G231gat), .A2(G233gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI211_X1 g022(.A(G231gat), .B(G233gat), .C1(new_n219), .C2(KEYINPUT21), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G127gat), .B(G155gat), .ZN(new_n226));
  XOR2_X1   g025(.A(new_n226), .B(KEYINPUT20), .Z(new_n227));
  AND2_X1   g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n225), .A2(new_n227), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(G183gat), .B(G211gat), .Z(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n231), .B1(new_n228), .B2(new_n229), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G15gat), .B(G22gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(KEYINPUT92), .ZN(new_n237));
  INV_X1    g036(.A(G1gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT92), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n236), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n238), .A2(KEYINPUT16), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G8gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n239), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n244), .B1(new_n239), .B2(new_n243), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n221), .B2(new_n220), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n249), .B(new_n250), .Z(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n233), .A2(new_n251), .A3(new_n234), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g054(.A1(G232gat), .A2(G233gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(KEYINPUT41), .ZN(new_n257));
  XNOR2_X1  g056(.A(G134gat), .B(G162gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G43gat), .B(G50gat), .Z(new_n261));
  INV_X1    g060(.A(KEYINPUT88), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT15), .ZN(new_n264));
  XNOR2_X1  g063(.A(G43gat), .B(G50gat), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n264), .B1(new_n265), .B2(KEYINPUT88), .ZN(new_n266));
  NAND2_X1  g065(.A1(G29gat), .A2(G36gat), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NOR3_X1   g068(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n267), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n263), .A2(new_n266), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT89), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n263), .A2(new_n266), .A3(KEYINPUT89), .A4(new_n271), .ZN(new_n275));
  OR3_X1    g074(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n269), .B1(new_n276), .B2(KEYINPUT91), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT91), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n270), .A2(new_n278), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n263), .A2(new_n266), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G43gat), .ZN(new_n281));
  OR2_X1    g080(.A1(new_n281), .A2(G50gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT90), .B(G50gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(G43gat), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n284), .A2(new_n264), .B1(G29gat), .B2(G36gat), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n274), .A2(new_n275), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n286), .A2(KEYINPUT17), .ZN(new_n287));
  NAND2_X1  g086(.A1(G85gat), .A2(G92gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(KEYINPUT7), .ZN(new_n289));
  NAND2_X1  g088(.A1(G99gat), .A2(G106gat), .ZN(new_n290));
  INV_X1    g089(.A(G85gat), .ZN(new_n291));
  INV_X1    g090(.A(G92gat), .ZN(new_n292));
  AOI22_X1  g091(.A1(KEYINPUT8), .A2(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(G99gat), .B(G106gat), .Z(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n286), .A2(KEYINPUT17), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(KEYINPUT94), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT94), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n299), .B1(new_n286), .B2(KEYINPUT17), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n287), .B(new_n296), .C1(new_n298), .C2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G190gat), .B(G218gat), .Z(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n286), .ZN(new_n304));
  INV_X1    g103(.A(new_n296), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n304), .A2(new_n305), .B1(KEYINPUT41), .B2(new_n256), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n301), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n303), .B1(new_n301), .B2(new_n306), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n260), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n309), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(new_n259), .A3(new_n307), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G120gat), .B(G148gat), .Z(new_n315));
  XNOR2_X1  g114(.A(G176gat), .B(G204gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT100), .ZN(new_n318));
  INV_X1    g117(.A(G230gat), .ZN(new_n319));
  INV_X1    g118(.A(G233gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n215), .A2(new_n296), .A3(new_n218), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT10), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n294), .A2(KEYINPUT99), .ZN(new_n324));
  INV_X1    g123(.A(new_n295), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n294), .A2(KEYINPUT99), .A3(new_n295), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n326), .B(new_n327), .C1(new_n214), .C2(new_n212), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n322), .A2(new_n323), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n219), .A2(KEYINPUT10), .A3(new_n305), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n321), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n321), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n332), .B1(new_n322), .B2(new_n328), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n318), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT101), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n329), .A2(new_n330), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n332), .ZN(new_n337));
  INV_X1    g136(.A(new_n333), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n317), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT101), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n340), .B(new_n318), .C1(new_n331), .C2(new_n333), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n335), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n255), .A2(new_n314), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G78gat), .B(G106gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(G22gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G228gat), .A2(G233gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(G141gat), .B(G148gat), .Z(new_n350));
  INV_X1    g149(.A(G155gat), .ZN(new_n351));
  INV_X1    g150(.A(G162gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(KEYINPUT2), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n350), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G141gat), .B(G148gat), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n354), .B(new_n353), .C1(new_n358), .C2(KEYINPUT2), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n361));
  XNOR2_X1  g160(.A(G211gat), .B(G218gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G197gat), .B(G204gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT22), .ZN(new_n364));
  INV_X1    g163(.A(G211gat), .ZN(new_n365));
  INV_X1    g164(.A(G218gat), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n362), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n362), .B1(new_n367), .B2(new_n363), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n361), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n360), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n363), .A2(new_n367), .ZN(new_n374));
  INV_X1    g173(.A(new_n362), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n368), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n357), .A2(new_n359), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n377), .B1(new_n379), .B2(new_n361), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n349), .B1(new_n373), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n378), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT82), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n382), .B1(new_n371), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT29), .B1(new_n376), .B2(new_n368), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT82), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n360), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n380), .A2(new_n349), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n381), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT83), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n357), .A2(new_n359), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n378), .B1(new_n385), .B2(KEYINPUT82), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n371), .A2(new_n383), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n380), .A2(new_n349), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT83), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n397), .A3(new_n381), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT31), .B(G50gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n390), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n400), .B1(new_n390), .B2(new_n398), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n347), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n390), .A2(new_n398), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n399), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(new_n401), .A3(new_n346), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(G226gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n410), .A2(new_n320), .ZN(new_n411));
  NAND2_X1  g210(.A1(G183gat), .A2(G190gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n412), .A2(KEYINPUT24), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G183gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G190gat), .ZN(new_n416));
  INV_X1    g215(.A(G190gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G183gat), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT24), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n414), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G169gat), .A2(G176gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT23), .ZN(new_n423));
  INV_X1    g222(.A(G169gat), .ZN(new_n424));
  INV_X1    g223(.A(G176gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT23), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n427), .B(KEYINPUT25), .C1(new_n428), .C2(new_n426), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n421), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT67), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n425), .ZN(new_n432));
  NAND2_X1  g231(.A1(KEYINPUT67), .A2(G176gat), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(KEYINPUT23), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n424), .A2(KEYINPUT66), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT66), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(G169gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n427), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT68), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(KEYINPUT68), .B(new_n427), .C1(new_n434), .C2(new_n438), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT65), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n420), .B1(new_n416), .B2(new_n418), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(new_n413), .ZN(new_n445));
  OAI211_X1 g244(.A(KEYINPUT65), .B(new_n414), .C1(new_n419), .C2(new_n420), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n441), .A2(new_n442), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT25), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n430), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n426), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT26), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n422), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT70), .B(KEYINPUT26), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(KEYINPUT71), .A3(new_n450), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT71), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n456), .B1(new_n453), .B2(new_n426), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n452), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT27), .B(G183gat), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT28), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n459), .A2(KEYINPUT69), .A3(new_n460), .A4(new_n417), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n459), .A2(new_n417), .ZN(new_n462));
  XOR2_X1   g261(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n463));
  OAI211_X1 g262(.A(new_n461), .B(new_n412), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n411), .B1(new_n449), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT76), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g267(.A(KEYINPUT76), .B(new_n411), .C1(new_n449), .C2(new_n465), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n361), .B1(new_n449), .B2(new_n465), .ZN(new_n471));
  INV_X1    g270(.A(new_n411), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n377), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n377), .A3(new_n466), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT77), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT77), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n468), .A2(new_n469), .B1(new_n472), .B2(new_n471), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n478), .B(new_n475), .C1(new_n479), .C2(new_n377), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n477), .A2(KEYINPUT37), .A3(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(KEYINPUT84), .B(KEYINPUT37), .Z(new_n482));
  OAI211_X1 g281(.A(new_n475), .B(new_n482), .C1(new_n479), .C2(new_n377), .ZN(new_n483));
  XNOR2_X1  g282(.A(G8gat), .B(G36gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(G64gat), .B(G92gat), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n484), .B(new_n485), .Z(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n481), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT38), .ZN(new_n490));
  XNOR2_X1  g289(.A(G1gat), .B(G29gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT0), .ZN(new_n492));
  XNOR2_X1  g291(.A(G57gat), .B(G85gat), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n492), .B(new_n493), .Z(new_n494));
  XOR2_X1   g293(.A(G127gat), .B(G134gat), .Z(new_n495));
  XNOR2_X1  g294(.A(G113gat), .B(G120gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n495), .B1(KEYINPUT1), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n495), .A2(KEYINPUT1), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT72), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G113gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(KEYINPUT72), .A3(G120gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n498), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n360), .A2(new_n497), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n507));
  OAI21_X1  g306(.A(new_n506), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G225gat), .A2(G233gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n503), .A2(new_n497), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n379), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n360), .A2(new_n372), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n508), .A2(new_n513), .A3(KEYINPUT5), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n510), .A2(new_n391), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n505), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n517), .B(KEYINPUT81), .C1(new_n516), .C2(new_n507), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n504), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n509), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n503), .A2(new_n497), .B1(new_n359), .B2(new_n357), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n516), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT5), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n494), .B(new_n515), .C1(new_n521), .C2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n494), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n525), .B1(new_n518), .B2(new_n520), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(new_n514), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT6), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n475), .B(new_n486), .C1(new_n479), .C2(new_n377), .ZN(new_n532));
  OAI211_X1 g331(.A(KEYINPUT6), .B(new_n527), .C1(new_n528), .C2(new_n514), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT37), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n473), .A2(new_n466), .ZN(new_n536));
  INV_X1    g335(.A(new_n377), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n470), .A2(new_n473), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n377), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT38), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n534), .B1(new_n488), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n409), .B1(new_n490), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT85), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n532), .B(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n477), .A2(new_n480), .A3(new_n487), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT78), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n477), .A2(KEYINPUT78), .A3(new_n480), .A4(new_n487), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n511), .A2(new_n512), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n522), .B1(new_n508), .B2(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n516), .A2(new_n523), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n553), .B(KEYINPUT39), .C1(new_n522), .C2(new_n554), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n555), .B(new_n494), .C1(KEYINPUT39), .C2(new_n553), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT40), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n557), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n529), .A3(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n543), .B(new_n544), .C1(new_n551), .C2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n551), .A2(new_n560), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n488), .A2(new_n541), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n531), .A2(new_n533), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n532), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT38), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n566), .B1(new_n481), .B2(new_n488), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n408), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT85), .B1(new_n562), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n561), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n447), .A2(new_n448), .ZN(new_n571));
  INV_X1    g370(.A(new_n430), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n465), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n510), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n510), .B1(new_n449), .B2(new_n465), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G227gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n579), .A2(new_n320), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT64), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n581), .A2(KEYINPUT34), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n575), .B(new_n576), .C1(new_n579), .C2(new_n320), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n578), .A2(new_n582), .B1(new_n583), .B2(KEYINPUT34), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G99gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT73), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(G15gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(new_n281), .ZN(new_n589));
  INV_X1    g388(.A(new_n581), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n590), .B1(new_n575), .B2(new_n576), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n589), .B1(new_n591), .B2(KEYINPUT33), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT32), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AOI221_X4 g394(.A(new_n593), .B1(KEYINPUT33), .B2(new_n589), .C1(new_n577), .C2(new_n581), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n585), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n576), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n449), .A2(new_n465), .A3(new_n510), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n581), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT32), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n601), .B(new_n589), .C1(KEYINPUT33), .C2(new_n591), .ZN(new_n602));
  INV_X1    g401(.A(new_n596), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(new_n603), .A3(new_n584), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT75), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n597), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n585), .B(KEYINPUT75), .C1(new_n595), .C2(new_n596), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT74), .B(KEYINPUT36), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n597), .A2(new_n604), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT36), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AOI211_X1 g411(.A(new_n564), .B(new_n546), .C1(new_n549), .C2(new_n550), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n612), .B1(new_n613), .B2(new_n408), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n570), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n606), .A2(new_n607), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n531), .A2(new_n533), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n409), .A2(KEYINPUT35), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n551), .A2(new_n617), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT35), .ZN(new_n621));
  AND4_X1   g420(.A1(new_n408), .A2(new_n597), .A3(new_n604), .A4(new_n618), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n621), .B1(new_n551), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n620), .B1(new_n623), .B2(KEYINPUT86), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT86), .ZN(new_n625));
  AOI211_X1 g424(.A(new_n625), .B(new_n621), .C1(new_n551), .C2(new_n622), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n616), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n629));
  XNOR2_X1  g428(.A(G113gat), .B(G141gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(G169gat), .B(G197gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(KEYINPUT12), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G229gat), .A2(G233gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n637), .B(KEYINPUT13), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n248), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n304), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n248), .A2(new_n286), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n298), .A2(new_n300), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT93), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n645), .B1(new_n246), .B2(new_n247), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n241), .A2(G1gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n242), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n237), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(G8gat), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(KEYINPUT93), .A3(new_n245), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n287), .A2(new_n646), .A3(new_n651), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n637), .B(new_n641), .C1(new_n644), .C2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT18), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n643), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n650), .A2(KEYINPUT93), .A3(new_n245), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT93), .B1(new_n650), .B2(new_n245), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n658), .B(new_n287), .C1(new_n300), .C2(new_n298), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n659), .A2(KEYINPUT18), .A3(new_n637), .A4(new_n641), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n636), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n653), .A2(new_n654), .ZN(new_n663));
  INV_X1    g462(.A(new_n643), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n660), .A2(new_n663), .A3(new_n664), .A4(new_n636), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n628), .A2(new_n629), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n614), .B1(new_n569), .B2(new_n561), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n624), .A2(new_n626), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT95), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n344), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n618), .B(KEYINPUT102), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  INV_X1    g474(.A(new_n551), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT16), .B(G8gat), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n672), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n244), .B1(new_n672), .B2(new_n676), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT42), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT42), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(G1325gat));
  INV_X1    g484(.A(G15gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n672), .A2(new_n686), .A3(new_n617), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n609), .A2(new_n611), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n672), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n689), .B2(new_n686), .ZN(G1326gat));
  NAND2_X1  g489(.A1(new_n672), .A2(new_n409), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  INV_X1    g492(.A(new_n342), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n255), .A2(new_n694), .A3(new_n314), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT103), .Z(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n667), .B2(new_n671), .ZN(new_n697));
  INV_X1    g496(.A(new_n673), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(G29gat), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n700), .A2(KEYINPUT45), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(KEYINPUT45), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n314), .B1(new_n668), .B2(new_n669), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g504(.A(KEYINPUT44), .B(new_n314), .C1(new_n668), .C2(new_n669), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n255), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n655), .A2(new_n660), .A3(new_n636), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n661), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n708), .A2(new_n710), .A3(new_n342), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n707), .A2(new_n673), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G29gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n701), .A2(new_n702), .A3(new_n713), .ZN(G1328gat));
  NOR2_X1   g513(.A1(new_n551), .A2(G36gat), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n697), .A2(new_n715), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n716), .A2(KEYINPUT46), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(KEYINPUT46), .ZN(new_n718));
  INV_X1    g517(.A(G36gat), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n707), .A2(new_n676), .A3(new_n711), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n717), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(G1329gat));
  NOR2_X1   g520(.A1(new_n612), .A2(new_n281), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n711), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(G43gat), .B1(new_n697), .B2(new_n617), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT47), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT47), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n697), .A2(new_n617), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n727), .B(new_n723), .C1(new_n728), .C2(G43gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n729), .ZN(G1330gat));
  NAND4_X1  g529(.A1(new_n705), .A2(new_n409), .A3(new_n706), .A4(new_n711), .ZN(new_n731));
  INV_X1    g530(.A(new_n283), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n696), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n408), .A2(new_n732), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT105), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n629), .B1(new_n628), .B2(new_n666), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n670), .A2(KEYINPUT95), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n734), .B(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT48), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  AOI211_X1 g542(.A(KEYINPUT104), .B(new_n743), .C1(new_n733), .C2(new_n739), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n742), .A2(new_n744), .ZN(G1331gat));
  NOR3_X1   g544(.A1(new_n666), .A2(new_n255), .A3(new_n314), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n342), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT106), .Z(new_n748));
  AND2_X1   g547(.A1(new_n628), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n673), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g550(.A1(new_n749), .A2(KEYINPUT107), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n628), .A2(new_n748), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n551), .B(KEYINPUT108), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n756), .B(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n756), .A2(new_n758), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(new_n759), .ZN(G1333gat));
  NAND4_X1  g562(.A1(new_n752), .A2(new_n755), .A3(G71gat), .A4(new_n688), .ZN(new_n764));
  INV_X1    g563(.A(G71gat), .ZN(new_n765));
  INV_X1    g564(.A(new_n617), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n753), .B2(new_n766), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n764), .A2(KEYINPUT50), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT50), .B1(new_n764), .B2(new_n767), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(G1334gat));
  NAND2_X1  g569(.A1(new_n756), .A2(new_n409), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G78gat), .ZN(new_n772));
  INV_X1    g571(.A(G78gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n756), .A2(new_n773), .A3(new_n409), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(G1335gat));
  NOR2_X1   g574(.A1(new_n708), .A2(new_n666), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n314), .B(new_n776), .C1(new_n668), .C2(new_n669), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n628), .A2(KEYINPUT51), .A3(new_n314), .A4(new_n776), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n777), .A2(new_n779), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n780), .B1(new_n783), .B2(new_n778), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT111), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n786), .B(new_n780), .C1(new_n783), .C2(new_n778), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n698), .A2(new_n694), .A3(G85gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n708), .A2(new_n666), .A3(new_n694), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n705), .A2(new_n673), .A3(new_n706), .A4(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n291), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n792), .B2(new_n791), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n789), .A2(new_n794), .ZN(G1336gat));
  NOR3_X1   g594(.A1(new_n757), .A2(G92gat), .A3(new_n694), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n784), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n705), .A2(new_n706), .A3(new_n758), .A4(new_n790), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G92gat), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n705), .A2(new_n676), .A3(new_n706), .A4(new_n790), .ZN(new_n803));
  AOI22_X1  g602(.A1(G92gat), .A2(new_n803), .B1(new_n783), .B2(new_n796), .ZN(new_n804));
  OAI22_X1  g603(.A1(new_n798), .A2(new_n802), .B1(new_n804), .B2(new_n801), .ZN(G1337gat));
  NOR3_X1   g604(.A1(new_n766), .A2(G99gat), .A3(new_n694), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n785), .A2(new_n787), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n707), .A2(new_n688), .A3(new_n790), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G99gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(G1338gat));
  NOR3_X1   g609(.A1(new_n408), .A2(G106gat), .A3(new_n694), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n784), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n705), .A2(new_n409), .A3(new_n706), .A4(new_n790), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G106gat), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI22_X1  g616(.A1(G106gat), .A2(new_n814), .B1(new_n783), .B2(new_n811), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n813), .A2(new_n817), .B1(new_n818), .B2(new_n816), .ZN(G1339gat));
  NAND2_X1  g618(.A1(new_n746), .A2(new_n694), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n329), .A2(new_n330), .A3(new_n321), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT112), .A4(new_n321), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n823), .A2(new_n337), .A3(KEYINPUT54), .A4(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n317), .B1(new_n331), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(KEYINPUT55), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n339), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT113), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(new_n831), .A3(new_n339), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n825), .A2(new_n827), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n830), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n637), .B1(new_n659), .B2(new_n641), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n641), .A2(new_n642), .A3(new_n639), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n634), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n665), .A2(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n836), .A2(new_n313), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n665), .A2(new_n839), .A3(new_n342), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n665), .A2(new_n839), .A3(KEYINPUT114), .A4(new_n342), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n844), .B(new_n845), .C1(new_n836), .C2(new_n710), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n841), .B1(new_n846), .B2(new_n313), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n820), .B1(new_n847), .B2(new_n708), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n408), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n758), .A2(new_n766), .A3(new_n698), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851), .B2(new_n710), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT115), .ZN(new_n853));
  AND4_X1   g652(.A1(new_n408), .A2(new_n848), .A3(new_n610), .A4(new_n673), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n757), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n666), .A2(new_n501), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(G1340gat));
  NAND3_X1  g656(.A1(new_n849), .A2(new_n342), .A3(new_n850), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n858), .A2(KEYINPUT116), .A3(G120gat), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT116), .B1(new_n858), .B2(G120gat), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n694), .A2(G120gat), .ZN(new_n861));
  OAI22_X1  g660(.A1(new_n859), .A2(new_n860), .B1(new_n855), .B2(new_n861), .ZN(G1341gat));
  OAI21_X1  g661(.A(G127gat), .B1(new_n851), .B2(new_n255), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n255), .A2(G127gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n855), .B2(new_n864), .ZN(G1342gat));
  OAI21_X1  g664(.A(G134gat), .B1(new_n851), .B2(new_n313), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT117), .ZN(new_n867));
  INV_X1    g666(.A(G134gat), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n676), .A2(new_n313), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  XOR2_X1   g669(.A(new_n870), .B(KEYINPUT56), .Z(new_n871));
  NAND2_X1  g670(.A1(new_n867), .A2(new_n871), .ZN(G1343gat));
  AND2_X1   g671(.A1(new_n848), .A2(new_n409), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n688), .A2(new_n698), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n757), .A3(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(G141gat), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n666), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT58), .B1(new_n878), .B2(KEYINPUT119), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n874), .A2(new_n757), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n828), .A2(new_n339), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n835), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n835), .A2(KEYINPUT118), .A3(new_n339), .A4(new_n828), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n666), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n314), .B1(new_n887), .B2(new_n842), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n255), .B1(new_n888), .B2(new_n841), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n408), .B1(new_n889), .B2(new_n820), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n881), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n848), .A2(new_n891), .A3(new_n409), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n876), .B1(new_n894), .B2(new_n666), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n880), .B1(new_n878), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(new_n878), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n879), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1344gat));
  OR3_X1    g698(.A1(new_n875), .A2(G148gat), .A3(new_n694), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G148gat), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n894), .B2(new_n342), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n848), .A2(KEYINPUT57), .A3(new_n409), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n886), .B1(new_n709), .B2(new_n661), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT118), .B1(new_n882), .B2(new_n835), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n842), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n841), .B1(new_n907), .B2(new_n313), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n820), .B1(new_n908), .B2(new_n708), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT57), .B1(new_n909), .B2(new_n409), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n342), .B(new_n881), .C1(new_n904), .C2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n901), .B1(new_n911), .B2(G148gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n900), .B1(new_n903), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT120), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n915), .B(new_n900), .C1(new_n903), .C2(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1345gat));
  INV_X1    g716(.A(new_n894), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n918), .A2(new_n351), .A3(new_n255), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n875), .A2(new_n255), .ZN(new_n920));
  AOI21_X1  g719(.A(G155gat), .B1(new_n920), .B2(KEYINPUT121), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n920), .A2(KEYINPUT121), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(G1346gat));
  OAI21_X1  g722(.A(G162gat), .B1(new_n918), .B2(new_n313), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n873), .A2(new_n352), .A3(new_n869), .A4(new_n874), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n551), .A2(new_n673), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n617), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT122), .Z(new_n929));
  NAND2_X1  g728(.A1(new_n849), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n710), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n848), .A2(new_n698), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n758), .A2(new_n408), .A3(new_n610), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n666), .A2(new_n435), .A3(new_n437), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(G1348gat));
  INV_X1    g736(.A(new_n935), .ZN(new_n938));
  AOI21_X1  g737(.A(G176gat), .B1(new_n938), .B2(new_n342), .ZN(new_n939));
  INV_X1    g738(.A(new_n930), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n694), .B1(new_n432), .B2(new_n433), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(G1349gat));
  OAI21_X1  g741(.A(G183gat), .B1(new_n930), .B2(new_n255), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n933), .A2(new_n459), .A3(new_n708), .A4(new_n934), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g748(.A1(new_n938), .A2(new_n417), .A3(new_n314), .ZN(new_n950));
  OAI21_X1  g749(.A(G190gat), .B1(new_n930), .B2(new_n313), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n951), .A2(KEYINPUT61), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(KEYINPUT61), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n950), .B1(new_n952), .B2(new_n953), .ZN(G1351gat));
  NAND2_X1  g753(.A1(new_n927), .A2(new_n612), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n956), .B1(new_n904), .B2(new_n910), .ZN(new_n957));
  OAI21_X1  g756(.A(G197gat), .B1(new_n957), .B2(new_n710), .ZN(new_n958));
  NOR4_X1   g757(.A1(new_n932), .A2(new_n408), .A3(new_n688), .A4(new_n757), .ZN(new_n959));
  INV_X1    g758(.A(G197gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n960), .A3(new_n666), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT124), .ZN(G1352gat));
  NOR2_X1   g762(.A1(new_n694), .A2(G204gat), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n965));
  AOI22_X1  g764(.A1(new_n959), .A2(new_n964), .B1(KEYINPUT125), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n965), .A2(KEYINPUT125), .ZN(new_n967));
  XOR2_X1   g766(.A(new_n966), .B(new_n967), .Z(new_n968));
  OAI21_X1  g767(.A(G204gat), .B1(new_n957), .B2(new_n694), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(G1353gat));
  NAND3_X1  g769(.A1(new_n959), .A2(new_n365), .A3(new_n708), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n708), .B(new_n956), .C1(new_n904), .C2(new_n910), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT63), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n365), .B1(KEYINPUT126), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n973), .A2(KEYINPUT126), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n972), .B2(new_n974), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n971), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI211_X1 g779(.A(KEYINPUT127), .B(new_n971), .C1(new_n976), .C2(new_n977), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1354gat));
  OAI21_X1  g781(.A(G218gat), .B1(new_n957), .B2(new_n313), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n959), .A2(new_n366), .A3(new_n314), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1355gat));
endmodule


