//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n523, new_n524, new_n525, new_n526, new_n527, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n539, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n591, new_n594, new_n596, new_n597, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1113, new_n1114;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n452), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n463), .A2(new_n465), .A3(G137), .A4(new_n461), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n462), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n463), .A2(new_n465), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n461), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  NAND4_X1  g057(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n461), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT68), .ZN(new_n484));
  XNOR2_X1  g059(.A(KEYINPUT3), .B(G2104), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n485), .A2(new_n486), .A3(G138), .A4(new_n461), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n484), .A2(new_n487), .A3(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n483), .A2(KEYINPUT68), .A3(new_n489), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n463), .A2(new_n465), .A3(G126), .A4(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n488), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G543), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n505), .A2(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  INV_X1    g088(.A(new_n507), .ZN(new_n514));
  AND2_X1   g089(.A1(G63), .A2(G651), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n514), .A2(G89), .B1(new_n502), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n509), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G51), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n516), .A2(new_n518), .A3(new_n520), .ZN(G286));
  INV_X1    g096(.A(G286), .ZN(G168));
  AOI22_X1  g097(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n504), .ZN(new_n524));
  INV_X1    g099(.A(G90), .ZN(new_n525));
  INV_X1    g100(.A(G52), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n507), .A2(new_n525), .B1(new_n509), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n524), .A2(new_n527), .ZN(G301));
  INV_X1    g103(.A(G301), .ZN(G171));
  AOI22_X1  g104(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n504), .ZN(new_n531));
  INV_X1    g106(.A(G81), .ZN(new_n532));
  INV_X1    g107(.A(G43), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n507), .A2(new_n532), .B1(new_n509), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT69), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(KEYINPUT69), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n531), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  AND3_X1   g113(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G36), .ZN(G176));
  XOR2_X1   g115(.A(KEYINPUT70), .B(KEYINPUT8), .Z(new_n541));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n539), .A2(new_n543), .ZN(G188));
  NAND3_X1  g119(.A1(new_n506), .A2(G53), .A3(G543), .ZN(new_n545));
  XOR2_X1   g120(.A(new_n545), .B(KEYINPUT9), .Z(new_n546));
  AOI22_X1  g121(.A1(new_n502), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G91), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n547), .A2(new_n504), .B1(new_n507), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(G299));
  NAND2_X1  g126(.A1(new_n514), .A2(G87), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n517), .A2(G49), .ZN(new_n553));
  OAI21_X1  g128(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(G288));
  NAND2_X1  g130(.A1(G73), .A2(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n499), .A2(new_n501), .ZN(new_n557));
  INV_X1    g132(.A(G61), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G651), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT71), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n559), .A2(new_n562), .A3(G651), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n561), .A2(new_n563), .B1(G48), .B2(new_n517), .ZN(new_n564));
  INV_X1    g139(.A(G86), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n565), .B2(new_n507), .ZN(G305));
  AOI22_X1  g141(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(new_n504), .ZN(new_n568));
  INV_X1    g143(.A(G85), .ZN(new_n569));
  INV_X1    g144(.A(G47), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n507), .A2(new_n569), .B1(new_n509), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G290));
  NAND2_X1  g148(.A1(G301), .A2(G868), .ZN(new_n574));
  INV_X1    g149(.A(G66), .ZN(new_n575));
  INV_X1    g150(.A(G79), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n557), .A2(new_n575), .B1(new_n576), .B2(new_n498), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI221_X1 g154(.A(KEYINPUT72), .B1(new_n576), .B2(new_n498), .C1(new_n557), .C2(new_n575), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n579), .A2(G651), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n517), .A2(G54), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT10), .B1(new_n514), .B2(G92), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT10), .ZN(new_n584));
  INV_X1    g159(.A(G92), .ZN(new_n585));
  NOR3_X1   g160(.A1(new_n507), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n581), .B(new_n582), .C1(new_n583), .C2(new_n586), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT73), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n574), .B1(new_n588), .B2(G868), .ZN(G284));
  OAI21_X1  g164(.A(new_n574), .B1(new_n588), .B2(G868), .ZN(G321));
  NAND2_X1  g165(.A1(G286), .A2(G868), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n591), .B1(G868), .B2(new_n550), .ZN(G297));
  OAI21_X1  g167(.A(new_n591), .B1(G868), .B2(new_n550), .ZN(G280));
  XNOR2_X1  g168(.A(KEYINPUT74), .B(G559), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n588), .B1(G860), .B2(new_n594), .ZN(G148));
  NAND2_X1  g170(.A1(new_n588), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G868), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(G868), .B2(new_n537), .ZN(G323));
  XOR2_X1   g173(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n599));
  XNOR2_X1  g174(.A(G323), .B(new_n599), .ZN(G282));
  NAND2_X1  g175(.A1(new_n477), .A2(G135), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n475), .A2(G123), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n461), .A2(G111), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT78), .Z(new_n604));
  OAI21_X1  g179(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n601), .B(new_n602), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  OAI22_X1  g181(.A1(new_n606), .A2(G2096), .B1(KEYINPUT77), .B2(G2100), .ZN(new_n607));
  NAND2_X1  g182(.A1(KEYINPUT77), .A2(G2100), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT76), .Z(new_n610));
  NAND2_X1  g185(.A1(new_n485), .A2(new_n470), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n610), .B(new_n612), .ZN(new_n613));
  AOI211_X1 g188(.A(new_n607), .B(new_n613), .C1(G2096), .C2(new_n606), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT79), .ZN(G156));
  XNOR2_X1  g190(.A(KEYINPUT15), .B(G2435), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT81), .B(G2438), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(G2427), .B(G2430), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT14), .ZN(new_n621));
  XOR2_X1   g196(.A(G2443), .B(G2446), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(G2451), .B(G2454), .Z(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n623), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G1341), .B(G1348), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G14), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT82), .ZN(G401));
  XOR2_X1   g206(.A(G2072), .B(G2078), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT83), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT17), .Z(new_n634));
  XOR2_X1   g209(.A(G2067), .B(G2678), .Z(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT84), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2084), .B(G2090), .ZN(new_n638));
  INV_X1    g213(.A(new_n633), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n637), .B(new_n638), .C1(new_n639), .C2(new_n636), .ZN(new_n640));
  OR3_X1    g215(.A1(new_n634), .A2(new_n638), .A3(new_n636), .ZN(new_n641));
  NOR3_X1   g216(.A1(new_n633), .A2(new_n638), .A3(new_n635), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT18), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2096), .B(G2100), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(G227));
  XNOR2_X1  g221(.A(G1971), .B(G1976), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n647), .B(new_n648), .Z(new_n649));
  XOR2_X1   g224(.A(G1956), .B(G2474), .Z(new_n650));
  XOR2_X1   g225(.A(G1961), .B(G1966), .Z(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT86), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n650), .A2(new_n651), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT20), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n653), .A2(new_n656), .ZN(new_n659));
  AOI211_X1 g234(.A(new_n655), .B(new_n658), .C1(new_n649), .C2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n661));
  INV_X1    g236(.A(G1986), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1991), .B(G1996), .ZN(new_n665));
  INV_X1    g240(.A(G1981), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT87), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n664), .B(new_n668), .ZN(G229));
  MUX2_X1   g244(.A(G6), .B(G305), .S(G16), .Z(new_n670));
  OR2_X1    g245(.A1(new_n670), .A2(KEYINPUT91), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(KEYINPUT91), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT32), .B(G1981), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(G16), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G22), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(G166), .B2(new_n677), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G1971), .ZN(new_n680));
  NOR2_X1   g255(.A1(G16), .A2(G23), .ZN(new_n681));
  INV_X1    g256(.A(G288), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(G16), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT33), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n671), .A2(new_n674), .A3(new_n672), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n676), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n689));
  NOR2_X1   g264(.A1(G25), .A2(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n477), .A2(G131), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT88), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n475), .A2(G119), .ZN(new_n693));
  OAI21_X1  g268(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n461), .A2(G107), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT89), .Z(new_n698));
  AOI21_X1  g273(.A(new_n690), .B1(new_n698), .B2(G29), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT35), .B(G1991), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n699), .B(new_n700), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n677), .A2(G24), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n572), .B2(new_n677), .ZN(new_n703));
  MUX2_X1   g278(.A(new_n702), .B(new_n703), .S(KEYINPUT90), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(new_n662), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT34), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n676), .A2(new_n706), .A3(new_n686), .A4(new_n687), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n689), .A2(new_n701), .A3(new_n705), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT36), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n677), .A2(G5), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G171), .B2(new_n677), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT103), .ZN(new_n712));
  INV_X1    g287(.A(G1961), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT95), .B(KEYINPUT24), .Z(new_n715));
  INV_X1    g290(.A(G34), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n717), .A2(new_n718), .A3(G29), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT96), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(G160), .A2(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(new_n720), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT97), .Z(new_n725));
  INV_X1    g300(.A(G2084), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OR2_X1    g302(.A1(G29), .A2(G32), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n475), .A2(G129), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT98), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n477), .A2(G141), .B1(G105), .B2(new_n470), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT99), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT26), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G29), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n728), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT27), .B(G1996), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT100), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n714), .A2(new_n727), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT104), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n677), .A2(G4), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n588), .B2(new_n677), .ZN(new_n747));
  INV_X1    g322(.A(G1348), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n737), .A2(G26), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n475), .A2(G128), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n477), .A2(G140), .ZN(new_n754));
  OR2_X1    g329(.A1(G104), .A2(G2105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n755), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n752), .B1(new_n758), .B2(new_n737), .ZN(new_n759));
  INV_X1    g334(.A(G2067), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(G29), .A2(G33), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n470), .A2(G103), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT93), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT25), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n477), .A2(G139), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n485), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n765), .B(new_n766), .C1(new_n461), .C2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(new_n737), .ZN(new_n769));
  INV_X1    g344(.A(G2072), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT30), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G28), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT102), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n774), .B(new_n737), .C1(new_n772), .C2(G28), .ZN(new_n775));
  AND4_X1   g350(.A1(new_n749), .A2(new_n761), .A3(new_n771), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n738), .A2(new_n741), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n769), .A2(new_n770), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT94), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n745), .A2(new_n776), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  OAI22_X1  g355(.A1(new_n712), .A2(new_n713), .B1(new_n725), .B2(new_n726), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n737), .A2(G35), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G162), .B2(new_n737), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT29), .Z(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(G2090), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n677), .A2(G19), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n537), .B2(new_n677), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n787), .A2(KEYINPUT106), .B1(G1341), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G1341), .B2(new_n789), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n787), .A2(KEYINPUT106), .ZN(new_n792));
  NOR4_X1   g367(.A1(new_n780), .A2(new_n781), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(G168), .A2(G16), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G16), .B2(G21), .ZN(new_n795));
  INV_X1    g370(.A(G1966), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT101), .ZN(new_n798));
  INV_X1    g373(.A(G11), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(KEYINPUT31), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(KEYINPUT31), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n606), .B2(new_n737), .ZN(new_n802));
  AOI211_X1 g377(.A(new_n800), .B(new_n802), .C1(new_n785), .C2(G2090), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n709), .A2(new_n793), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n795), .A2(new_n796), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n677), .A2(KEYINPUT23), .A3(G20), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT23), .ZN(new_n808));
  INV_X1    g383(.A(G20), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(G16), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n807), .B(new_n810), .C1(new_n550), .C2(new_n677), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1956), .ZN(new_n812));
  NOR2_X1   g387(.A1(G27), .A2(G29), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G164), .B2(G29), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT105), .B(G2078), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NOR4_X1   g392(.A1(new_n804), .A2(new_n806), .A3(new_n812), .A4(new_n817), .ZN(G311));
  NOR2_X1   g393(.A1(new_n804), .A2(new_n817), .ZN(new_n819));
  INV_X1    g394(.A(new_n812), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n819), .A2(new_n805), .A3(new_n820), .ZN(G150));
  AOI22_X1  g396(.A1(new_n514), .A2(G93), .B1(G55), .B2(new_n517), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(new_n504), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G860), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n588), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT39), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n537), .B(new_n826), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n830), .B(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n828), .B1(new_n834), .B2(G860), .ZN(G145));
  XNOR2_X1  g410(.A(new_n736), .B(new_n768), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n758), .B(new_n496), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT109), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n697), .B(new_n612), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n477), .A2(G142), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n475), .A2(G130), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n461), .A2(G118), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT108), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n841), .B(new_n842), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n840), .B(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n838), .A2(new_n839), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n481), .B(G160), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(new_n606), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n838), .B(new_n847), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n848), .B(new_n850), .C1(new_n851), .C2(new_n839), .ZN(new_n852));
  INV_X1    g427(.A(G37), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n852), .B(new_n853), .C1(new_n851), .C2(new_n850), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g430(.A(G868), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n826), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n596), .B(new_n831), .Z(new_n858));
  XOR2_X1   g433(.A(new_n550), .B(new_n587), .Z(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT110), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n859), .B(KEYINPUT41), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT42), .Z(new_n864));
  XNOR2_X1  g439(.A(G305), .B(G288), .ZN(new_n865));
  XNOR2_X1  g440(.A(G290), .B(G303), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n864), .B(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n857), .B1(new_n868), .B2(new_n856), .ZN(G295));
  OAI21_X1  g444(.A(new_n857), .B1(new_n868), .B2(new_n856), .ZN(G331));
  XOR2_X1   g445(.A(G286), .B(G301), .Z(new_n871));
  AOI21_X1  g446(.A(KEYINPUT111), .B1(new_n831), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n831), .B(new_n871), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n872), .B1(new_n873), .B2(KEYINPUT111), .ZN(new_n874));
  INV_X1    g449(.A(new_n859), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n874), .A2(new_n875), .B1(new_n862), .B2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n853), .B1(new_n876), .B2(new_n867), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(KEYINPUT112), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n867), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT112), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n880), .B(new_n853), .C1(new_n876), .C2(new_n867), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n878), .A2(KEYINPUT43), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(new_n853), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n873), .A2(KEYINPUT111), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n862), .B1(new_n885), .B2(new_n872), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n860), .A2(new_n873), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n867), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n883), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n884), .A2(new_n888), .A3(new_n883), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n893), .B1(new_n883), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n892), .B1(new_n895), .B2(new_n891), .ZN(G397));
  INV_X1    g471(.A(KEYINPUT122), .ZN(new_n897));
  NAND2_X1  g472(.A1(G303), .A2(G8), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(G1971), .ZN(new_n901));
  INV_X1    g476(.A(G40), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n468), .A2(new_n472), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n483), .A2(KEYINPUT68), .A3(new_n489), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n905), .A2(new_n494), .ZN(new_n906));
  AOI21_X1  g481(.A(G1384), .B1(new_n906), .B2(new_n488), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n904), .B1(new_n907), .B2(KEYINPUT45), .ZN(new_n908));
  INV_X1    g483(.A(G1384), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n484), .A2(new_n487), .A3(KEYINPUT4), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n490), .A2(new_n493), .A3(new_n492), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT45), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT115), .B1(new_n908), .B2(new_n914), .ZN(new_n915));
  OAI211_X1 g490(.A(KEYINPUT45), .B(new_n909), .C1(new_n910), .C2(new_n911), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n903), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT115), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT45), .B1(new_n496), .B2(new_n909), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n901), .B1(new_n915), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT116), .ZN(new_n922));
  XNOR2_X1  g497(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n909), .B(new_n924), .C1(new_n910), .C2(new_n911), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT50), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n925), .B(new_n903), .C1(new_n907), .C2(new_n926), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n927), .A2(G2090), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n918), .B1(new_n917), .B2(new_n919), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n914), .A2(KEYINPUT115), .A3(new_n903), .A4(new_n916), .ZN(new_n930));
  AOI21_X1  g505(.A(G1971), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT116), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n922), .A2(new_n928), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n900), .B1(new_n934), .B2(G8), .ZN(new_n935));
  INV_X1    g510(.A(G8), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n907), .B2(new_n903), .ZN(new_n937));
  INV_X1    g512(.A(G1976), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n937), .B(KEYINPUT118), .C1(new_n938), .C2(G288), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(new_n938), .A3(G288), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT52), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(new_n942), .A3(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(KEYINPUT119), .B(G86), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n564), .B1(new_n507), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(G1981), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n564), .B(new_n666), .C1(new_n565), .C2(new_n507), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT49), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n949), .A2(KEYINPUT49), .A3(new_n950), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n937), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n946), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n897), .B1(new_n935), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n956), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n929), .A2(new_n930), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n932), .B1(new_n959), .B2(new_n901), .ZN(new_n960));
  AOI211_X1 g535(.A(KEYINPUT116), .B(G1971), .C1(new_n929), .C2(new_n930), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n936), .B1(new_n962), .B2(new_n928), .ZN(new_n963));
  OAI211_X1 g538(.A(KEYINPUT122), .B(new_n958), .C1(new_n963), .C2(new_n900), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n934), .A2(G8), .A3(new_n900), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n904), .B1(new_n912), .B2(KEYINPUT50), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(new_n726), .A3(new_n925), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n796), .B1(new_n917), .B2(new_n919), .ZN(new_n968));
  AOI211_X1 g543(.A(new_n936), .B(G286), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n957), .A2(new_n964), .A3(new_n965), .A4(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT63), .ZN(new_n971));
  INV_X1    g546(.A(G2078), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n929), .A2(new_n972), .A3(new_n930), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n974));
  AOI22_X1  g549(.A1(new_n973), .A2(new_n974), .B1(new_n713), .B2(new_n927), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n908), .A2(KEYINPUT53), .A3(new_n972), .A4(new_n914), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(G301), .B(KEYINPUT54), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n967), .A2(new_n968), .A3(G168), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(G8), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT51), .ZN(new_n981));
  AOI21_X1  g556(.A(G168), .B1(new_n967), .B2(new_n968), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n983));
  OAI211_X1 g558(.A(G8), .B(new_n979), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n977), .A2(new_n978), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n903), .B1(new_n912), .B2(KEYINPUT50), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n907), .A2(new_n924), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n986), .A2(new_n987), .A3(G2090), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n931), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(G8), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n899), .ZN(new_n991));
  AND4_X1   g566(.A1(new_n965), .A2(new_n985), .A3(new_n958), .A4(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n912), .B(KEYINPUT113), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n993), .A2(KEYINPUT45), .ZN(new_n994));
  OR4_X1    g569(.A1(new_n974), .A2(new_n994), .A3(G2078), .A4(new_n917), .ZN(new_n995));
  INV_X1    g570(.A(new_n978), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(new_n975), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n927), .A2(new_n748), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT123), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n907), .A2(new_n999), .A3(new_n903), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n496), .A2(new_n909), .A3(new_n903), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT123), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n1002), .A3(new_n760), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n588), .B1(new_n1004), .B2(KEYINPUT60), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT73), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n587), .B(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n1003), .B2(new_n998), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT125), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1004), .A2(new_n588), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT125), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT60), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n998), .B2(new_n1003), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1010), .B(new_n1011), .C1(new_n588), .C2(new_n1013), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1009), .A2(KEYINPUT60), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT60), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT124), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n904), .B1(new_n907), .B2(new_n926), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n912), .A2(new_n923), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1956), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT56), .B(G2072), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n917), .A2(new_n919), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1017), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n550), .A2(KEYINPUT57), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n546), .B2(new_n549), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1956), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n986), .B2(new_n987), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n908), .A2(new_n914), .A3(new_n1021), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n1032), .A3(KEYINPUT124), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1024), .A2(new_n1029), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT61), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(new_n1028), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1029), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1028), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1035), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT58), .B(G1341), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1042), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n917), .A2(G1996), .A3(new_n919), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n537), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT59), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1047), .B(new_n537), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1038), .A2(new_n1041), .A3(new_n1049), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1015), .A2(new_n1016), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1034), .B1(new_n1010), .B2(new_n1039), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n992), .B(new_n997), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n900), .B1(new_n989), .B2(G8), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n963), .B2(new_n900), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1055), .A2(KEYINPUT121), .A3(new_n958), .A4(new_n969), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT63), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n965), .A2(new_n991), .A3(new_n958), .A4(new_n969), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1056), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n955), .A2(new_n938), .A3(new_n682), .ZN(new_n1062));
  XOR2_X1   g637(.A(new_n950), .B(KEYINPUT120), .Z(new_n1063));
  AND2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1001), .A2(G8), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1064), .A2(new_n1065), .B1(new_n965), .B2(new_n956), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n965), .A2(new_n958), .A3(new_n991), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n981), .A2(new_n984), .ZN(new_n1068));
  OAI211_X1 g643(.A(G171), .B(new_n977), .C1(new_n1068), .C2(KEYINPUT62), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1068), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT126), .B1(new_n1068), .B2(KEYINPUT62), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1066), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n971), .A2(new_n1053), .A3(new_n1061), .A4(new_n1074), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n993), .A2(KEYINPUT45), .A3(new_n904), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(G1996), .A3(new_n736), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(KEYINPUT114), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1077), .A2(KEYINPUT114), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n757), .B(new_n760), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n736), .B2(G1996), .ZN(new_n1081));
  AOI211_X1 g656(.A(new_n1078), .B(new_n1079), .C1(new_n1076), .C2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1076), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n697), .B(new_n700), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n572), .A2(new_n662), .ZN(new_n1086));
  NAND2_X1  g661(.A1(G290), .A2(G1986), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1083), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1075), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1083), .A2(G1996), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT46), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1091), .B(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n732), .A2(new_n1080), .A3(new_n735), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1083), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT47), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1095), .B(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT48), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1085), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n698), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(new_n700), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1082), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n758), .A2(new_n760), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1083), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1097), .A2(new_n1100), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1090), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT127), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT127), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1090), .A2(new_n1106), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g686(.A1(new_n882), .A2(new_n854), .A3(G319), .A4(new_n889), .ZN(new_n1113));
  OR2_X1    g687(.A1(G401), .A2(G227), .ZN(new_n1114));
  NOR3_X1   g688(.A1(new_n1113), .A2(G229), .A3(new_n1114), .ZN(G308));
  INV_X1    g689(.A(G308), .ZN(G225));
endmodule


