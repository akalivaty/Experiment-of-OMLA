//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G176gat), .B(G204gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  NAND2_X1  g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT7), .ZN(new_n206));
  INV_X1    g005(.A(G99gat), .ZN(new_n207));
  INV_X1    g006(.A(G106gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT8), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(KEYINPUT99), .B(G85gat), .Z(new_n210));
  OAI211_X1 g009(.A(new_n206), .B(new_n209), .C1(G92gat), .C2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G99gat), .B(G106gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214));
  XNOR2_X1  g013(.A(G57gat), .B(G64gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(KEYINPUT96), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(KEYINPUT96), .B2(new_n215), .ZN(new_n217));
  OR2_X1    g016(.A1(G71gat), .A2(G78gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G71gat), .A2(G78gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n215), .B(KEYINPUT97), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n218), .B2(new_n214), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n217), .A2(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n213), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n213), .A2(new_n223), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT101), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n224), .B1(new_n227), .B2(KEYINPUT10), .ZN(new_n228));
  NAND2_X1  g027(.A1(G230gat), .A2(G233gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT10), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n232), .A2(KEYINPUT104), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(KEYINPUT104), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n213), .A2(new_n223), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n229), .B1(new_n236), .B2(new_n225), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(KEYINPUT103), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n204), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT105), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT106), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n232), .A2(KEYINPUT102), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n232), .A2(KEYINPUT102), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n243), .A2(new_n244), .A3(new_n204), .A4(new_n238), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n241), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n242), .B1(new_n241), .B2(new_n245), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G43gat), .B(G50gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT89), .B(KEYINPUT15), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(KEYINPUT15), .ZN(new_n253));
  NAND2_X1  g052(.A1(G29gat), .A2(G36gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT14), .ZN(new_n255));
  INV_X1    g054(.A(G29gat), .ZN(new_n256));
  INV_X1    g055(.A(G36gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n252), .A2(new_n253), .A3(new_n254), .A4(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n258), .A2(KEYINPUT87), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT87), .ZN(new_n263));
  NOR2_X1   g062(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n263), .B1(new_n264), .B2(new_n257), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n259), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT88), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n254), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n266), .A2(new_n267), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n261), .B1(new_n271), .B2(new_n253), .ZN(new_n272));
  NAND2_X1  g071(.A1(KEYINPUT90), .A2(KEYINPUT17), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(KEYINPUT90), .A2(KEYINPUT17), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n213), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G190gat), .B(G218gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT100), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT41), .ZN(new_n281));
  NAND2_X1  g080(.A1(G232gat), .A2(G233gat), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n283), .B1(new_n272), .B2(new_n213), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n279), .A2(KEYINPUT100), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G134gat), .B(G162gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n282), .A2(new_n281), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n288), .B(new_n289), .Z(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n287), .A2(new_n291), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n223), .A2(KEYINPUT21), .ZN(new_n296));
  NAND2_X1  g095(.A1(G231gat), .A2(G233gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G127gat), .B(G155gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT98), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n298), .B(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G183gat), .B(G211gat), .Z(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G8gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(G15gat), .B(G22gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT91), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n306), .A2(G1gat), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n304), .B1(new_n307), .B2(KEYINPUT92), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT16), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n306), .B1(new_n309), .B2(G1gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n311), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(KEYINPUT21), .B2(new_n223), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n303), .B(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n295), .A2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n249), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT95), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n314), .A2(new_n272), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT93), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n276), .A2(new_n312), .A3(new_n313), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G229gat), .A2(G233gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(KEYINPUT18), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n324), .B1(new_n272), .B2(new_n314), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(new_n327), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n324), .A2(new_n327), .A3(new_n325), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT18), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n328), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G113gat), .B(G141gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(G197gat), .ZN(new_n338));
  XOR2_X1   g137(.A(KEYINPUT11), .B(G169gat), .Z(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n340), .B(KEYINPUT12), .Z(new_n341));
  NAND2_X1  g140(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n341), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n328), .A2(new_n343), .A3(new_n332), .A4(new_n335), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n348));
  NAND2_X1  g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT2), .ZN(new_n350));
  INV_X1    g149(.A(G141gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(G148gat), .ZN(new_n352));
  INV_X1    g151(.A(G148gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n353), .A2(G141gat), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n348), .B(new_n350), .C1(new_n352), .C2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G155gat), .B(G162gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n353), .A2(G141gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n351), .A2(G148gat), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT75), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n361), .A2(new_n356), .A3(new_n350), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT3), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n358), .A2(new_n365), .A3(new_n362), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(G127gat), .A2(G134gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(G127gat), .A2(G134gat), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT1), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  AND2_X1   g170(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n373));
  INV_X1    g172(.A(G120gat), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(G113gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT70), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  OR2_X1    g177(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(G120gat), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT70), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n382), .A3(new_n376), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n371), .B1(new_n378), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G113gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G120gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n376), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT1), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT68), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(G134gat), .ZN(new_n391));
  INV_X1    g190(.A(G134gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(KEYINPUT68), .ZN(new_n393));
  OAI21_X1  g192(.A(G127gat), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n389), .A2(new_n394), .A3(new_n368), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n384), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n347), .B1(new_n367), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n398), .A2(KEYINPUT5), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n358), .A3(new_n362), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n381), .A2(new_n382), .A3(new_n376), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n382), .B1(new_n381), .B2(new_n376), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n370), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT4), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT76), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n406), .B1(new_n384), .B2(new_n400), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n359), .A2(new_n360), .ZN(new_n408));
  AND4_X1   g207(.A1(new_n348), .A2(new_n408), .A3(new_n356), .A4(new_n350), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n356), .B1(new_n361), .B2(new_n350), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n404), .A2(new_n411), .A3(KEYINPUT76), .A4(new_n395), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n405), .B1(new_n413), .B2(KEYINPUT4), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT77), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n413), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n398), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT4), .B1(new_n407), .B2(new_n412), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n384), .A2(new_n400), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT77), .B1(new_n422), .B2(new_n417), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT5), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n363), .B1(new_n384), .B2(new_n396), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n407), .A2(new_n412), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n347), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(KEYINPUT78), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT78), .B1(new_n427), .B2(new_n428), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n415), .B1(new_n425), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G1gat), .B(G29gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT0), .ZN(new_n435));
  XNOR2_X1  g234(.A(G57gat), .B(G85gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(KEYINPUT6), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT6), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n433), .A2(new_n437), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT79), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n437), .B1(new_n399), .B2(new_n414), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n442), .B(new_n443), .C1(new_n425), .C2(new_n432), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n427), .A2(new_n428), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT78), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n429), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n418), .B(new_n419), .C1(new_n421), .C2(new_n423), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(KEYINPUT5), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n442), .B1(new_n451), .B2(new_n443), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n440), .B(new_n441), .C1(new_n445), .C2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n439), .B1(new_n453), .B2(KEYINPUT80), .ZN(new_n454));
  INV_X1    g253(.A(new_n452), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n444), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT80), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n440), .A4(new_n441), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G197gat), .B(G204gat), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT22), .ZN(new_n461));
  INV_X1    g260(.A(G211gat), .ZN(new_n462));
  INV_X1    g261(.A(G218gat), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(G211gat), .B(G218gat), .Z(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G226gat), .A2(G233gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT73), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G190gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT65), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT65), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(G190gat), .ZN(new_n474));
  INV_X1    g273(.A(G183gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT27), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT27), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(G183gat), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n472), .A2(new_n474), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(KEYINPUT66), .B(KEYINPUT28), .Z(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT67), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n472), .A2(new_n474), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT27), .B(G183gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT28), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT67), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n479), .A2(new_n486), .A3(new_n480), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G183gat), .A2(G190gat), .ZN(new_n489));
  INV_X1    g288(.A(G169gat), .ZN(new_n490));
  INV_X1    g289(.A(G176gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT26), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G169gat), .A2(G176gat), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT26), .B1(new_n490), .B2(new_n491), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT24), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n489), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n475), .A2(new_n471), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT23), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT23), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(G169gat), .B2(G176gat), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n502), .A2(new_n495), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT25), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT64), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n500), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n509), .A2(new_n499), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n503), .A2(new_n505), .A3(new_n495), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(KEYINPUT25), .A3(new_n514), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n488), .A2(new_n497), .B1(new_n508), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n470), .B1(new_n516), .B2(KEYINPUT29), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT74), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n487), .A2(new_n485), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n486), .B1(new_n479), .B2(new_n480), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n497), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n515), .A2(new_n508), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n518), .B1(new_n523), .B2(new_n469), .ZN(new_n524));
  AOI211_X1 g323(.A(KEYINPUT74), .B(new_n470), .C1(new_n521), .C2(new_n522), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n467), .B(new_n517), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n467), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT29), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n469), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n516), .A2(new_n470), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G8gat), .B(G36gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(G64gat), .B(G92gat), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n532), .B(new_n533), .Z(new_n534));
  AND3_X1   g333(.A1(new_n526), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n534), .B1(new_n526), .B2(new_n531), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n526), .A2(new_n531), .ZN(new_n539));
  INV_X1    g338(.A(new_n534), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n539), .A2(KEYINPUT30), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n459), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G50gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n366), .A2(new_n528), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n527), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT3), .B1(new_n467), .B2(new_n528), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(new_n548), .B2(new_n411), .ZN(new_n549));
  INV_X1    g348(.A(G228gat), .ZN(new_n550));
  INV_X1    g349(.A(G233gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT81), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n465), .A2(new_n555), .A3(new_n466), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n528), .B(new_n556), .C1(new_n467), .C2(new_n555), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n411), .B1(new_n557), .B2(new_n365), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n545), .B1(new_n554), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G78gat), .B(G106gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G22gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n545), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n553), .B(new_n564), .C1(new_n558), .C2(new_n559), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n561), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n563), .B1(new_n561), .B2(new_n565), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n544), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n516), .B1(new_n384), .B2(new_n396), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n523), .A2(new_n397), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G227gat), .A2(G233gat), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT71), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n571), .A2(G227gat), .A3(G233gat), .A4(new_n572), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT32), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n577), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT33), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G15gat), .B(G43gat), .Z(new_n583));
  XNOR2_X1  g382(.A(G71gat), .B(G99gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n587), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n582), .A2(new_n590), .A3(new_n585), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n580), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n588), .A2(new_n578), .A3(new_n579), .A4(new_n591), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n593), .A2(KEYINPUT36), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT36), .B1(new_n593), .B2(new_n594), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n407), .A2(new_n412), .A3(new_n426), .A4(new_n347), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT83), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n364), .B(new_n366), .C1(new_n384), .C2(new_n396), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n414), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n600), .B(KEYINPUT39), .C1(new_n602), .C2(new_n347), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n437), .B(KEYINPUT82), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n347), .B1(new_n414), .B2(new_n601), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n603), .A2(KEYINPUT40), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT40), .B1(new_n603), .B2(new_n607), .ZN(new_n609));
  INV_X1    g408(.A(new_n604), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n610), .B1(new_n451), .B2(new_n415), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n569), .B1(new_n612), .B2(new_n542), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n433), .A2(new_n604), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n440), .B(new_n614), .C1(new_n445), .C2(new_n452), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n540), .B1(new_n539), .B2(KEYINPUT37), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT37), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n617), .B1(new_n526), .B2(new_n531), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT38), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n517), .B(new_n467), .C1(new_n470), .C2(new_n516), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT74), .B1(new_n516), .B2(new_n470), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n523), .A2(new_n518), .A3(new_n469), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n529), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI211_X1 g422(.A(KEYINPUT84), .B(new_n620), .C1(new_n623), .C2(new_n467), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n529), .A2(new_n530), .A3(new_n527), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT84), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n617), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT38), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n526), .A2(new_n531), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n534), .B1(new_n629), .B2(new_n617), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n535), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n615), .A2(new_n438), .A3(new_n619), .A4(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n613), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT85), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n597), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n613), .A2(KEYINPUT85), .A3(new_n632), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n570), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n593), .A2(new_n568), .A3(new_n594), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(KEYINPUT35), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT86), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n615), .A2(new_n438), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n640), .B1(new_n641), .B2(new_n543), .ZN(new_n642));
  AOI211_X1 g441(.A(KEYINPUT86), .B(new_n542), .C1(new_n615), .C2(new_n438), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI211_X1 g443(.A(new_n542), .B(new_n638), .C1(new_n454), .C2(new_n458), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT35), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI211_X1 g446(.A(new_n321), .B(new_n346), .C1(new_n637), .C2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n415), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT5), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n398), .B1(new_n421), .B2(new_n416), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n413), .A2(new_n417), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n401), .A2(new_n404), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n416), .B1(new_n653), .B2(KEYINPUT4), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n650), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n649), .B1(new_n656), .B2(new_n449), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n440), .B1(new_n657), .B2(new_n610), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n658), .B1(new_n455), .B2(new_n444), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n628), .A2(new_n630), .ZN(new_n660));
  INV_X1    g459(.A(new_n535), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(new_n619), .A3(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n659), .A2(new_n662), .A3(new_n439), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n603), .A2(new_n607), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n603), .A2(KEYINPUT40), .A3(new_n607), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n614), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n568), .B1(new_n668), .B2(new_n543), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n634), .B1(new_n663), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n597), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(new_n636), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n542), .B1(new_n454), .B2(new_n458), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n568), .ZN(new_n674));
  INV_X1    g473(.A(new_n638), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n646), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n646), .ZN(new_n677));
  INV_X1    g476(.A(new_n658), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n439), .B1(new_n456), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT86), .B1(new_n679), .B2(new_n542), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n641), .A2(new_n640), .A3(new_n543), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n677), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI22_X1  g481(.A1(new_n672), .A2(new_n674), .B1(new_n676), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT95), .B1(new_n683), .B2(new_n345), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n320), .B1(new_n648), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT107), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n687), .B(new_n320), .C1(new_n648), .C2(new_n684), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n459), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g491(.A(KEYINPUT16), .B(G8gat), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n689), .A2(new_n542), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n304), .A2(KEYINPUT42), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n693), .A2(new_n694), .ZN(new_n699));
  AND4_X1   g498(.A1(KEYINPUT108), .A2(new_n689), .A3(new_n542), .A4(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n543), .B1(new_n686), .B2(new_n688), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT108), .B1(new_n701), .B2(new_n699), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n698), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT109), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g504(.A(KEYINPUT109), .B(new_n698), .C1(new_n700), .C2(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1325gat));
  INV_X1    g506(.A(new_n689), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n593), .A2(new_n594), .ZN(new_n709));
  OR3_X1    g508(.A1(new_n708), .A2(G15gat), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(G15gat), .B1(new_n708), .B2(new_n671), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1326gat));
  XNOR2_X1  g511(.A(KEYINPUT43), .B(G22gat), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n689), .A2(new_n569), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT110), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n715), .A2(KEYINPUT110), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n714), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n718), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(new_n716), .A3(new_n713), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(G1327gat));
  OR2_X1    g521(.A1(new_n648), .A2(new_n684), .ZN(new_n723));
  INV_X1    g522(.A(new_n249), .ZN(new_n724));
  INV_X1    g523(.A(new_n318), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n724), .A2(new_n725), .A3(new_n294), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(new_n256), .A3(new_n690), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT45), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n294), .B1(new_n637), .B2(new_n647), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n731), .A2(KEYINPUT44), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(KEYINPUT44), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n724), .A2(new_n346), .A3(new_n725), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n737), .A2(new_n690), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n730), .B1(new_n256), .B2(new_n739), .ZN(G1328gat));
  NOR3_X1   g539(.A1(new_n727), .A2(G36gat), .A3(new_n543), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT46), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n737), .A2(new_n542), .A3(new_n738), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n257), .B2(new_n743), .ZN(G1329gat));
  NOR3_X1   g543(.A1(new_n727), .A2(G43gat), .A3(new_n709), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G43gat), .B1(new_n735), .B2(new_n671), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n746), .A2(KEYINPUT47), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n737), .A2(new_n597), .A3(new_n738), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n745), .B1(new_n749), .B2(G43gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n750), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g550(.A1(new_n727), .A2(G50gat), .A3(new_n568), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G50gat), .B1(new_n735), .B2(new_n568), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(KEYINPUT48), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n737), .A2(new_n569), .A3(new_n738), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n752), .B1(new_n756), .B2(G50gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n757), .B2(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g557(.A1(new_n346), .A2(new_n724), .A3(new_n683), .A4(new_n319), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n690), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n542), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n763));
  XOR2_X1   g562(.A(KEYINPUT49), .B(G64gat), .Z(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n762), .B2(new_n764), .ZN(G1333gat));
  NAND2_X1  g564(.A1(new_n759), .A2(new_n597), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n709), .A2(G71gat), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n766), .A2(G71gat), .B1(new_n759), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1334gat));
  NAND2_X1  g569(.A1(new_n759), .A2(new_n569), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g571(.A1(new_n345), .A2(new_n725), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n731), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT114), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT51), .B1(new_n731), .B2(new_n773), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n731), .A2(new_n779), .A3(KEYINPUT51), .A4(new_n773), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n776), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(KEYINPUT115), .Z(new_n782));
  NOR3_X1   g581(.A1(new_n249), .A2(new_n459), .A3(new_n210), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n732), .A2(new_n724), .A3(new_n733), .A4(new_n773), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n785), .A2(KEYINPUT113), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(KEYINPUT113), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(new_n690), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n210), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n784), .A2(new_n789), .ZN(G1336gat));
  NOR3_X1   g589(.A1(new_n249), .A2(G92gat), .A3(new_n543), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n781), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(G92gat), .B1(new_n785), .B2(new_n543), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n786), .A2(new_n542), .A3(new_n787), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n774), .A2(new_n775), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n797), .A2(new_n777), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n796), .A2(G92gat), .B1(new_n798), .B2(new_n791), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n795), .B1(new_n799), .B2(new_n794), .ZN(G1337gat));
  NOR3_X1   g599(.A1(new_n249), .A2(G99gat), .A3(new_n709), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n782), .A2(new_n801), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n786), .A2(new_n597), .A3(new_n787), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n207), .B2(new_n803), .ZN(G1338gat));
  NOR3_X1   g603(.A1(new_n249), .A2(G106gat), .A3(new_n568), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n781), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(G106gat), .B1(new_n785), .B2(new_n568), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT117), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n805), .B1(new_n797), .B2(new_n777), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n786), .A2(new_n569), .A3(new_n787), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(G106gat), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n810), .B1(new_n815), .B2(new_n808), .ZN(G1339gat));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n228), .A2(new_n231), .ZN(new_n818));
  INV_X1    g617(.A(new_n229), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n243), .A2(new_n244), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n204), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n821), .B(new_n822), .C1(KEYINPUT54), .C2(new_n235), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n245), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n326), .A2(new_n327), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n329), .A2(new_n331), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n340), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n344), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n295), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n318), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n344), .B(new_n830), .C1(new_n247), .C2(new_n248), .ZN(new_n834));
  INV_X1    g633(.A(new_n827), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n295), .B1(new_n835), .B2(new_n345), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n833), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n294), .A2(new_n725), .ZN(new_n838));
  NOR4_X1   g637(.A1(new_n247), .A2(new_n248), .A3(new_n838), .A4(new_n345), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n690), .A2(new_n543), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n840), .A2(new_n638), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n345), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n843), .B1(new_n379), .B2(new_n380), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(new_n385), .B2(new_n843), .ZN(G1340gat));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n724), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g646(.A1(new_n842), .A2(new_n725), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g648(.A1(new_n840), .A2(new_n638), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n294), .A2(new_n542), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n459), .A2(new_n391), .A3(new_n393), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(KEYINPUT56), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT118), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n850), .A2(new_n690), .A3(new_n851), .ZN(new_n856));
  AOI22_X1  g655(.A1(KEYINPUT56), .A2(new_n853), .B1(new_n856), .B2(G134gat), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(G1343gat));
  NAND2_X1  g657(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n837), .A2(new_n839), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n841), .A2(new_n597), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n569), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n345), .A2(new_n351), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n865), .B1(new_n840), .B2(new_n568), .ZN(new_n866));
  OAI211_X1 g665(.A(KEYINPUT57), .B(new_n569), .C1(new_n837), .C2(new_n839), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n861), .B(KEYINPUT119), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n868), .A2(new_n345), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n864), .B1(new_n871), .B2(G141gat), .ZN(new_n872));
  NOR2_X1   g671(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  AOI211_X1 g674(.A(new_n873), .B(new_n864), .C1(new_n871), .C2(G141gat), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(G1344gat));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n866), .A2(new_n879), .A3(new_n867), .ZN(new_n880));
  OAI211_X1 g679(.A(KEYINPUT122), .B(new_n865), .C1(new_n840), .C2(new_n568), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n869), .B(KEYINPUT121), .Z(new_n882));
  NAND4_X1  g681(.A1(new_n880), .A2(new_n724), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n878), .B1(new_n883), .B2(G148gat), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n869), .B1(new_n866), .B2(new_n867), .ZN(new_n885));
  AOI211_X1 g684(.A(KEYINPUT59), .B(new_n353), .C1(new_n885), .C2(new_n724), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n724), .A2(new_n353), .ZN(new_n887));
  OAI22_X1  g686(.A1(new_n884), .A2(new_n886), .B1(new_n862), .B2(new_n887), .ZN(G1345gat));
  NAND3_X1  g687(.A1(new_n885), .A2(G155gat), .A3(new_n725), .ZN(new_n889));
  INV_X1    g688(.A(G155gat), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n860), .A2(new_n569), .A3(new_n725), .A4(new_n861), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n889), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n889), .B(KEYINPUT124), .C1(new_n893), .C2(new_n894), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1346gat));
  INV_X1    g698(.A(G162gat), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n900), .B1(new_n885), .B2(new_n295), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n851), .A2(new_n900), .A3(new_n671), .ZN(new_n902));
  NOR4_X1   g701(.A1(new_n840), .A2(new_n459), .A3(new_n568), .A4(new_n902), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n901), .A2(new_n903), .ZN(G1347gat));
  NOR3_X1   g703(.A1(new_n690), .A2(new_n543), .A3(new_n638), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n860), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  OAI22_X1  g706(.A1(new_n907), .A2(new_n346), .B1(KEYINPUT125), .B2(G169gat), .ZN(new_n908));
  NAND2_X1  g707(.A1(KEYINPUT125), .A2(G169gat), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT126), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n908), .B(new_n910), .ZN(G1348gat));
  NAND2_X1  g710(.A1(new_n906), .A2(new_n724), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g712(.A1(new_n906), .A2(new_n725), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n914), .A2(G183gat), .B1(new_n915), .B2(KEYINPUT60), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n915), .A2(KEYINPUT60), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n906), .A2(new_n484), .A3(new_n725), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n917), .B1(new_n916), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(G1350gat));
  AOI21_X1  g720(.A(new_n471), .B1(new_n906), .B2(new_n295), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n922), .A2(KEYINPUT61), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(KEYINPUT61), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n483), .A3(new_n295), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G1351gat));
  NOR3_X1   g725(.A1(new_n690), .A2(new_n543), .A3(new_n597), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n860), .A2(new_n569), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(G197gat), .B1(new_n928), .B2(new_n345), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n880), .A2(new_n881), .A3(new_n927), .ZN(new_n930));
  INV_X1    g729(.A(G197gat), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n346), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n929), .B1(new_n930), .B2(new_n932), .ZN(G1352gat));
  INV_X1    g732(.A(G204gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n928), .A2(new_n934), .A3(new_n724), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT62), .Z(new_n936));
  NAND2_X1  g735(.A1(new_n930), .A2(new_n724), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G204gat), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1353gat));
  NAND3_X1  g738(.A1(new_n928), .A2(new_n462), .A3(new_n725), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n880), .A2(new_n725), .A3(new_n881), .A4(new_n927), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n941), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT63), .B1(new_n941), .B2(G211gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(G1354gat));
  NAND3_X1  g743(.A1(new_n928), .A2(new_n463), .A3(new_n295), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n930), .A2(new_n295), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n946), .B2(new_n463), .ZN(G1355gat));
endmodule


