

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581;

  XOR2_X1 U323 ( .A(n355), .B(n298), .Z(n291) );
  INV_X1 U324 ( .A(KEYINPUT71), .ZN(n302) );
  XNOR2_X1 U325 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U326 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n408) );
  XNOR2_X1 U327 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U328 ( .A(n409), .B(n408), .ZN(n530) );
  NOR2_X1 U329 ( .A1(n471), .A2(n444), .ZN(n563) );
  NOR2_X1 U330 ( .A1(n517), .A2(n508), .ZN(n514) );
  XNOR2_X1 U331 ( .A(KEYINPUT28), .B(n468), .ZN(n534) );
  XNOR2_X1 U332 ( .A(n445), .B(G176GAT), .ZN(n446) );
  XNOR2_X1 U333 ( .A(n447), .B(n446), .ZN(G1349GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n293) );
  XNOR2_X1 U335 ( .A(G71GAT), .B(G57GAT), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n393) );
  XOR2_X1 U337 ( .A(G64GAT), .B(G92GAT), .Z(n295) );
  XNOR2_X1 U338 ( .A(G176GAT), .B(G204GAT), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n295), .B(n294), .ZN(n417) );
  XNOR2_X1 U340 ( .A(n393), .B(n417), .ZN(n307) );
  XOR2_X1 U341 ( .A(G99GAT), .B(G85GAT), .Z(n355) );
  XOR2_X1 U342 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n297) );
  XNOR2_X1 U343 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n298) );
  NAND2_X1 U345 ( .A1(G230GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n291), .B(n299), .ZN(n305) );
  XOR2_X1 U347 ( .A(G78GAT), .B(G148GAT), .Z(n301) );
  XNOR2_X1 U348 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n335) );
  XNOR2_X1 U350 ( .A(n335), .B(KEYINPUT33), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n307), .B(n306), .ZN(n455) );
  XNOR2_X1 U352 ( .A(KEYINPUT41), .B(n455), .ZN(n549) );
  XNOR2_X1 U353 ( .A(KEYINPUT108), .B(n549), .ZN(n537) );
  XOR2_X1 U354 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n309) );
  XNOR2_X1 U355 ( .A(KEYINPUT82), .B(G183GAT), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U357 ( .A(KEYINPUT17), .B(n310), .Z(n414) );
  XOR2_X1 U358 ( .A(KEYINPUT65), .B(G99GAT), .Z(n312) );
  XNOR2_X1 U359 ( .A(G43GAT), .B(G190GAT), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U361 ( .A(G176GAT), .B(KEYINPUT20), .Z(n314) );
  XNOR2_X1 U362 ( .A(KEYINPUT83), .B(KEYINPUT81), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U364 ( .A(n316), .B(n315), .Z(n321) );
  XOR2_X1 U365 ( .A(G15GAT), .B(G71GAT), .Z(n318) );
  NAND2_X1 U366 ( .A1(G227GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U368 ( .A(G169GAT), .B(n319), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n414), .B(n322), .ZN(n326) );
  XOR2_X1 U371 ( .A(G127GAT), .B(G134GAT), .Z(n324) );
  XNOR2_X1 U372 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U374 ( .A(G113GAT), .B(n325), .Z(n427) );
  XNOR2_X1 U375 ( .A(n326), .B(n427), .ZN(n531) );
  INV_X1 U376 ( .A(n531), .ZN(n471) );
  XNOR2_X1 U377 ( .A(G211GAT), .B(KEYINPUT87), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n327), .B(KEYINPUT21), .ZN(n328) );
  XOR2_X1 U379 ( .A(n328), .B(KEYINPUT86), .Z(n330) );
  XNOR2_X1 U380 ( .A(G197GAT), .B(G218GAT), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n413) );
  XOR2_X1 U382 ( .A(KEYINPUT84), .B(G204GAT), .Z(n332) );
  NAND2_X1 U383 ( .A1(G228GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U385 ( .A(n333), .B(KEYINPUT85), .Z(n337) );
  XNOR2_X1 U386 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n334), .B(KEYINPUT2), .ZN(n437) );
  XNOR2_X1 U388 ( .A(n335), .B(n437), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U390 ( .A(KEYINPUT24), .B(KEYINPUT88), .Z(n339) );
  XNOR2_X1 U391 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n338) );
  XNOR2_X1 U392 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U393 ( .A(n341), .B(n340), .Z(n343) );
  XOR2_X1 U394 ( .A(G141GAT), .B(G22GAT), .Z(n362) );
  XOR2_X1 U395 ( .A(G50GAT), .B(G162GAT), .Z(n356) );
  XNOR2_X1 U396 ( .A(n362), .B(n356), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n413), .B(n344), .ZN(n468) );
  XOR2_X1 U399 ( .A(KEYINPUT9), .B(KEYINPUT74), .Z(n346) );
  XNOR2_X1 U400 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n360) );
  XOR2_X1 U402 ( .A(G36GAT), .B(G190GAT), .Z(n419) );
  XOR2_X1 U403 ( .A(G29GAT), .B(G43GAT), .Z(n348) );
  XNOR2_X1 U404 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n348), .B(n347), .ZN(n364) );
  XOR2_X1 U406 ( .A(n419), .B(n364), .Z(n350) );
  NAND2_X1 U407 ( .A1(G232GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U409 ( .A(G92GAT), .B(KEYINPUT10), .Z(n352) );
  XNOR2_X1 U410 ( .A(G134GAT), .B(G106GAT), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U412 ( .A(n354), .B(n353), .Z(n358) );
  XNOR2_X1 U413 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n564) );
  XNOR2_X1 U416 ( .A(G15GAT), .B(G1GAT), .ZN(n361) );
  XNOR2_X1 U417 ( .A(n361), .B(KEYINPUT67), .ZN(n394) );
  XNOR2_X1 U418 ( .A(n362), .B(n394), .ZN(n363) );
  XOR2_X1 U419 ( .A(G169GAT), .B(G8GAT), .Z(n420) );
  XNOR2_X1 U420 ( .A(n363), .B(n420), .ZN(n368) );
  XOR2_X1 U421 ( .A(n364), .B(KEYINPUT30), .Z(n366) );
  NAND2_X1 U422 ( .A1(G229GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U424 ( .A(n368), .B(n367), .Z(n376) );
  XOR2_X1 U425 ( .A(G197GAT), .B(G113GAT), .Z(n370) );
  XNOR2_X1 U426 ( .A(G36GAT), .B(G50GAT), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U428 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n372) );
  XNOR2_X1 U429 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n570) );
  NAND2_X1 U433 ( .A1(n570), .A2(n549), .ZN(n377) );
  XNOR2_X1 U434 ( .A(KEYINPUT46), .B(n377), .ZN(n397) );
  XOR2_X1 U435 ( .A(G78GAT), .B(G211GAT), .Z(n379) );
  XNOR2_X1 U436 ( .A(G183GAT), .B(G127GAT), .ZN(n378) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U438 ( .A(KEYINPUT76), .B(G64GAT), .Z(n381) );
  XNOR2_X1 U439 ( .A(G22GAT), .B(G155GAT), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U441 ( .A(n383), .B(n382), .Z(n388) );
  XOR2_X1 U442 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n385) );
  NAND2_X1 U443 ( .A1(G231GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U445 ( .A(KEYINPUT12), .B(n386), .ZN(n387) );
  XNOR2_X1 U446 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U447 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n390) );
  XNOR2_X1 U448 ( .A(G8GAT), .B(KEYINPUT75), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U450 ( .A(n392), .B(n391), .Z(n396) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n396), .B(n395), .ZN(n490) );
  NAND2_X1 U453 ( .A1(n397), .A2(n490), .ZN(n398) );
  XNOR2_X1 U454 ( .A(KEYINPUT112), .B(n398), .ZN(n399) );
  NOR2_X1 U455 ( .A1(n564), .A2(n399), .ZN(n401) );
  XNOR2_X1 U456 ( .A(KEYINPUT113), .B(KEYINPUT47), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n401), .B(n400), .ZN(n407) );
  INV_X1 U458 ( .A(n564), .ZN(n456) );
  XNOR2_X1 U459 ( .A(n456), .B(KEYINPUT36), .ZN(n578) );
  NOR2_X1 U460 ( .A1(n490), .A2(n578), .ZN(n402) );
  XNOR2_X1 U461 ( .A(KEYINPUT45), .B(n402), .ZN(n403) );
  NAND2_X1 U462 ( .A1(n403), .A2(n455), .ZN(n404) );
  NOR2_X1 U463 ( .A1(n570), .A2(n404), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n405), .B(KEYINPUT114), .ZN(n406) );
  NOR2_X1 U465 ( .A1(n407), .A2(n406), .ZN(n409) );
  XOR2_X1 U466 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n411) );
  NAND2_X1 U467 ( .A1(G226GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U469 ( .A(n412), .B(KEYINPUT94), .Z(n416) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n416), .B(n415), .ZN(n418) );
  XOR2_X1 U472 ( .A(n418), .B(n417), .Z(n422) );
  XNOR2_X1 U473 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U474 ( .A(n422), .B(n421), .ZN(n479) );
  NOR2_X1 U475 ( .A1(n530), .A2(n479), .ZN(n423) );
  XNOR2_X1 U476 ( .A(n423), .B(KEYINPUT54), .ZN(n442) );
  XOR2_X1 U477 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n425) );
  XNOR2_X1 U478 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n441) );
  XOR2_X1 U481 ( .A(G57GAT), .B(G148GAT), .Z(n429) );
  XNOR2_X1 U482 ( .A(G29GAT), .B(G141GAT), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U484 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n431) );
  XNOR2_X1 U485 ( .A(G1GAT), .B(KEYINPUT89), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U487 ( .A(n433), .B(n432), .Z(n439) );
  XOR2_X1 U488 ( .A(G85GAT), .B(G162GAT), .Z(n435) );
  NAND2_X1 U489 ( .A1(G225GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n469) );
  NAND2_X1 U494 ( .A1(n442), .A2(n469), .ZN(n449) );
  NOR2_X1 U495 ( .A1(n468), .A2(n449), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n443), .B(KEYINPUT55), .ZN(n444) );
  NAND2_X1 U497 ( .A1(n537), .A2(n563), .ZN(n447) );
  XOR2_X1 U498 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n445) );
  INV_X1 U499 ( .A(G204GAT), .ZN(n454) );
  XOR2_X1 U500 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n452) );
  NAND2_X1 U501 ( .A1(n468), .A2(n471), .ZN(n448) );
  XOR2_X1 U502 ( .A(n448), .B(KEYINPUT26), .Z(n547) );
  INV_X1 U503 ( .A(n547), .ZN(n450) );
  NOR2_X1 U504 ( .A1(n450), .A2(n449), .ZN(n573) );
  INV_X1 U505 ( .A(n573), .ZN(n577) );
  OR2_X1 U506 ( .A1(n577), .A2(n455), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n454), .B(n453), .ZN(G1353GAT) );
  XOR2_X1 U509 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n477) );
  NAND2_X1 U510 ( .A1(n570), .A2(n455), .ZN(n494) );
  INV_X1 U511 ( .A(n490), .ZN(n574) );
  NAND2_X1 U512 ( .A1(n574), .A2(n456), .ZN(n459) );
  XNOR2_X1 U513 ( .A(KEYINPUT16), .B(KEYINPUT80), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n457), .B(KEYINPUT79), .ZN(n458) );
  XNOR2_X1 U515 ( .A(n459), .B(n458), .ZN(n475) );
  NOR2_X1 U516 ( .A1(n479), .A2(n471), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n460), .B(KEYINPUT96), .ZN(n461) );
  NOR2_X1 U518 ( .A1(n468), .A2(n461), .ZN(n462) );
  XOR2_X1 U519 ( .A(n462), .B(KEYINPUT97), .Z(n463) );
  XNOR2_X1 U520 ( .A(KEYINPUT25), .B(n463), .ZN(n466) );
  XOR2_X1 U521 ( .A(n479), .B(KEYINPUT27), .Z(n470) );
  NAND2_X1 U522 ( .A1(n470), .A2(n547), .ZN(n464) );
  XOR2_X1 U523 ( .A(KEYINPUT95), .B(n464), .Z(n465) );
  NAND2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U525 ( .A1(n467), .A2(n469), .ZN(n474) );
  INV_X1 U526 ( .A(n469), .ZN(n519) );
  NAND2_X1 U527 ( .A1(n470), .A2(n519), .ZN(n529) );
  NOR2_X1 U528 ( .A1(n534), .A2(n529), .ZN(n472) );
  NAND2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U530 ( .A1(n474), .A2(n473), .ZN(n489) );
  NAND2_X1 U531 ( .A1(n475), .A2(n489), .ZN(n508) );
  NOR2_X1 U532 ( .A1(n494), .A2(n508), .ZN(n486) );
  NAND2_X1 U533 ( .A1(n486), .A2(n519), .ZN(n476) );
  XNOR2_X1 U534 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U535 ( .A(G1GAT), .B(n478), .Z(G1324GAT) );
  XOR2_X1 U536 ( .A(G8GAT), .B(KEYINPUT99), .Z(n481) );
  INV_X1 U537 ( .A(n479), .ZN(n521) );
  NAND2_X1 U538 ( .A1(n486), .A2(n521), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n483) );
  NAND2_X1 U541 ( .A1(n486), .A2(n531), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n485) );
  XOR2_X1 U543 ( .A(G15GAT), .B(KEYINPUT100), .Z(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NAND2_X1 U545 ( .A1(n486), .A2(n534), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n487), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT39), .Z(n498) );
  XNOR2_X1 U548 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n488), .B(KEYINPUT38), .ZN(n496) );
  NAND2_X1 U550 ( .A1(n490), .A2(n489), .ZN(n491) );
  NOR2_X1 U551 ( .A1(n491), .A2(n578), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(KEYINPUT102), .ZN(n493) );
  XNOR2_X1 U553 ( .A(KEYINPUT37), .B(n493), .ZN(n518) );
  NOR2_X1 U554 ( .A1(n518), .A2(n494), .ZN(n495) );
  XOR2_X1 U555 ( .A(n496), .B(n495), .Z(n504) );
  NAND2_X1 U556 ( .A1(n504), .A2(n519), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n504), .A2(n521), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(n499), .ZN(G1329GAT) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n503) );
  XOR2_X1 U561 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n501) );
  NAND2_X1 U562 ( .A1(n504), .A2(n531), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(G1330GAT) );
  XOR2_X1 U565 ( .A(G50GAT), .B(KEYINPUT107), .Z(n506) );
  NAND2_X1 U566 ( .A1(n504), .A2(n534), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n506), .B(n505), .ZN(G1331GAT) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n510) );
  INV_X1 U569 ( .A(n570), .ZN(n507) );
  NAND2_X1 U570 ( .A1(n537), .A2(n507), .ZN(n517) );
  NAND2_X1 U571 ( .A1(n514), .A2(n519), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n510), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n521), .A2(n514), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U575 ( .A(G71GAT), .B(KEYINPUT109), .Z(n513) );
  NAND2_X1 U576 ( .A1(n514), .A2(n531), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U579 ( .A1(n514), .A2(n534), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NOR2_X1 U581 ( .A1(n518), .A2(n517), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n524), .A2(n519), .ZN(n520) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n521), .A2(n524), .ZN(n522) );
  XNOR2_X1 U585 ( .A(n522), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n524), .A2(n531), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n528) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n526) );
  NAND2_X1 U590 ( .A1(n524), .A2(n534), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(G1339GAT) );
  NOR2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n546) );
  NAND2_X1 U594 ( .A1(n531), .A2(n546), .ZN(n532) );
  XOR2_X1 U595 ( .A(KEYINPUT115), .B(n532), .Z(n533) );
  NOR2_X1 U596 ( .A1(n534), .A2(n533), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n542), .A2(n570), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n535), .B(KEYINPUT116), .ZN(n536) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n536), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U601 ( .A1(n542), .A2(n537), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  NAND2_X1 U603 ( .A1(n574), .A2(n542), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n540), .B(KEYINPUT50), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U607 ( .A1(n542), .A2(n564), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U609 ( .A(G134GAT), .B(n545), .Z(G1343GAT) );
  AND2_X1 U610 ( .A1(n547), .A2(n546), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n570), .A2(n556), .ZN(n548) );
  XNOR2_X1 U612 ( .A(G141GAT), .B(n548), .ZN(G1344GAT) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n553) );
  XOR2_X1 U614 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n551) );
  NAND2_X1 U615 ( .A1(n556), .A2(n549), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  XOR2_X1 U618 ( .A(G155GAT), .B(KEYINPUT119), .Z(n555) );
  NAND2_X1 U619 ( .A1(n556), .A2(n574), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n564), .A2(n556), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(KEYINPUT120), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G162GAT), .B(n558), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n570), .A2(n563), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(n559), .ZN(G1348GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n561) );
  NAND2_X1 U627 ( .A1(n563), .A2(n574), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(G183GAT), .B(n562), .ZN(G1350GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT58), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(n566), .ZN(G1351GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n568) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U636 ( .A(KEYINPUT123), .B(n569), .Z(n572) );
  NAND2_X1 U637 ( .A1(n573), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT126), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(n576), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

