

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581;

  XNOR2_X1 U325 ( .A(n353), .B(n377), .ZN(n354) );
  INV_X1 U326 ( .A(KEYINPUT68), .ZN(n318) );
  XNOR2_X1 U327 ( .A(n319), .B(n318), .ZN(n353) );
  XOR2_X1 U328 ( .A(KEYINPUT81), .B(n552), .Z(n560) );
  INV_X1 U329 ( .A(G183GAT), .ZN(n447) );
  XNOR2_X1 U330 ( .A(n447), .B(KEYINPUT124), .ZN(n448) );
  XNOR2_X1 U331 ( .A(n449), .B(n448), .ZN(G1350GAT) );
  XOR2_X1 U332 ( .A(G1GAT), .B(G8GAT), .Z(n309) );
  XOR2_X1 U333 ( .A(G22GAT), .B(G155GAT), .Z(n415) );
  XOR2_X1 U334 ( .A(n415), .B(KEYINPUT12), .Z(n294) );
  NAND2_X1 U335 ( .A1(G231GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U337 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n296) );
  XNOR2_X1 U338 ( .A(G64GAT), .B(KEYINPUT82), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U340 ( .A(n298), .B(n297), .Z(n303) );
  XOR2_X1 U341 ( .A(G15GAT), .B(G127GAT), .Z(n433) );
  XOR2_X1 U342 ( .A(G78GAT), .B(G211GAT), .Z(n300) );
  XNOR2_X1 U343 ( .A(G183GAT), .B(G71GAT), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n433), .B(n301), .ZN(n302) );
  XNOR2_X1 U346 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U347 ( .A(n309), .B(n304), .ZN(n305) );
  XOR2_X1 U348 ( .A(G57GAT), .B(KEYINPUT13), .Z(n329) );
  XNOR2_X1 U349 ( .A(n305), .B(n329), .ZN(n574) );
  XOR2_X1 U350 ( .A(G15GAT), .B(G113GAT), .Z(n307) );
  XNOR2_X1 U351 ( .A(G36GAT), .B(G50GAT), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U353 ( .A(n309), .B(n308), .Z(n311) );
  NAND2_X1 U354 ( .A1(G229GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U355 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U356 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n313) );
  XNOR2_X1 U357 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n312) );
  XNOR2_X1 U358 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U359 ( .A(n315), .B(n314), .Z(n324) );
  XOR2_X1 U360 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n317) );
  XNOR2_X1 U361 ( .A(G43GAT), .B(G29GAT), .ZN(n316) );
  XNOR2_X1 U362 ( .A(n317), .B(n316), .ZN(n319) );
  XOR2_X1 U363 ( .A(G22GAT), .B(G141GAT), .Z(n321) );
  XNOR2_X1 U364 ( .A(G169GAT), .B(G197GAT), .ZN(n320) );
  XNOR2_X1 U365 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U366 ( .A(n353), .B(n322), .ZN(n323) );
  XNOR2_X1 U367 ( .A(n324), .B(n323), .ZN(n567) );
  XOR2_X1 U368 ( .A(G78GAT), .B(G148GAT), .Z(n326) );
  XNOR2_X1 U369 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n325) );
  XNOR2_X1 U370 ( .A(n326), .B(n325), .ZN(n423) );
  XOR2_X1 U371 ( .A(KEYINPUT74), .B(G85GAT), .Z(n328) );
  XNOR2_X1 U372 ( .A(G99GAT), .B(G106GAT), .ZN(n327) );
  XNOR2_X1 U373 ( .A(n328), .B(n327), .ZN(n359) );
  XOR2_X1 U374 ( .A(n423), .B(n359), .Z(n342) );
  XOR2_X1 U375 ( .A(G176GAT), .B(G64GAT), .Z(n381) );
  XNOR2_X1 U376 ( .A(n381), .B(n329), .ZN(n331) );
  AND2_X1 U377 ( .A1(G230GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U378 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U379 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n333) );
  XNOR2_X1 U380 ( .A(KEYINPUT71), .B(KEYINPUT70), .ZN(n332) );
  XNOR2_X1 U381 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U382 ( .A(n335), .B(n334), .Z(n340) );
  XOR2_X1 U383 ( .A(G120GAT), .B(G71GAT), .Z(n432) );
  XOR2_X1 U384 ( .A(KEYINPUT31), .B(KEYINPUT75), .Z(n337) );
  XNOR2_X1 U385 ( .A(G204GAT), .B(G92GAT), .ZN(n336) );
  XNOR2_X1 U386 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U387 ( .A(n432), .B(n338), .ZN(n339) );
  XNOR2_X1 U388 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U389 ( .A(n342), .B(n341), .ZN(n571) );
  XOR2_X1 U390 ( .A(n571), .B(KEYINPUT64), .Z(n343) );
  XNOR2_X1 U391 ( .A(n343), .B(KEYINPUT41), .ZN(n555) );
  NOR2_X1 U392 ( .A1(n567), .A2(n555), .ZN(n344) );
  XNOR2_X1 U393 ( .A(n344), .B(KEYINPUT46), .ZN(n363) );
  NAND2_X1 U394 ( .A1(G232GAT), .A2(G233GAT), .ZN(n350) );
  XOR2_X1 U395 ( .A(KEYINPUT80), .B(KEYINPUT78), .Z(n346) );
  XNOR2_X1 U396 ( .A(KEYINPUT10), .B(KEYINPUT79), .ZN(n345) );
  XNOR2_X1 U397 ( .A(n346), .B(n345), .ZN(n348) );
  XOR2_X1 U398 ( .A(G134GAT), .B(KEYINPUT9), .Z(n347) );
  XNOR2_X1 U399 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U400 ( .A(n350), .B(n349), .ZN(n357) );
  XOR2_X1 U401 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n355) );
  XOR2_X1 U402 ( .A(G92GAT), .B(G218GAT), .Z(n352) );
  XNOR2_X1 U403 ( .A(G36GAT), .B(G190GAT), .ZN(n351) );
  XNOR2_X1 U404 ( .A(n352), .B(n351), .ZN(n377) );
  XNOR2_X1 U405 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U406 ( .A(n357), .B(n356), .ZN(n361) );
  XNOR2_X1 U407 ( .A(G50GAT), .B(KEYINPUT77), .ZN(n358) );
  XNOR2_X1 U408 ( .A(n358), .B(G162GAT), .ZN(n418) );
  XNOR2_X1 U409 ( .A(n418), .B(n359), .ZN(n360) );
  XNOR2_X1 U410 ( .A(n361), .B(n360), .ZN(n552) );
  NAND2_X1 U411 ( .A1(n574), .A2(n552), .ZN(n362) );
  OR2_X1 U412 ( .A1(n363), .A2(n362), .ZN(n364) );
  XNOR2_X1 U413 ( .A(KEYINPUT47), .B(n364), .ZN(n370) );
  XNOR2_X1 U414 ( .A(KEYINPUT36), .B(n560), .ZN(n579) );
  NOR2_X1 U415 ( .A1(n574), .A2(n579), .ZN(n366) );
  XNOR2_X1 U416 ( .A(KEYINPUT45), .B(KEYINPUT117), .ZN(n365) );
  XNOR2_X1 U417 ( .A(n366), .B(n365), .ZN(n368) );
  NAND2_X1 U418 ( .A1(n567), .A2(n571), .ZN(n367) );
  NOR2_X1 U419 ( .A1(n368), .A2(n367), .ZN(n369) );
  NOR2_X1 U420 ( .A1(n370), .A2(n369), .ZN(n371) );
  XNOR2_X1 U421 ( .A(n371), .B(KEYINPUT48), .ZN(n525) );
  XOR2_X1 U422 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n373) );
  NAND2_X1 U423 ( .A1(G226GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U424 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U425 ( .A(n374), .B(KEYINPUT91), .Z(n379) );
  XOR2_X1 U426 ( .A(G204GAT), .B(G211GAT), .Z(n376) );
  XNOR2_X1 U427 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n375) );
  XNOR2_X1 U428 ( .A(n376), .B(n375), .ZN(n424) );
  XNOR2_X1 U429 ( .A(n424), .B(n377), .ZN(n378) );
  XNOR2_X1 U430 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U431 ( .A(n380), .B(KEYINPUT94), .Z(n383) );
  XNOR2_X1 U432 ( .A(G8GAT), .B(n381), .ZN(n382) );
  XNOR2_X1 U433 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U434 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n385) );
  XNOR2_X1 U435 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n384) );
  XNOR2_X1 U436 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U437 ( .A(G169GAT), .B(n386), .ZN(n444) );
  XNOR2_X1 U438 ( .A(n387), .B(n444), .ZN(n515) );
  XNOR2_X1 U439 ( .A(n515), .B(KEYINPUT122), .ZN(n388) );
  NOR2_X1 U440 ( .A1(n525), .A2(n388), .ZN(n389) );
  XNOR2_X1 U441 ( .A(n389), .B(KEYINPUT54), .ZN(n410) );
  XOR2_X1 U442 ( .A(KEYINPUT88), .B(KEYINPUT90), .Z(n391) );
  XNOR2_X1 U443 ( .A(G1GAT), .B(KEYINPUT89), .ZN(n390) );
  XNOR2_X1 U444 ( .A(n391), .B(n390), .ZN(n409) );
  XOR2_X1 U445 ( .A(G162GAT), .B(G148GAT), .Z(n393) );
  XNOR2_X1 U446 ( .A(G127GAT), .B(G120GAT), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U448 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n395) );
  XNOR2_X1 U449 ( .A(G155GAT), .B(G57GAT), .ZN(n394) );
  XNOR2_X1 U450 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U451 ( .A(n397), .B(n396), .Z(n403) );
  XNOR2_X1 U452 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n398) );
  XNOR2_X1 U453 ( .A(n398), .B(KEYINPUT2), .ZN(n414) );
  XOR2_X1 U454 ( .A(G85GAT), .B(n414), .Z(n400) );
  NAND2_X1 U455 ( .A1(G225GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U457 ( .A(G29GAT), .B(n401), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U459 ( .A(n404), .B(KEYINPUT5), .Z(n407) );
  XNOR2_X1 U460 ( .A(G113GAT), .B(G134GAT), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n405), .B(KEYINPUT0), .ZN(n441) );
  XNOR2_X1 U462 ( .A(n441), .B(KEYINPUT4), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n511) );
  NAND2_X1 U465 ( .A1(n410), .A2(n511), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n411), .B(KEYINPUT65), .ZN(n566) );
  XOR2_X1 U467 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n413) );
  XNOR2_X1 U468 ( .A(KEYINPUT87), .B(KEYINPUT86), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n428) );
  XOR2_X1 U470 ( .A(n415), .B(n414), .Z(n417) );
  XNOR2_X1 U471 ( .A(G218GAT), .B(G106GAT), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n422) );
  XOR2_X1 U473 ( .A(n418), .B(KEYINPUT23), .Z(n420) );
  NAND2_X1 U474 ( .A1(G228GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U476 ( .A(n422), .B(n421), .Z(n426) );
  XNOR2_X1 U477 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U478 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U479 ( .A(n428), .B(n427), .Z(n459) );
  NAND2_X1 U480 ( .A1(n566), .A2(n459), .ZN(n429) );
  XNOR2_X1 U481 ( .A(n429), .B(KEYINPUT55), .ZN(n446) );
  XOR2_X1 U482 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n431) );
  XNOR2_X1 U483 ( .A(G99GAT), .B(G176GAT), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n437) );
  XOR2_X1 U485 ( .A(G190GAT), .B(n432), .Z(n435) );
  XNOR2_X1 U486 ( .A(G43GAT), .B(n433), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U488 ( .A(n437), .B(n436), .Z(n439) );
  NAND2_X1 U489 ( .A1(G227GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U491 ( .A(n440), .B(KEYINPUT84), .Z(n443) );
  XNOR2_X1 U492 ( .A(n441), .B(KEYINPUT83), .ZN(n442) );
  XNOR2_X1 U493 ( .A(n443), .B(n442), .ZN(n445) );
  XNOR2_X1 U494 ( .A(n445), .B(n444), .ZN(n528) );
  NAND2_X1 U495 ( .A1(n446), .A2(n528), .ZN(n561) );
  NOR2_X1 U496 ( .A1(n574), .A2(n561), .ZN(n449) );
  NOR2_X1 U497 ( .A1(n459), .A2(n528), .ZN(n450) );
  XNOR2_X1 U498 ( .A(n450), .B(KEYINPUT26), .ZN(n565) );
  XOR2_X1 U499 ( .A(n515), .B(KEYINPUT27), .Z(n457) );
  NAND2_X1 U500 ( .A1(n565), .A2(n457), .ZN(n454) );
  INV_X1 U501 ( .A(n528), .ZN(n518) );
  OR2_X1 U502 ( .A1(n518), .A2(n515), .ZN(n451) );
  NAND2_X1 U503 ( .A1(n459), .A2(n451), .ZN(n452) );
  XOR2_X1 U504 ( .A(KEYINPUT25), .B(n452), .Z(n453) );
  NAND2_X1 U505 ( .A1(n454), .A2(n453), .ZN(n455) );
  NAND2_X1 U506 ( .A1(n455), .A2(n511), .ZN(n456) );
  XNOR2_X1 U507 ( .A(n456), .B(KEYINPUT95), .ZN(n461) );
  INV_X1 U508 ( .A(n457), .ZN(n458) );
  NOR2_X1 U509 ( .A1(n511), .A2(n458), .ZN(n540) );
  XNOR2_X1 U510 ( .A(n459), .B(KEYINPUT28), .ZN(n521) );
  NAND2_X1 U511 ( .A1(n540), .A2(n521), .ZN(n526) );
  NOR2_X1 U512 ( .A1(n526), .A2(n528), .ZN(n460) );
  NOR2_X1 U513 ( .A1(n461), .A2(n460), .ZN(n478) );
  INV_X1 U514 ( .A(n574), .ZN(n549) );
  NAND2_X1 U515 ( .A1(n560), .A2(n549), .ZN(n462) );
  XNOR2_X1 U516 ( .A(KEYINPUT16), .B(n462), .ZN(n463) );
  NOR2_X1 U517 ( .A1(n478), .A2(n463), .ZN(n496) );
  INV_X1 U518 ( .A(n567), .ZN(n542) );
  AND2_X1 U519 ( .A1(n571), .A2(n542), .ZN(n464) );
  XNOR2_X1 U520 ( .A(n464), .B(KEYINPUT76), .ZN(n481) );
  NAND2_X1 U521 ( .A1(n496), .A2(n481), .ZN(n475) );
  NOR2_X1 U522 ( .A1(n511), .A2(n475), .ZN(n466) );
  XNOR2_X1 U523 ( .A(KEYINPUT34), .B(KEYINPUT96), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U525 ( .A(G1GAT), .B(n467), .Z(G1324GAT) );
  NOR2_X1 U526 ( .A1(n515), .A2(n475), .ZN(n469) );
  XNOR2_X1 U527 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U529 ( .A(G8GAT), .B(n470), .ZN(G1325GAT) );
  NOR2_X1 U530 ( .A1(n475), .A2(n518), .ZN(n474) );
  XOR2_X1 U531 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n472) );
  XNOR2_X1 U532 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n471) );
  XNOR2_X1 U533 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n474), .B(n473), .ZN(G1326GAT) );
  NOR2_X1 U535 ( .A1(n521), .A2(n475), .ZN(n477) );
  XNOR2_X1 U536 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(G1327GAT) );
  NOR2_X1 U538 ( .A1(n579), .A2(n478), .ZN(n479) );
  NAND2_X1 U539 ( .A1(n574), .A2(n479), .ZN(n480) );
  XNOR2_X1 U540 ( .A(KEYINPUT37), .B(n480), .ZN(n510) );
  NAND2_X1 U541 ( .A1(n510), .A2(n481), .ZN(n482) );
  XNOR2_X1 U542 ( .A(KEYINPUT38), .B(n482), .ZN(n492) );
  NOR2_X1 U543 ( .A1(n511), .A2(n492), .ZN(n486) );
  XOR2_X1 U544 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n484) );
  XNOR2_X1 U545 ( .A(G29GAT), .B(KEYINPUT102), .ZN(n483) );
  XNOR2_X1 U546 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(G1328GAT) );
  NOR2_X1 U548 ( .A1(n515), .A2(n492), .ZN(n487) );
  XOR2_X1 U549 ( .A(KEYINPUT104), .B(n487), .Z(n488) );
  XNOR2_X1 U550 ( .A(G36GAT), .B(n488), .ZN(G1329GAT) );
  NOR2_X1 U551 ( .A1(n492), .A2(n518), .ZN(n490) );
  XNOR2_X1 U552 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(n491), .ZN(G1330GAT) );
  NOR2_X1 U555 ( .A1(n492), .A2(n521), .ZN(n493) );
  XOR2_X1 U556 ( .A(KEYINPUT106), .B(n493), .Z(n494) );
  XNOR2_X1 U557 ( .A(G50GAT), .B(n494), .ZN(G1331GAT) );
  NOR2_X1 U558 ( .A1(n542), .A2(n555), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n495), .B(KEYINPUT108), .ZN(n509) );
  NAND2_X1 U560 ( .A1(n496), .A2(n509), .ZN(n504) );
  NOR2_X1 U561 ( .A1(n511), .A2(n504), .ZN(n498) );
  XNOR2_X1 U562 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(n499), .ZN(G1332GAT) );
  NOR2_X1 U565 ( .A1(n515), .A2(n504), .ZN(n501) );
  XNOR2_X1 U566 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(G1333GAT) );
  NOR2_X1 U568 ( .A1(n518), .A2(n504), .ZN(n502) );
  XOR2_X1 U569 ( .A(KEYINPUT110), .B(n502), .Z(n503) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(n503), .ZN(G1334GAT) );
  NOR2_X1 U571 ( .A1(n504), .A2(n521), .ZN(n508) );
  XOR2_X1 U572 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n506) );
  XNOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT112), .ZN(n505) );
  XNOR2_X1 U574 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  NAND2_X1 U576 ( .A1(n510), .A2(n509), .ZN(n520) );
  NOR2_X1 U577 ( .A1(n511), .A2(n520), .ZN(n513) );
  XNOR2_X1 U578 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NOR2_X1 U581 ( .A1(n515), .A2(n520), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G92GAT), .B(KEYINPUT115), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(G1337GAT) );
  NOR2_X1 U584 ( .A1(n518), .A2(n520), .ZN(n519) );
  XOR2_X1 U585 ( .A(G99GAT), .B(n519), .Z(G1338GAT) );
  NOR2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n523) );
  XNOR2_X1 U587 ( .A(KEYINPUT44), .B(KEYINPUT116), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U589 ( .A(G106GAT), .B(n524), .Z(G1339GAT) );
  NOR2_X1 U590 ( .A1(n525), .A2(n526), .ZN(n527) );
  NAND2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n536) );
  NOR2_X1 U592 ( .A1(n567), .A2(n536), .ZN(n529) );
  XOR2_X1 U593 ( .A(G113GAT), .B(n529), .Z(G1340GAT) );
  NOR2_X1 U594 ( .A1(n555), .A2(n536), .ZN(n531) );
  XNOR2_X1 U595 ( .A(KEYINPUT118), .B(KEYINPUT49), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G120GAT), .B(n532), .ZN(G1341GAT) );
  NOR2_X1 U598 ( .A1(n574), .A2(n536), .ZN(n534) );
  XNOR2_X1 U599 ( .A(KEYINPUT119), .B(KEYINPUT50), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  NOR2_X1 U602 ( .A1(n560), .A2(n536), .ZN(n538) );
  XNOR2_X1 U603 ( .A(KEYINPUT120), .B(KEYINPUT51), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(n539), .ZN(G1343GAT) );
  NAND2_X1 U606 ( .A1(n540), .A2(n565), .ZN(n541) );
  NOR2_X1 U607 ( .A1(n525), .A2(n541), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n542), .A2(n548), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n543), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT53), .Z(n545) );
  INV_X1 U611 ( .A(n548), .ZN(n551) );
  OR2_X1 U612 ( .A1(n551), .A2(n555), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n547) );
  XOR2_X1 U614 ( .A(KEYINPUT121), .B(KEYINPUT52), .Z(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  NAND2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n550), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U619 ( .A(G162GAT), .B(n553), .Z(G1347GAT) );
  NOR2_X1 U620 ( .A1(n561), .A2(n567), .ZN(n554) );
  XOR2_X1 U621 ( .A(G169GAT), .B(n554), .Z(G1348GAT) );
  NOR2_X1 U622 ( .A1(n561), .A2(n555), .ZN(n559) );
  XOR2_X1 U623 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n557) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U628 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(n564), .ZN(G1351GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n578) );
  NOR2_X1 U632 ( .A1(n567), .A2(n578), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(n570), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n578), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n578), .ZN(n575) );
  XOR2_X1 U640 ( .A(G211GAT), .B(n575), .Z(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n577) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n581) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(n581), .B(n580), .Z(G1355GAT) );
endmodule

