//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G469), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT4), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G104), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n196));
  INV_X1    g010(.A(G104), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(KEYINPUT3), .A3(G104), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n195), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n193), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n195), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n194), .A2(KEYINPUT3), .A3(G104), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT3), .B1(new_n194), .B2(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G101), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XOR2_X1   g025(.A(KEYINPUT0), .B(G128), .Z(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(new_n209), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n206), .A2(new_n193), .A3(G101), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n208), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT79), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n197), .B2(G107), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT80), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(new_n194), .B2(G104), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n194), .A2(KEYINPUT79), .A3(G104), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n197), .A2(KEYINPUT80), .A3(G107), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n217), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G101), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G143), .ZN(new_n225));
  INV_X1    g039(.A(G143), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G146), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n225), .A2(new_n227), .A3(new_n228), .A4(G128), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(new_n225), .B2(KEYINPUT1), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n229), .B1(new_n231), .B2(new_n209), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n200), .A2(new_n201), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n223), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT10), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(KEYINPUT81), .A3(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n215), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G134), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(G137), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n240), .A2(KEYINPUT11), .B1(new_n238), .B2(G137), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT11), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT64), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n239), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT11), .A3(G134), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT65), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n248), .A2(new_n245), .A3(KEYINPUT11), .A4(G134), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(G131), .B1(new_n244), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n239), .ZN(new_n252));
  OAI22_X1  g066(.A1(KEYINPUT64), .A2(new_n242), .B1(new_n245), .B2(G134), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n240), .A2(KEYINPUT11), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G131), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n255), .A2(new_n256), .A3(new_n247), .A4(new_n249), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n251), .A2(new_n257), .A3(KEYINPUT68), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n234), .A2(new_n235), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT81), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT1), .B1(new_n226), .B2(G146), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT66), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT67), .B(G128), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT66), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n225), .A2(new_n269), .A3(KEYINPUT1), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n225), .A2(new_n227), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n229), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT82), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n223), .A2(new_n275), .A3(new_n233), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n275), .B1(new_n223), .B2(new_n233), .ZN(new_n277));
  OAI211_X1 g091(.A(KEYINPUT10), .B(new_n274), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n237), .A2(new_n262), .A3(new_n265), .A4(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G953), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G227), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(G140), .ZN(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT78), .B(G110), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n282), .B(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n251), .A2(new_n257), .A3(KEYINPUT68), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT68), .B1(new_n251), .B2(new_n257), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n272), .A2(new_n230), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n271), .A2(new_n272), .B1(new_n289), .B2(new_n228), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n223), .A2(new_n233), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n234), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT12), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(KEYINPUT12), .A3(new_n258), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n285), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n278), .A2(new_n265), .A3(new_n236), .A4(new_n215), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n288), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n284), .B1(new_n300), .B2(new_n279), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n192), .B(new_n189), .C1(new_n298), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT84), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n300), .A2(new_n279), .ZN(new_n304));
  OAI22_X1  g118(.A1(new_n304), .A2(new_n284), .B1(new_n285), .B2(new_n297), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT84), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n192), .A4(new_n189), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n284), .ZN(new_n309));
  INV_X1    g123(.A(new_n279), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n309), .B1(new_n297), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n300), .A2(new_n279), .A3(new_n284), .ZN(new_n312));
  AOI21_X1  g126(.A(G902), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT83), .B1(new_n313), .B2(new_n192), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT83), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT12), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n292), .A2(new_n234), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n262), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n295), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n284), .B1(new_n319), .B2(new_n279), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n300), .A2(new_n279), .A3(new_n284), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n315), .B(G469), .C1(new_n322), .C2(G902), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n314), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n191), .B1(new_n308), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G214), .B1(G237), .B2(G902), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n213), .A2(G125), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(new_n290), .B2(G125), .ZN(new_n328));
  INV_X1    g142(.A(G224), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(G953), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n328), .B(new_n331), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT2), .B(G113), .Z(new_n333));
  XNOR2_X1  g147(.A(G116), .B(G119), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n208), .A2(new_n335), .A3(new_n214), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT85), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G116), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n339), .A2(KEYINPUT5), .A3(G119), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n340), .B1(new_n334), .B2(KEYINPUT5), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n341), .A2(G113), .B1(new_n334), .B2(new_n333), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(new_n276), .B2(new_n277), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n208), .A2(KEYINPUT85), .A3(new_n335), .A4(new_n214), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n338), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT86), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XOR2_X1   g161(.A(G110), .B(G122), .Z(new_n348));
  NAND4_X1  g162(.A1(new_n338), .A2(new_n343), .A3(KEYINPUT86), .A4(new_n344), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OR2_X1    g166(.A1(new_n345), .A2(new_n348), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n351), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n332), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(G210), .B1(G237), .B2(G902), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n330), .A2(KEYINPUT87), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n331), .A2(KEYINPUT7), .ZN(new_n358));
  OR3_X1    g172(.A1(new_n328), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  XOR2_X1   g173(.A(new_n291), .B(new_n342), .Z(new_n360));
  XOR2_X1   g174(.A(new_n348), .B(KEYINPUT8), .Z(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT87), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n358), .B1(new_n328), .B2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n353), .A2(new_n359), .A3(new_n362), .A4(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n189), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n355), .A2(new_n356), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n356), .B1(new_n355), .B2(new_n367), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n326), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n325), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT22), .B(G137), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n280), .A2(G221), .A3(G234), .ZN(new_n373));
  XOR2_X1   g187(.A(new_n372), .B(new_n373), .Z(new_n374));
  AND2_X1   g188(.A1(new_n230), .A2(KEYINPUT67), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n230), .A2(KEYINPUT67), .ZN(new_n376));
  OAI211_X1 g190(.A(KEYINPUT23), .B(G119), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G119), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G128), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT23), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT73), .B1(new_n378), .B2(G128), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT73), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n230), .A3(G119), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G110), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n377), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT74), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n379), .B1(new_n268), .B2(new_n378), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT24), .B(G110), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n377), .A2(new_n384), .A3(KEYINPUT74), .A4(new_n385), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n388), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT75), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(G125), .A2(G140), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(G125), .A2(G140), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT16), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G125), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n400), .A2(KEYINPUT16), .A3(G140), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n402), .A3(G146), .ZN(new_n403));
  INV_X1    g217(.A(G140), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n396), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n224), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT76), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT76), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(new_n409), .A3(new_n224), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n388), .A2(KEYINPUT75), .A3(new_n391), .A4(new_n392), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n395), .A2(new_n403), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT16), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n414), .B1(new_n405), .B2(new_n396), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n224), .B1(new_n415), .B2(new_n401), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n403), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n377), .A2(new_n384), .ZN(new_n418));
  OAI221_X1 g232(.A(new_n417), .B1(new_n389), .B2(new_n390), .C1(new_n418), .C2(new_n385), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n374), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n413), .A2(new_n419), .A3(new_n374), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n189), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT77), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT25), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G217), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n427), .B1(G234), .B2(new_n189), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT77), .B1(new_n423), .B2(new_n425), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n413), .A2(new_n419), .A3(new_n374), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n430), .A2(new_n420), .A3(G902), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(KEYINPUT25), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n426), .B(new_n428), .C1(new_n429), .C2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n423), .B2(new_n428), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n260), .A2(new_n261), .A3(new_n213), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n245), .A2(G134), .ZN(new_n436));
  OAI21_X1  g250(.A(G131), .B1(new_n239), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n274), .A2(new_n257), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(KEYINPUT30), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT30), .ZN(new_n440));
  INV_X1    g254(.A(new_n438), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n258), .A2(new_n213), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(new_n443), .A3(new_n335), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n335), .B(KEYINPUT69), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n435), .A2(new_n438), .A3(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(G237), .A2(G953), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G210), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(new_n201), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n444), .A2(new_n446), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT31), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n444), .A2(KEYINPUT31), .A3(new_n446), .A4(new_n452), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT28), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n446), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n335), .B1(new_n441), .B2(new_n442), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n446), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n459), .B1(new_n461), .B2(new_n458), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n451), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT70), .B1(G472), .B2(G902), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NOR3_X1   g280(.A1(KEYINPUT70), .A2(G472), .A3(G902), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT32), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n455), .A2(new_n456), .B1(new_n462), .B2(new_n451), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT32), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n471), .A2(new_n472), .A3(new_n468), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n446), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n445), .B1(new_n435), .B2(new_n438), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT28), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n459), .A2(KEYINPUT71), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n452), .A2(KEYINPUT29), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT71), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n446), .A2(new_n480), .A3(new_n458), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n477), .A2(new_n478), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n189), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT72), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n444), .A2(new_n446), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT29), .B1(new_n485), .B2(new_n451), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n462), .B2(new_n451), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT72), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n482), .A2(new_n488), .A3(new_n189), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n484), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G472), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n434), .B1(new_n474), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT93), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n339), .A2(G122), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n493), .B1(new_n494), .B2(KEYINPUT14), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n339), .A2(G122), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(KEYINPUT14), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT14), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n498), .A2(new_n339), .A3(KEYINPUT93), .A4(G122), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n495), .A2(new_n496), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G107), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT94), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n496), .A2(new_n194), .A3(new_n494), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(KEYINPUT94), .A3(G107), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n226), .A2(G128), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(new_n268), .B2(new_n226), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G134), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n238), .B(new_n506), .C1(new_n268), .C2(new_n226), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n503), .A2(new_n504), .A3(new_n505), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT95), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n501), .A2(new_n502), .B1(new_n508), .B2(new_n509), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT95), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n504), .A4(new_n505), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n496), .A2(new_n494), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G107), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n504), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT91), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT13), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n506), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n226), .A2(KEYINPUT13), .A3(G128), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n522), .B(new_n523), .C1(new_n268), .C2(new_n226), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G134), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT92), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT92), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(new_n527), .A3(G134), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n520), .A2(new_n509), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n188), .A2(G217), .A3(new_n280), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n516), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n530), .B1(new_n516), .B2(new_n529), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n189), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G478), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT96), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n539), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n189), .B(new_n541), .C1(new_n531), .C2(new_n532), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n447), .A2(G214), .ZN(new_n544));
  NAND2_X1  g358(.A1(KEYINPUT88), .A2(G143), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT88), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n226), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n447), .A2(new_n546), .A3(new_n226), .A4(G214), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n548), .A2(KEYINPUT17), .A3(G131), .A4(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(new_n416), .A3(new_n403), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT89), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n548), .A2(new_n549), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n256), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n548), .A2(G131), .A3(new_n549), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n550), .A2(new_n403), .A3(new_n416), .A4(KEYINPUT89), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n553), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n406), .A2(new_n224), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n408), .B2(new_n410), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT18), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n557), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(KEYINPUT18), .A2(G131), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n554), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n563), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(G113), .B(G122), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(new_n197), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n560), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n571), .ZN(new_n573));
  INV_X1    g387(.A(new_n568), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n574), .A2(new_n562), .A3(new_n565), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT19), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n406), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n405), .A2(KEYINPUT19), .A3(new_n396), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n224), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n403), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n557), .B2(new_n555), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n573), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n572), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(G475), .A2(G902), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT90), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT20), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT20), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n583), .A2(new_n588), .A3(new_n585), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G475), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n560), .A2(new_n569), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(new_n571), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(G902), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n590), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(G234), .A2(G237), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(G952), .A3(new_n280), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT97), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT21), .B(G898), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n596), .A2(G902), .A3(G953), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n598), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(new_n602), .B(KEYINPUT98), .Z(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n543), .A2(new_n595), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n371), .A2(new_n492), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT99), .B(G101), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G3));
  INV_X1    g422(.A(new_n326), .ZN(new_n609));
  INV_X1    g423(.A(new_n356), .ZN(new_n610));
  INV_X1    g424(.A(new_n332), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n350), .A2(new_n353), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT6), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n350), .A2(new_n351), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n610), .B1(new_n615), .B2(new_n366), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n355), .A2(new_n356), .A3(new_n367), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n609), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n303), .A2(new_n307), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n314), .A3(new_n323), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(new_n191), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n464), .A2(KEYINPUT100), .A3(new_n189), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n471), .B2(G902), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(new_n624), .A3(G472), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n423), .A2(new_n428), .ZN(new_n626));
  INV_X1    g440(.A(new_n428), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n424), .B1(new_n431), .B2(KEYINPUT25), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n423), .A2(new_n425), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n626), .B1(new_n630), .B2(new_n426), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n464), .A2(new_n469), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n625), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n621), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n534), .B(new_n189), .C1(new_n531), .C2(new_n532), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT33), .B1(new_n530), .B2(KEYINPUT101), .ZN(new_n637));
  OR3_X1    g451(.A1(new_n531), .A2(new_n532), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n637), .B1(new_n531), .B2(new_n532), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n636), .B1(new_n640), .B2(G478), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n534), .A2(new_n189), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n641), .A2(new_n595), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n604), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n634), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NOR2_X1   g462(.A1(new_n594), .A2(new_n591), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n589), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n589), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n587), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n543), .A2(new_n650), .A3(new_n603), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT103), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n634), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT35), .B(G107), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NAND4_X1  g473(.A1(new_n618), .A2(new_n605), .A3(new_n191), .A4(new_n620), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n625), .A2(new_n632), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n413), .A2(new_n419), .ZN(new_n662));
  INV_X1    g476(.A(new_n374), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(KEYINPUT36), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT104), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n662), .B(new_n665), .Z(new_n666));
  NOR2_X1   g480(.A1(new_n428), .A2(G902), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n630), .A2(new_n426), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n660), .A2(new_n661), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT37), .B(G110), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G12));
  AOI21_X1  g485(.A(new_n668), .B1(new_n474), .B2(new_n491), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n371), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n543), .A2(new_n650), .A3(new_n654), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n598), .B(KEYINPUT105), .ZN(new_n676));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n676), .B1(new_n677), .B2(new_n601), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT106), .B(G128), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G30));
  XOR2_X1   g496(.A(new_n678), .B(KEYINPUT39), .Z(new_n683));
  NAND3_X1  g497(.A1(new_n620), .A2(new_n191), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n684), .B(KEYINPUT108), .Z(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(KEYINPUT40), .Z(new_n686));
  NAND2_X1  g500(.A1(new_n616), .A2(new_n617), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT38), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n543), .A2(new_n595), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n464), .A2(KEYINPUT32), .A3(new_n469), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n472), .B1(new_n471), .B2(new_n468), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n475), .A2(new_n476), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n189), .B1(new_n692), .B2(new_n452), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n451), .B1(new_n444), .B2(new_n446), .ZN(new_n694));
  OAI21_X1  g508(.A(G472), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n690), .A2(new_n691), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT107), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n697), .A2(new_n326), .A3(new_n668), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n686), .A2(new_n688), .A3(new_n689), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G143), .ZN(G45));
  NOR2_X1   g514(.A1(new_n644), .A2(new_n678), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n674), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  NAND2_X1  g517(.A1(new_n305), .A2(new_n189), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n619), .A2(new_n191), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n370), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n492), .A2(new_n645), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT41), .B(G113), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G15));
  NAND3_X1  g524(.A1(new_n492), .A2(new_n656), .A3(new_n707), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  NAND2_X1  g526(.A1(new_n474), .A2(new_n491), .ZN(new_n713));
  INV_X1    g527(.A(new_n668), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n707), .A2(new_n713), .A3(new_n605), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  OAI21_X1  g530(.A(G472), .B1(new_n471), .B2(G902), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n477), .A2(new_n478), .A3(new_n481), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n455), .A2(new_n456), .B1(new_n718), .B2(new_n451), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n468), .B(KEYINPUT109), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n717), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n434), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n543), .A2(new_n595), .ZN(new_n723));
  AOI211_X1 g537(.A(new_n609), .B(new_n723), .C1(new_n616), .C2(new_n617), .ZN(new_n724));
  INV_X1    g538(.A(new_n706), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n722), .A2(new_n724), .A3(new_n603), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  NOR2_X1   g541(.A1(new_n668), .A2(new_n721), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n707), .A2(new_n728), .A3(new_n701), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  OR2_X1    g544(.A1(new_n690), .A2(KEYINPUT112), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n690), .A2(KEYINPUT112), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n731), .A2(new_n691), .A3(new_n491), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n631), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n616), .A2(new_n326), .A3(new_n617), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n735), .A2(new_n644), .A3(new_n678), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  OAI21_X1  g552(.A(G469), .B1(new_n322), .B2(G902), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT110), .B1(new_n619), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n619), .A2(KEYINPUT110), .A3(new_n739), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n191), .A3(new_n742), .ZN(new_n743));
  NOR4_X1   g557(.A1(new_n734), .A2(new_n737), .A3(new_n738), .A4(new_n743), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n619), .A2(KEYINPUT110), .A3(new_n739), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n745), .A2(new_n740), .A3(new_n190), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n368), .A2(new_n369), .A3(new_n609), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n746), .A2(new_n492), .A3(new_n701), .A4(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT111), .B1(new_n748), .B2(new_n738), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(KEYINPUT111), .A3(new_n738), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n744), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n256), .ZN(G33));
  INV_X1    g567(.A(G472), .ZN(new_n754));
  INV_X1    g568(.A(new_n489), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n488), .B1(new_n482), .B2(new_n189), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n754), .B1(new_n757), .B2(new_n487), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n690), .A2(new_n691), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n747), .B(new_n631), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n743), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT113), .B1(new_n761), .B2(new_n679), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n746), .A2(new_n492), .A3(new_n679), .A4(new_n747), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n238), .ZN(G36));
  XOR2_X1   g581(.A(new_n322), .B(KEYINPUT45), .Z(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(G469), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT114), .ZN(new_n770));
  NAND2_X1  g584(.A1(G469), .A2(G902), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n619), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n772), .A2(new_n773), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n191), .B(new_n683), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n595), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n641), .A2(new_n779), .A3(new_n643), .ZN(new_n780));
  XOR2_X1   g594(.A(new_n780), .B(KEYINPUT43), .Z(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n661), .A3(new_n714), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n735), .B1(new_n783), .B2(KEYINPUT44), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n778), .B(new_n784), .C1(KEYINPUT44), .C2(new_n783), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G137), .ZN(G39));
  OAI21_X1  g600(.A(new_n191), .B1(new_n775), .B2(new_n776), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT47), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g603(.A(KEYINPUT47), .B(new_n191), .C1(new_n775), .C2(new_n776), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n713), .A2(new_n631), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n736), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  AND3_X1   g608(.A1(new_n781), .A2(new_n676), .A3(new_n722), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n619), .A2(new_n705), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n191), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n747), .B(new_n795), .C1(new_n791), .C2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n688), .A2(new_n326), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n795), .A2(new_n725), .A3(new_n799), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT50), .Z(new_n801));
  NOR2_X1   g615(.A1(new_n697), .A2(new_n434), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n735), .A2(new_n706), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n802), .A2(new_n598), .A3(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n804), .A2(new_n779), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n641), .A2(new_n643), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n781), .A2(new_n676), .A3(new_n803), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n805), .A2(new_n806), .B1(new_n728), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n798), .A2(new_n801), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  INV_X1    g627(.A(new_n734), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT48), .B1(new_n808), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(G952), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n815), .A2(new_n816), .A3(G953), .ZN(new_n817));
  INV_X1    g631(.A(new_n644), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n804), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n808), .A2(KEYINPUT48), .A3(new_n814), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n812), .A2(new_n813), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n795), .A2(new_n707), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n595), .A2(new_n604), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n543), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n621), .A2(new_n633), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT117), .B1(new_n669), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n825), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n634), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n830));
  INV_X1    g644(.A(new_n661), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n371), .A3(new_n605), .A4(new_n714), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n606), .A2(new_n827), .A3(new_n833), .A4(new_n646), .ZN(new_n834));
  INV_X1    g648(.A(new_n744), .ZN(new_n835));
  INV_X1    g649(.A(new_n751), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n835), .B1(new_n836), .B2(new_n749), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n325), .A2(new_n678), .A3(new_n735), .ZN(new_n838));
  INV_X1    g652(.A(new_n654), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n839), .A2(new_n543), .A3(new_n649), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n672), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n746), .A2(new_n728), .A3(new_n736), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n762), .B2(new_n765), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n711), .A2(new_n715), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n708), .A2(new_n726), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n708), .A2(new_n711), .A3(new_n715), .A4(new_n726), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT116), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n834), .A2(new_n837), .A3(new_n845), .A4(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n326), .B(new_n689), .C1(new_n368), .C2(new_n369), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n696), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n678), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n746), .A2(new_n855), .A3(new_n668), .A4(new_n856), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n371), .B(new_n672), .C1(new_n679), .C2(new_n701), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n729), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT52), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT52), .A4(new_n729), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n861), .A2(KEYINPUT118), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT118), .B1(new_n861), .B2(new_n862), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n853), .A2(new_n865), .A3(KEYINPUT53), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n861), .A2(new_n862), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n853), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n866), .B1(KEYINPUT53), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT54), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT53), .B1(new_n850), .B2(KEYINPUT119), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n844), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n850), .A2(KEYINPUT119), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n873), .A2(new_n837), .A3(new_n834), .A4(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT120), .B1(new_n876), .B2(new_n865), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(new_n853), .B2(new_n868), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n867), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n861), .A2(KEYINPUT118), .A3(new_n862), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n827), .A2(new_n833), .A3(new_n606), .A4(new_n646), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n752), .A2(new_n885), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n844), .A2(new_n874), .A3(new_n872), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n883), .A2(new_n884), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n877), .A2(new_n879), .A3(new_n888), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n889), .A2(KEYINPUT54), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n822), .A2(new_n823), .A3(new_n871), .A4(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(G952), .B2(G953), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n802), .A2(new_n326), .A3(new_n191), .ZN(new_n893));
  INV_X1    g707(.A(new_n796), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT49), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n780), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(new_n895), .B2(new_n894), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n893), .A2(new_n897), .A3(new_n688), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT115), .Z(new_n899));
  NAND2_X1  g713(.A1(new_n892), .A2(new_n899), .ZN(G75));
  NAND2_X1  g714(.A1(new_n889), .A2(G902), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT56), .B1(new_n902), .B2(G210), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n352), .A2(new_n354), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(new_n332), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n903), .A2(new_n906), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n280), .A2(G952), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(G51));
  NAND2_X1  g724(.A1(new_n889), .A2(KEYINPUT54), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT121), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n889), .A2(new_n913), .A3(KEYINPUT54), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n912), .A2(new_n890), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n771), .B(KEYINPUT57), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n305), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n901), .A2(new_n770), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n909), .B1(new_n918), .B2(new_n919), .ZN(G54));
  INV_X1    g734(.A(new_n909), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n923));
  INV_X1    g737(.A(new_n583), .ZN(new_n924));
  OR3_X1    g738(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n922), .A2(new_n924), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n923), .B1(new_n922), .B2(new_n924), .ZN(new_n927));
  AND4_X1   g741(.A1(new_n921), .A2(new_n925), .A3(new_n926), .A4(new_n927), .ZN(G60));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n929));
  INV_X1    g743(.A(new_n640), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n642), .B(KEYINPUT59), .Z(new_n931));
  AND2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n915), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n929), .B1(new_n933), .B2(new_n921), .ZN(new_n934));
  AOI211_X1 g748(.A(KEYINPUT123), .B(new_n909), .C1(new_n915), .C2(new_n932), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n871), .A2(new_n890), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n930), .B1(new_n936), .B2(new_n931), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(G63));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT60), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n889), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n420), .B2(new_n430), .ZN(new_n942));
  INV_X1    g756(.A(new_n666), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n942), .B(new_n921), .C1(new_n943), .C2(new_n941), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g759(.A(G953), .B1(new_n599), .B2(new_n329), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n885), .B1(new_n851), .B2(new_n849), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(G953), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n904), .B1(G898), .B2(new_n280), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G69));
  NAND2_X1  g764(.A1(new_n439), .A2(new_n443), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n577), .A2(new_n578), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n793), .A2(new_n785), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n818), .B1(new_n543), .B2(new_n779), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT124), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n685), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n760), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n957), .B(new_n958), .C1(new_n956), .C2(new_n955), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n858), .A2(new_n729), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT62), .B1(new_n699), .B2(new_n960), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n699), .A2(KEYINPUT62), .A3(new_n960), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n954), .B(new_n959), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n953), .B1(new_n964), .B2(G953), .ZN(new_n965));
  INV_X1    g779(.A(new_n953), .ZN(new_n966));
  NAND2_X1  g780(.A1(G900), .A2(G953), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n778), .A2(new_n724), .A3(new_n814), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n752), .A2(new_n766), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n954), .A2(new_n960), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n966), .B(new_n967), .C1(new_n970), .C2(G953), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n965), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n280), .B1(G227), .B2(G900), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n971), .B2(KEYINPUT125), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n965), .B(new_n971), .C1(KEYINPUT125), .C2(new_n973), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(G72));
  INV_X1    g791(.A(new_n694), .ZN(new_n978));
  XNOR2_X1  g792(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n754), .A2(new_n189), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n979), .B(new_n980), .Z(new_n981));
  NAND3_X1  g795(.A1(new_n444), .A2(new_n446), .A3(new_n451), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n870), .A2(new_n978), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT127), .Z(new_n984));
  INV_X1    g798(.A(new_n981), .ZN(new_n985));
  INV_X1    g799(.A(new_n970), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(new_n947), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n921), .B1(new_n987), .B2(new_n982), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n964), .A2(new_n947), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n978), .B1(new_n989), .B2(new_n981), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n984), .A2(new_n988), .A3(new_n990), .ZN(G57));
endmodule


