//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT76), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  INV_X1    g004(.A(G227), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G953), .ZN(new_n192));
  XOR2_X1   g006(.A(new_n190), .B(new_n192), .Z(new_n193));
  XOR2_X1   g007(.A(new_n193), .B(KEYINPUT77), .Z(new_n194));
  INV_X1    g008(.A(KEYINPUT79), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT64), .A2(G146), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT64), .A2(G146), .ZN(new_n197));
  OAI21_X1  g011(.A(G143), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n198), .A2(new_n201), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT1), .B1(new_n205), .B2(G146), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n198), .A2(new_n201), .B1(G128), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT78), .A2(G107), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT78), .A2(G107), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n209), .B(G104), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  INV_X1    g027(.A(G104), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT3), .ZN(new_n215));
  OAI21_X1  g029(.A(G107), .B1(new_n214), .B2(KEYINPUT3), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n212), .A2(new_n213), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n214), .B1(new_n210), .B2(new_n211), .ZN(new_n218));
  NAND2_X1  g032(.A1(G104), .A2(G107), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(G101), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n195), .B1(new_n208), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n198), .A2(new_n201), .A3(new_n203), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT64), .B(G146), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n200), .B1(new_n224), .B2(G143), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n206), .A2(G128), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n223), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n227), .A2(KEYINPUT79), .A3(new_n217), .A4(new_n220), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  OR2_X1    g043(.A1(KEYINPUT64), .A2(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT64), .A2(G146), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n205), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT1), .ZN(new_n233));
  OAI21_X1  g047(.A(G128), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n205), .A2(G146), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n224), .B2(G143), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n234), .A2(new_n237), .B1(new_n225), .B2(new_n203), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n221), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n229), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT11), .ZN(new_n241));
  INV_X1    g055(.A(G134), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(G137), .ZN(new_n243));
  INV_X1    g057(.A(G137), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT11), .A3(G134), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(G137), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G131), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n243), .A2(new_n245), .A3(new_n249), .A4(new_n246), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n240), .A2(KEYINPUT12), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT12), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n222), .A2(new_n228), .B1(new_n238), .B2(new_n221), .ZN(new_n254));
  INV_X1    g068(.A(new_n251), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT10), .B1(new_n222), .B2(new_n228), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n209), .A2(G104), .ZN(new_n260));
  INV_X1    g074(.A(new_n211), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT78), .A2(G107), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n216), .A2(new_n215), .ZN(new_n264));
  OAI21_X1  g078(.A(G101), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n217), .A3(KEYINPUT4), .ZN(new_n266));
  AND2_X1   g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n237), .A2(new_n269), .B1(new_n225), .B2(new_n267), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n271), .B(G101), .C1(new_n263), .C2(new_n264), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n266), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT10), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n238), .A2(new_n275), .A3(new_n221), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n259), .A2(new_n255), .A3(new_n274), .A4(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n194), .B1(new_n257), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n276), .B1(new_n229), .B2(new_n275), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n255), .B1(new_n280), .B2(new_n274), .ZN(new_n281));
  NOR4_X1   g095(.A1(new_n258), .A2(new_n251), .A3(new_n273), .A4(new_n276), .ZN(new_n282));
  INV_X1    g096(.A(new_n193), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT80), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n279), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT12), .B1(new_n240), .B2(new_n251), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n254), .A2(new_n253), .A3(new_n255), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n278), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n194), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n282), .A2(new_n283), .ZN(new_n292));
  INV_X1    g106(.A(new_n281), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT80), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G469), .B1(new_n286), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G469), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n283), .B1(new_n281), .B2(new_n282), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n278), .B(new_n193), .C1(new_n287), .C2(new_n288), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n299), .B1(new_n302), .B2(new_n297), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n189), .B1(new_n296), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G125), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n238), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n198), .A2(new_n201), .A3(new_n267), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n196), .A2(new_n197), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n235), .B1(new_n310), .B2(new_n205), .ZN(new_n311));
  INV_X1    g125(.A(new_n269), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G125), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT83), .B(G224), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n317), .A2(G953), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n315), .B(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(KEYINPUT82), .A2(KEYINPUT6), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n217), .A2(new_n220), .ZN(new_n321));
  INV_X1    g135(.A(G119), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G116), .ZN(new_n323));
  INV_X1    g137(.A(G116), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G119), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT2), .B(G113), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G116), .B(G119), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT5), .ZN(new_n330));
  INV_X1    g144(.A(G113), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n324), .A2(G119), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT5), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n321), .A2(KEYINPUT81), .A3(new_n328), .A4(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n327), .B(new_n329), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n266), .A2(new_n338), .A3(new_n272), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n217), .A2(new_n335), .A3(new_n328), .A4(new_n220), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT81), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n336), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  XOR2_X1   g157(.A(G110), .B(G122), .Z(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n344), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n336), .A2(new_n339), .A3(new_n346), .A4(new_n342), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n320), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n343), .A2(new_n344), .B1(KEYINPUT82), .B2(KEYINPUT6), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n319), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n318), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n308), .A2(KEYINPUT7), .A3(new_n314), .A4(new_n351), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n334), .A2(KEYINPUT85), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n334), .A2(KEYINPUT85), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n330), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n321), .B(new_n328), .C1(new_n354), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n335), .A2(new_n328), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n221), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT86), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n221), .A2(new_n358), .A3(KEYINPUT86), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n357), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  XOR2_X1   g177(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n364));
  XNOR2_X1  g178(.A(new_n344), .B(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT7), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n315), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n315), .A2(new_n318), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n353), .A2(new_n366), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n350), .A2(new_n298), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G210), .B1(G237), .B2(G902), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(KEYINPUT87), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n373), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n350), .A2(new_n298), .A3(new_n375), .A4(new_n370), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n306), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G113), .B(G122), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(new_n214), .ZN(new_n379));
  INV_X1    g193(.A(G140), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G125), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n307), .A2(G140), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT69), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n381), .A2(new_n382), .A3(new_n383), .A4(KEYINPUT16), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n381), .A2(new_n382), .A3(KEYINPUT16), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT69), .B1(new_n381), .B2(KEYINPUT16), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G146), .ZN(new_n388));
  NOR2_X1   g202(.A1(G237), .A2(G953), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(G143), .A3(G214), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(G143), .B1(new_n389), .B2(G214), .ZN(new_n392));
  OAI21_X1  g206(.A(G131), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n392), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n249), .A3(new_n390), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n381), .A2(new_n382), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n397), .A2(KEYINPUT19), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(KEYINPUT19), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n224), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n388), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(G146), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n397), .A2(new_n310), .A3(KEYINPUT71), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT71), .ZN(new_n404));
  XNOR2_X1  g218(.A(G125), .B(G140), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n224), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n402), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n394), .A2(KEYINPUT18), .A3(G131), .A4(new_n390), .ZN(new_n408));
  NAND2_X1  g222(.A1(KEYINPUT18), .A2(G131), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n391), .B2(new_n392), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n379), .B1(new_n401), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT88), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI211_X1 g229(.A(KEYINPUT88), .B(new_n379), .C1(new_n401), .C2(new_n412), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT17), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n393), .A2(new_n395), .A3(new_n417), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n199), .B(new_n384), .C1(new_n385), .C2(new_n386), .ZN(new_n419));
  OAI211_X1 g233(.A(KEYINPUT17), .B(G131), .C1(new_n391), .C2(new_n392), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n418), .A2(new_n388), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n421), .A2(new_n379), .A3(new_n412), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n415), .A2(new_n416), .A3(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(G475), .A2(G902), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT89), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT90), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n413), .A2(new_n414), .ZN(new_n427));
  INV_X1    g241(.A(new_n422), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n413), .A2(new_n414), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT90), .ZN(new_n431));
  INV_X1    g245(.A(new_n425), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n426), .A2(new_n433), .A3(KEYINPUT20), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n379), .B1(new_n421), .B2(new_n412), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n298), .B1(new_n422), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT91), .ZN(new_n437));
  OR2_X1    g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n437), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(G475), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n441));
  OAI211_X1 g255(.A(KEYINPUT90), .B(new_n441), .C1(new_n423), .C2(new_n425), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n434), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G122), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT14), .B1(new_n444), .B2(G116), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT14), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n324), .A3(G122), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(G116), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n445), .A2(new_n447), .A3(KEYINPUT92), .A4(new_n448), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n445), .A2(new_n448), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n449), .B(G107), .C1(new_n450), .C2(KEYINPUT92), .ZN(new_n451));
  XNOR2_X1  g265(.A(G128), .B(G143), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(new_n242), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n261), .A2(new_n262), .ZN(new_n454));
  XNOR2_X1  g268(.A(G116), .B(G122), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n451), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n205), .A2(G128), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n202), .A2(G143), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT13), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n460), .B(G134), .C1(KEYINPUT13), .C2(new_n458), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n452), .A2(new_n242), .ZN(new_n462));
  INV_X1    g276(.A(new_n456), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n454), .A2(new_n455), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n461), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n457), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G217), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n187), .A2(new_n467), .A3(G953), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n457), .A2(new_n465), .A3(new_n468), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(KEYINPUT93), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT93), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n466), .A2(new_n473), .A3(new_n469), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(new_n298), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G478), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n477));
  XOR2_X1   g291(.A(new_n475), .B(new_n477), .Z(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G953), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n480), .A2(G952), .ZN(new_n481));
  NAND2_X1  g295(.A1(G234), .A2(G237), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  XOR2_X1   g298(.A(KEYINPUT21), .B(G898), .Z(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n482), .A2(G902), .A3(G953), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n484), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n443), .A2(new_n479), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n304), .A2(KEYINPUT94), .A3(new_n377), .A4(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT94), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n434), .A2(new_n440), .A3(new_n442), .ZN(new_n493));
  INV_X1    g307(.A(new_n489), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n377), .A2(new_n478), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n189), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n285), .B1(new_n279), .B2(new_n284), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n291), .A2(new_n294), .A3(KEYINPUT80), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n297), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n300), .A2(new_n301), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n297), .A3(new_n298), .ZN(new_n501));
  INV_X1    g315(.A(new_n299), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n496), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n492), .B1(new_n495), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT75), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n467), .B1(G234), .B2(new_n298), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n480), .A2(G221), .A3(G234), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(G137), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT73), .B(KEYINPUT22), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT23), .B1(new_n202), .B2(G119), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n202), .A2(G119), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(KEYINPUT68), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT68), .ZN(new_n516));
  OAI211_X1 g330(.A(G119), .B(new_n202), .C1(new_n516), .C2(KEYINPUT23), .ZN(new_n517));
  INV_X1    g331(.A(G110), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT70), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XOR2_X1   g335(.A(KEYINPUT24), .B(G110), .Z(new_n522));
  XNOR2_X1  g336(.A(G119), .B(G128), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n515), .A2(new_n517), .A3(KEYINPUT70), .A4(new_n518), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n224), .A2(new_n405), .A3(new_n404), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT71), .B1(new_n397), .B2(new_n310), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n387), .A2(G146), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT72), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT72), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n526), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n388), .A2(new_n419), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n518), .B1(new_n515), .B2(new_n517), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n523), .B2(new_n522), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n512), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n526), .A2(new_n532), .A3(new_n529), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n532), .B1(new_n526), .B2(new_n529), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n538), .B(new_n512), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n298), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT25), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n547));
  INV_X1    g361(.A(new_n512), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n542), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(KEYINPUT25), .A3(new_n298), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n508), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n507), .A2(G902), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(KEYINPUT74), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n506), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT25), .B1(new_n550), .B2(new_n298), .ZN(new_n558));
  AOI211_X1 g372(.A(new_n545), .B(G902), .C1(new_n549), .C2(new_n542), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n507), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(KEYINPUT75), .A3(new_n555), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g376(.A(KEYINPUT66), .B(KEYINPUT27), .Z(new_n563));
  NAND2_X1  g377(.A1(new_n389), .A2(G210), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT26), .B(G101), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT30), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n568), .A2(KEYINPUT65), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(KEYINPUT65), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n255), .A2(new_n313), .ZN(new_n571));
  INV_X1    g385(.A(new_n246), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n242), .A2(G137), .ZN(new_n573));
  OAI21_X1  g387(.A(G131), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n250), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n233), .B1(new_n224), .B2(G143), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n237), .B1(new_n576), .B2(new_n202), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n575), .B1(new_n577), .B2(new_n223), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n270), .A2(new_n251), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n202), .B1(new_n198), .B2(KEYINPUT1), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n223), .B1(new_n581), .B2(new_n311), .ZN(new_n582));
  INV_X1    g396(.A(new_n575), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n580), .A2(new_n584), .A3(KEYINPUT65), .A4(new_n568), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n337), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n580), .A2(new_n584), .A3(new_n337), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n567), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT67), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT67), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n591), .B(new_n567), .C1(new_n586), .C2(new_n588), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n251), .A2(new_n270), .B1(new_n582), .B2(new_n583), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT28), .B1(new_n593), .B2(new_n337), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n338), .B1(new_n571), .B2(new_n578), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n587), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n596), .B2(KEYINPUT28), .ZN(new_n597));
  INV_X1    g411(.A(new_n567), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT29), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n590), .A2(new_n592), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n597), .A2(KEYINPUT29), .A3(new_n598), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n298), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT32), .ZN(new_n604));
  NOR4_X1   g418(.A1(new_n586), .A2(KEYINPUT31), .A3(new_n588), .A4(new_n567), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n586), .A2(new_n588), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n598), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT31), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n597), .B2(new_n598), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n605), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(G472), .A2(G902), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n604), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n609), .A2(new_n607), .ZN(new_n614));
  OAI211_X1 g428(.A(KEYINPUT32), .B(new_n611), .C1(new_n614), .C2(new_n605), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n603), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n562), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n491), .A2(new_n505), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  OAI21_X1  g433(.A(G472), .B1(new_n610), .B2(G902), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n611), .B1(new_n614), .B2(new_n605), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n304), .A2(new_n562), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT95), .B(KEYINPUT33), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n472), .A2(new_n474), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n471), .A2(KEYINPUT96), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT96), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n457), .A2(new_n465), .A3(new_n628), .A4(new_n468), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n627), .A2(new_n470), .A3(KEYINPUT33), .A4(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n626), .A2(new_n298), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(G478), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n475), .A2(G478), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT97), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n632), .A2(new_n636), .A3(new_n633), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n443), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n489), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n371), .A2(new_n372), .ZN(new_n641));
  INV_X1    g455(.A(new_n372), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n350), .A2(new_n298), .A3(new_n642), .A4(new_n370), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n641), .A2(new_n305), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n624), .A2(new_n640), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NAND4_X1  g462(.A1(new_n479), .A2(new_n440), .A3(new_n442), .A4(new_n434), .ZN(new_n649));
  OAI21_X1  g463(.A(KEYINPUT98), .B1(new_n649), .B2(new_n489), .ZN(new_n650));
  OR3_X1    g464(.A1(new_n649), .A2(KEYINPUT98), .A3(new_n489), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n624), .A2(new_n645), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NOR2_X1   g468(.A1(new_n512), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n547), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n554), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n560), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n491), .A2(new_n505), .A3(new_n623), .A4(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  INV_X1    g475(.A(new_n616), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n496), .B(new_n658), .C1(new_n499), .C2(new_n503), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n662), .A2(new_n663), .A3(new_n644), .ZN(new_n664));
  INV_X1    g478(.A(G900), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n488), .A2(KEYINPUT99), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n667), .B1(new_n487), .B2(G900), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n666), .A2(new_n483), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n649), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n664), .A2(KEYINPUT100), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n304), .A2(new_n616), .A3(new_n645), .A4(new_n658), .ZN(new_n674));
  INV_X1    g488(.A(new_n671), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT101), .B(G128), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G30));
  XOR2_X1   g493(.A(new_n669), .B(KEYINPUT39), .Z(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n304), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n683), .A2(new_n478), .A3(new_n493), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n615), .A2(new_n613), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n606), .A2(new_n567), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n298), .B1(new_n596), .B2(new_n598), .ZN(new_n687));
  OAI21_X1  g501(.A(G472), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n658), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n306), .B1(new_n682), .B2(KEYINPUT40), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n374), .A2(new_n376), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n693), .B(new_n694), .Z(new_n695));
  NAND4_X1  g509(.A1(new_n684), .A2(new_n691), .A3(new_n692), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G143), .ZN(G45));
  NAND2_X1  g511(.A1(new_n635), .A2(new_n637), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n698), .A2(new_n493), .A3(new_n670), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n664), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  NOR2_X1   g515(.A1(new_n302), .A2(new_n297), .ZN(new_n702));
  AOI211_X1 g516(.A(G469), .B(G902), .C1(new_n300), .C2(new_n301), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n645), .A2(new_n704), .A3(new_n496), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n617), .A2(new_n706), .A3(new_n640), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND4_X1  g523(.A1(new_n617), .A2(new_n706), .A3(new_n650), .A4(new_n651), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  NAND4_X1  g525(.A1(new_n706), .A2(new_n616), .A3(new_n490), .A4(new_n658), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  NOR2_X1   g527(.A1(new_n493), .A2(new_n478), .ZN(new_n714));
  XOR2_X1   g528(.A(new_n611), .B(KEYINPUT103), .Z(new_n715));
  OAI21_X1  g529(.A(new_n620), .B1(new_n610), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n560), .A2(new_n555), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n706), .A2(new_n494), .A3(new_n714), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G122), .ZN(G24));
  NAND3_X1  g534(.A1(new_n638), .A2(new_n443), .A3(new_n669), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n658), .B(new_n620), .C1(new_n610), .C2(new_n715), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n705), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n307), .ZN(G27));
  INV_X1    g538(.A(KEYINPUT42), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n189), .A2(new_n306), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n279), .A2(new_n284), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(G469), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n727), .B1(new_n303), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n562), .A2(new_n616), .A3(new_n693), .A4(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n725), .B1(new_n731), .B2(new_n721), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g548(.A(KEYINPUT104), .B(new_n725), .C1(new_n731), .C2(new_n721), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n717), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n616), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n730), .A2(new_n693), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(KEYINPUT42), .A3(new_n699), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  NAND3_X1  g557(.A1(new_n617), .A2(new_n671), .A3(new_n740), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G134), .ZN(G36));
  NAND2_X1  g559(.A1(new_n728), .A2(KEYINPUT45), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT105), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n497), .A2(new_n498), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n728), .A2(new_n750), .A3(KEYINPUT45), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n747), .A2(G469), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT106), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n299), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n703), .B1(new_n756), .B2(KEYINPUT46), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n752), .B(new_n753), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n502), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n496), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n680), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n693), .A2(new_n305), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n638), .A2(new_n493), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT107), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n766), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n769), .A2(new_n622), .A3(new_n658), .A4(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n771), .A2(new_n772), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n764), .A2(new_n765), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G137), .ZN(G39));
  NOR2_X1   g592(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n763), .A2(new_n780), .ZN(new_n781));
  XOR2_X1   g595(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n501), .B1(new_n759), .B2(new_n760), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n756), .A2(KEYINPUT46), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n496), .B(new_n783), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n765), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n787), .A2(new_n562), .A3(new_n616), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n781), .A2(new_n699), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  INV_X1    g604(.A(new_n704), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n726), .B1(new_n791), .B2(KEYINPUT49), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n766), .B(new_n792), .C1(KEYINPUT49), .C2(new_n791), .ZN(new_n793));
  INV_X1    g607(.A(new_n695), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n793), .A2(new_n737), .A3(new_n690), .A4(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n769), .A2(new_n770), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(new_n484), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n704), .A2(new_n496), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n787), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(KEYINPUT114), .A3(new_n739), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n800), .B2(new_n738), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(KEYINPUT48), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n481), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n704), .A2(new_n189), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n779), .B1(new_n762), .B2(new_n496), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n189), .B(new_n782), .C1(new_n757), .C2(new_n761), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n796), .A2(new_n484), .A3(new_n718), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n765), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n798), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n811), .A2(new_n306), .A3(new_n794), .A4(new_n813), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n814), .B(KEYINPUT50), .Z(new_n815));
  NAND4_X1  g629(.A1(new_n799), .A2(new_n562), .A3(new_n484), .A4(new_n690), .ZN(new_n816));
  OR3_X1    g630(.A1(new_n816), .A2(new_n443), .A3(new_n638), .ZN(new_n817));
  INV_X1    g631(.A(new_n658), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n716), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n801), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n812), .A2(new_n815), .A3(new_n817), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n806), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n723), .B1(new_n664), .B2(new_n699), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n670), .B(new_n658), .C1(new_n303), .C2(new_n729), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n644), .A2(new_n493), .A3(new_n478), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n825), .A2(new_n496), .A3(new_n689), .A4(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT100), .B1(new_n664), .B2(new_n671), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n674), .A2(new_n673), .A3(new_n675), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n824), .B(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT52), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n710), .A2(new_n712), .A3(new_n719), .A4(new_n707), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(new_n736), .B2(new_n741), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n649), .B1(new_n698), .B2(new_n493), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n834), .A2(new_n377), .A3(new_n494), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n624), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n659), .A2(new_n618), .A3(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n819), .A2(new_n699), .A3(new_n693), .A4(new_n730), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT110), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n740), .A2(KEYINPUT110), .A3(new_n699), .A4(new_n819), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n840), .A2(new_n744), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n493), .A2(new_n478), .A3(new_n669), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n787), .A2(new_n662), .A3(new_n663), .A4(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n837), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n677), .A2(new_n846), .A3(new_n824), .A4(new_n827), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n831), .A2(new_n833), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT54), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n189), .B1(new_n757), .B2(new_n761), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n786), .B1(new_n852), .B2(new_n779), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n787), .B1(new_n853), .B2(new_n807), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n854), .A2(new_n811), .B1(new_n819), .B2(new_n801), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(KEYINPUT51), .A3(new_n817), .A4(new_n815), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n848), .A2(new_n849), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT111), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n831), .A2(new_n845), .A3(new_n847), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT112), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n849), .B1(new_n833), .B2(new_n860), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n833), .A2(new_n860), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n859), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT111), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n848), .A2(new_n865), .A3(new_n849), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n858), .A2(new_n863), .A3(new_n864), .A4(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n823), .A2(new_n851), .A3(new_n856), .A4(new_n867), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n804), .A2(KEYINPUT48), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n811), .A2(new_n645), .A3(new_n813), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT113), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n816), .A2(new_n639), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n868), .A2(new_n870), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(G952), .A2(G953), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n795), .B1(new_n874), .B2(new_n875), .ZN(G75));
  AND3_X1   g690(.A1(new_n848), .A2(new_n865), .A3(new_n849), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n865), .B1(new_n848), .B2(new_n849), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n298), .B1(new_n879), .B2(new_n863), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT56), .B1(new_n880), .B2(G210), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n348), .A2(new_n349), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(new_n319), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT55), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n884), .B1(KEYINPUT115), .B2(KEYINPUT56), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n881), .A2(new_n886), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n480), .A2(G952), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(G51));
  XNOR2_X1  g704(.A(new_n299), .B(KEYINPUT57), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n864), .B1(new_n879), .B2(new_n863), .ZN(new_n892));
  INV_X1    g706(.A(new_n867), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n500), .B(KEYINPUT116), .Z(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(KEYINPUT117), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n898));
  INV_X1    g712(.A(new_n891), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n858), .A2(new_n863), .A3(new_n866), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT54), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n899), .B1(new_n901), .B2(new_n867), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n898), .B1(new_n902), .B2(new_n895), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n880), .A2(new_n755), .A3(new_n754), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n897), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n889), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(G54));
  NAND2_X1  g721(.A1(KEYINPUT58), .A2(G475), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT118), .Z(new_n909));
  NAND4_X1  g723(.A1(new_n900), .A2(G902), .A3(new_n430), .A4(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n910), .A2(new_n906), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n900), .A2(G902), .A3(new_n909), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n912), .A2(KEYINPUT119), .A3(new_n423), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT119), .B1(new_n912), .B2(new_n423), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT120), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT120), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n917), .B(new_n911), .C1(new_n913), .C2(new_n914), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(G60));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT59), .Z(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n851), .B2(new_n867), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n626), .A2(new_n630), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n906), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n923), .B(new_n921), .C1(new_n901), .C2(new_n867), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(G63));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT60), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n900), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n930), .A2(new_n542), .A3(new_n549), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n900), .A2(new_n656), .A3(new_n929), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n931), .A2(KEYINPUT61), .A3(new_n906), .A4(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT122), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n932), .A2(new_n934), .ZN(new_n936));
  AND4_X1   g750(.A1(new_n906), .A2(new_n935), .A3(new_n931), .A4(new_n936), .ZN(new_n937));
  XOR2_X1   g751(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n938));
  OAI21_X1  g752(.A(new_n933), .B1(new_n937), .B2(new_n938), .ZN(G66));
  OR2_X1    g753(.A1(new_n837), .A2(new_n832), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n480), .ZN(new_n941));
  OAI21_X1  g755(.A(G953), .B1(new_n486), .B2(new_n317), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n882), .B1(G898), .B2(new_n480), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  XOR2_X1   g759(.A(KEYINPUT123), .B(KEYINPUT124), .Z(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G69));
  NAND2_X1  g761(.A1(new_n579), .A2(new_n585), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n398), .A2(new_n399), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n480), .A2(G900), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT127), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n852), .A2(new_n681), .A3(new_n739), .A4(new_n826), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n677), .A2(new_n824), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n955), .A2(new_n742), .A3(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n957), .A2(new_n777), .A3(new_n789), .A4(new_n744), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n954), .B1(new_n958), .B2(new_n480), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n951), .B(new_n953), .C1(new_n959), .C2(new_n952), .ZN(new_n960));
  INV_X1    g774(.A(new_n682), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n961), .A2(new_n617), .A3(new_n765), .A4(new_n834), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n956), .A2(new_n696), .ZN(new_n963));
  XNOR2_X1  g777(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n777), .A2(new_n789), .A3(new_n962), .A4(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n963), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n968), .A2(new_n480), .A3(new_n950), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT126), .B1(new_n960), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(G953), .B1(new_n191), .B2(new_n665), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  AOI211_X1 g787(.A(KEYINPUT126), .B(new_n971), .C1(new_n960), .C2(new_n969), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(G72));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n958), .B2(new_n940), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n606), .A3(new_n567), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n590), .A2(new_n607), .A3(new_n592), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n850), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n979), .A2(new_n906), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n977), .B1(new_n968), .B2(new_n940), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n983), .B2(new_n686), .ZN(G57));
endmodule


