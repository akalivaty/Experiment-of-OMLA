//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  INV_X1    g0007(.A(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT1), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  AND2_X1   g0027(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n229));
  NOR3_X1   g0029(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT65), .Z(new_n232));
  AOI21_X1  g0032(.A(new_n207), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n212), .B(new_n219), .C1(new_n220), .C2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n233), .A2(new_n220), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT67), .Z(new_n236));
  NOR2_X1   g0036(.A1(new_n234), .A2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n250), .B(new_n251), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  AND2_X1   g0054(.A1(G1), .A2(G13), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G226), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n256), .A2(G1), .A3(G13), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n259), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n263), .B1(new_n271), .B2(new_n224), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G222), .A2(G1698), .ZN(new_n273));
  XOR2_X1   g0073(.A(KEYINPUT70), .B(G223), .Z(new_n274));
  AOI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(G1698), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n272), .B1(new_n275), .B2(new_n271), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n266), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G179), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n279), .B(KEYINPUT71), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n216), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n222), .A2(KEYINPUT8), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT8), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n217), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n287), .A2(new_n289), .B1(G150), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n203), .A2(G20), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n283), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n283), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n258), .A2(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G50), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n295), .A2(new_n297), .B1(G50), .B2(new_n294), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n299), .B1(new_n278), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n280), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g0102(.A(new_n302), .B(KEYINPUT72), .Z(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT3), .B(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n223), .A2(G1698), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n304), .B(new_n305), .C1(G226), .C2(G1698), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G97), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n263), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G238), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n261), .B1(new_n309), .B2(new_n264), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(KEYINPUT76), .A2(KEYINPUT13), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n311), .B(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G179), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT75), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n311), .A2(new_n315), .A3(KEYINPUT13), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n315), .A2(KEYINPUT13), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(KEYINPUT13), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n317), .B(new_n318), .C1(new_n308), .C2(new_n310), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(G169), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT14), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT14), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n316), .A2(new_n322), .A3(G169), .A4(new_n319), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n314), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G68), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n290), .A2(G50), .B1(G20), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n224), .B2(new_n288), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n327), .A2(new_n282), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(KEYINPUT11), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(KEYINPUT11), .ZN(new_n330));
  INV_X1    g0130(.A(new_n294), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n325), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT12), .ZN(new_n333));
  INV_X1    g0133(.A(new_n295), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(G68), .A3(new_n296), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n329), .A2(new_n330), .A3(new_n333), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n324), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(new_n313), .B2(G190), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n316), .A2(G200), .A3(new_n319), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT9), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n299), .B(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n278), .A2(G200), .ZN(new_n345));
  INV_X1    g0145(.A(G190), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n344), .B(new_n345), .C1(new_n346), .C2(new_n278), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT10), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n296), .A2(G77), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n295), .A2(new_n349), .B1(G77), .B2(new_n294), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n287), .B(KEYINPUT74), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n290), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT15), .B(G87), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n352), .B1(new_n217), .B2(new_n224), .C1(new_n288), .C2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n350), .B1(new_n354), .B2(new_n282), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G179), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n261), .B1(new_n225), .B2(new_n264), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G1698), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n304), .A2(G232), .A3(new_n360), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n361), .B(KEYINPUT73), .ZN(new_n362));
  INV_X1    g0162(.A(G107), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n304), .A2(new_n363), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n271), .A2(new_n309), .A3(new_n360), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n362), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n357), .B(new_n359), .C1(new_n366), .C2(new_n263), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n263), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n368), .A2(new_n358), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n356), .B(new_n367), .C1(new_n369), .C2(G169), .ZN(new_n370));
  OAI211_X1 g0170(.A(G190), .B(new_n359), .C1(new_n366), .C2(new_n263), .ZN(new_n371));
  INV_X1    g0171(.A(G200), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n355), .B(new_n371), .C1(new_n369), .C2(new_n372), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n303), .A2(new_n342), .A3(new_n348), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n287), .A2(new_n296), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT79), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n334), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n377), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n378), .A2(new_n380), .B1(new_n294), .B2(new_n287), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n222), .A2(new_n325), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n382), .A2(new_n201), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(G20), .B1(G159), .B2(new_n290), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n271), .A2(new_n217), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT7), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(G20), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n386), .A2(new_n387), .B1(new_n271), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT77), .B1(new_n389), .B2(new_n325), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n387), .B1(new_n304), .B2(G20), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n271), .A2(new_n388), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n325), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT77), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n385), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n283), .B1(new_n396), .B2(KEYINPUT16), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT78), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n268), .A2(new_n270), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n267), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n388), .ZN(new_n401));
  AOI21_X1  g0201(.A(G20), .B1(new_n268), .B2(new_n270), .ZN(new_n402));
  OAI22_X1  g0202(.A1(new_n399), .A2(new_n401), .B1(new_n402), .B2(KEYINPUT7), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n384), .B1(new_n404), .B2(new_n325), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n381), .B1(new_n397), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n262), .A2(G1698), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n304), .B(new_n409), .C1(G223), .C2(G1698), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G87), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n263), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n261), .B1(new_n223), .B2(new_n264), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(new_n300), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n412), .A2(new_n413), .A3(new_n357), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT18), .B1(new_n408), .B2(new_n417), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n389), .A2(KEYINPUT77), .A3(new_n325), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n393), .A2(new_n394), .ZN(new_n420));
  OAI211_X1 g0220(.A(KEYINPUT16), .B(new_n384), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(new_n407), .A3(new_n282), .ZN(new_n422));
  INV_X1    g0222(.A(new_n381), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n417), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT18), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n414), .A2(new_n372), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(G190), .B2(new_n414), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n408), .A2(KEYINPUT17), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n422), .A2(new_n428), .A3(new_n423), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n418), .A2(new_n426), .A3(new_n429), .A4(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n375), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n263), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n258), .A2(G45), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT5), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n437), .B1(new_n438), .B2(G41), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT81), .B1(new_n438), .B2(G41), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT81), .ZN(new_n441));
  INV_X1    g0241(.A(G41), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT5), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n436), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G270), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n439), .A2(new_n257), .A3(new_n444), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT84), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT84), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n446), .A2(new_n450), .A3(new_n447), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G264), .A2(G1698), .ZN(new_n452));
  INV_X1    g0252(.A(G257), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n452), .B1(new_n453), .B2(G1698), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n304), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G303), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(new_n304), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT85), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n263), .B1(new_n457), .B2(new_n458), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n449), .A2(new_n451), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  INV_X1    g0262(.A(G97), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n217), .C1(G33), .C2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G116), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G20), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n282), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT20), .ZN(new_n468));
  XNOR2_X1  g0268(.A(new_n467), .B(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n294), .A2(G116), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n258), .A2(G33), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n283), .A2(new_n294), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n470), .B1(new_n472), .B2(G116), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G169), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT21), .B1(new_n461), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n459), .A2(new_n460), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n446), .A2(new_n450), .A3(new_n447), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n450), .B1(new_n446), .B2(new_n447), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT21), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n480), .A2(new_n481), .A3(G169), .A4(new_n474), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(G200), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n469), .A2(new_n473), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n484), .B(new_n485), .C1(new_n346), .C2(new_n480), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n357), .B1(new_n469), .B2(new_n473), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n487), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n483), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n225), .A2(G1698), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(new_n268), .A3(new_n270), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n360), .A2(KEYINPUT4), .A3(G244), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G250), .A2(G1698), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n304), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n462), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT80), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n462), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n502), .B1(new_n492), .B2(new_n493), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(KEYINPUT80), .A3(new_n498), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n263), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n445), .A2(G257), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n447), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G190), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n403), .A2(G107), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n290), .A2(G77), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT6), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n463), .A2(new_n363), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G97), .A2(G107), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n363), .A2(KEYINPUT6), .A3(G97), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n512), .B1(new_n519), .B2(G20), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n283), .B1(new_n510), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n294), .A2(G97), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n472), .B2(G97), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(G200), .B1(new_n505), .B2(new_n507), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n509), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT82), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n506), .A2(new_n357), .A3(new_n447), .ZN(new_n529));
  OAI22_X1  g0329(.A1(new_n505), .A2(new_n529), .B1(new_n521), .B2(new_n524), .ZN(new_n530));
  AND4_X1   g0330(.A1(KEYINPUT80), .A2(new_n494), .A3(new_n462), .A4(new_n498), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT80), .B1(new_n503), .B2(new_n498), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n436), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n507), .ZN(new_n534));
  AOI21_X1  g0334(.A(G169), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n528), .B1(new_n530), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n506), .A2(new_n357), .A3(new_n447), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n388), .B(new_n400), .C1(new_n271), .C2(KEYINPUT78), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n363), .B1(new_n538), .B2(new_n391), .ZN(new_n539));
  XNOR2_X1  g0339(.A(G97), .B(G107), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n517), .B1(new_n540), .B2(new_n513), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n511), .B1(new_n541), .B2(new_n217), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n282), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n533), .A2(new_n537), .B1(new_n543), .B2(new_n523), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n300), .B1(new_n505), .B2(new_n507), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT82), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n527), .A2(new_n536), .A3(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n268), .A2(new_n270), .A3(new_n217), .A4(G87), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT22), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT22), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n304), .A2(new_n550), .A3(new_n217), .A4(G87), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT23), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n217), .B2(G107), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n363), .A2(KEYINPUT23), .A3(G20), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n267), .A2(new_n465), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n558), .B2(G20), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n552), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT24), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n552), .A2(KEYINPUT24), .A3(new_n560), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n564), .A3(new_n282), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n472), .A2(G107), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT86), .ZN(new_n567));
  OR3_X1    g0367(.A1(new_n294), .A2(KEYINPUT25), .A3(G107), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT25), .B1(new_n294), .B2(G107), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n283), .A2(new_n294), .A3(new_n471), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n568), .B(new_n569), .C1(new_n571), .C2(new_n363), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT86), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n565), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n445), .A2(G264), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n453), .A2(G1698), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(G250), .B2(G1698), .ZN(new_n578));
  INV_X1    g0378(.A(G294), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n578), .A2(new_n271), .B1(new_n267), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n436), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n576), .A2(new_n447), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n300), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n582), .A2(G179), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n575), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n217), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT83), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(KEYINPUT83), .A3(new_n217), .ZN(new_n591));
  INV_X1    g0391(.A(G87), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n463), .A3(new_n363), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n304), .A2(new_n217), .A3(G68), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT19), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n288), .B2(new_n463), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n598), .A2(new_n282), .B1(new_n331), .B2(new_n353), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n472), .A2(G87), .ZN(new_n600));
  INV_X1    g0400(.A(G45), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(G1), .ZN(new_n602));
  INV_X1    g0402(.A(G250), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n258), .B2(G45), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n257), .A2(new_n602), .B1(new_n263), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(G238), .A2(G1698), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n225), .B2(G1698), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n557), .B1(new_n607), .B2(new_n304), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n605), .B(G190), .C1(new_n608), .C2(new_n263), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n309), .A2(new_n360), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n225), .A2(G1698), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n268), .A2(new_n610), .A3(new_n270), .A4(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n263), .B1(new_n612), .B2(new_n558), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n263), .A2(G274), .A3(new_n602), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n604), .A2(new_n263), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(G200), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n599), .A2(new_n600), .A3(new_n609), .A4(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n595), .A2(new_n597), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n282), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n353), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n472), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n353), .A2(new_n331), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(G169), .B1(new_n613), .B2(new_n616), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n605), .B(G179), .C1(new_n608), .C2(new_n263), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n618), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n582), .A2(G200), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n576), .A2(new_n581), .A3(G190), .A4(new_n447), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n565), .A2(new_n574), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n586), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n490), .A2(new_n547), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n435), .A2(new_n636), .ZN(G372));
  INV_X1    g0437(.A(new_n340), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n337), .B1(new_n638), .B2(new_n370), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n429), .A2(new_n432), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n424), .A2(new_n425), .ZN(new_n642));
  AOI211_X1 g0442(.A(KEYINPUT18), .B(new_n417), .C1(new_n422), .C2(new_n423), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n348), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n646), .A2(new_n303), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT90), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n630), .B1(new_n536), .B2(new_n546), .ZN(new_n649));
  XOR2_X1   g0449(.A(KEYINPUT89), .B(KEYINPUT26), .Z(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT88), .B1(new_n530), .B2(new_n535), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n621), .A2(new_n624), .A3(new_n600), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n617), .A2(new_n609), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT87), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n628), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n626), .A2(new_n627), .A3(KEYINPUT87), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n655), .B1(new_n659), .B2(new_n625), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT88), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n544), .A2(new_n545), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n652), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n649), .A2(new_n651), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n626), .A2(new_n627), .A3(KEYINPUT87), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT87), .B1(new_n626), .B2(new_n627), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n625), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n648), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n663), .A2(new_n664), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n530), .A2(new_n535), .A3(new_n528), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT82), .B1(new_n544), .B2(new_n545), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n631), .B(new_n651), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n669), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT90), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n483), .A2(new_n488), .A3(new_n586), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n634), .A2(new_n618), .A3(new_n668), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(new_n547), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n670), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n647), .B1(new_n435), .B2(new_n681), .ZN(G369));
  NAND2_X1  g0482(.A1(new_n483), .A2(new_n488), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n258), .A2(new_n217), .A3(G13), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n485), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n683), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n489), .B2(new_n691), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n575), .A2(new_n689), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT91), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT91), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n697), .A2(new_n634), .A3(new_n586), .A4(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n586), .B2(new_n690), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n683), .A2(new_n690), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n699), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n586), .A2(new_n689), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n701), .A2(new_n705), .ZN(G399));
  NOR2_X1   g0506(.A1(new_n209), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n593), .A2(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n214), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT31), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n576), .A2(new_n581), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n627), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n461), .A2(new_n508), .A3(new_n714), .A4(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(new_n534), .A3(new_n533), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT30), .B1(new_n718), .B2(new_n480), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n582), .B(new_n357), .C1(new_n613), .C2(new_n616), .ZN(new_n721));
  OR3_X1    g0521(.A1(new_n461), .A2(new_n508), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n720), .A2(KEYINPUT92), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT92), .B1(new_n720), .B2(new_n722), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n713), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n726), .A2(new_n689), .B1(new_n636), .B2(KEYINPUT31), .ZN(new_n727));
  AOI211_X1 g0527(.A(new_n713), .B(new_n690), .C1(new_n720), .C2(new_n722), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT29), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n680), .A2(new_n731), .A3(new_n690), .ZN(new_n732));
  INV_X1    g0532(.A(new_n488), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n584), .B1(new_n300), .B2(new_n582), .ZN(new_n734));
  AOI221_X4 g0534(.A(new_n733), .B1(new_n734), .B2(new_n575), .C1(new_n476), .C2(new_n482), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n678), .A2(new_n527), .A3(new_n536), .A4(new_n546), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n649), .A2(new_n651), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n663), .A2(new_n664), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n668), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n737), .B1(new_n740), .B2(KEYINPUT93), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT93), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n742), .B(new_n668), .C1(new_n738), .C2(new_n739), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n689), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n732), .B1(new_n744), .B2(new_n731), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n730), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n712), .B1(new_n747), .B2(G1), .ZN(G364));
  NOR2_X1   g0548(.A1(new_n208), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n258), .B1(new_n749), .B2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n707), .A2(new_n751), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n693), .A2(G330), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n752), .B1(new_n753), .B2(new_n694), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G13), .A2(G33), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n216), .B1(G20), .B2(new_n300), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT95), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n252), .A2(new_n601), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n762), .A2(KEYINPUT94), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(KEYINPUT94), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n209), .A2(new_n304), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n601), .B2(new_n215), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n763), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n209), .A2(new_n271), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n769), .A2(G355), .B1(new_n465), .B2(new_n209), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n760), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(G20), .A2(G179), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT96), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n372), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(G200), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G50), .A2(new_n775), .B1(new_n776), .B2(G58), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n773), .A2(new_n346), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G200), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n777), .B1(new_n224), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT97), .ZN(new_n782));
  NOR4_X1   g0582(.A1(new_n217), .A2(new_n372), .A3(G179), .A4(G190), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n271), .B1(new_n783), .B2(G107), .ZN(new_n784));
  NOR4_X1   g0584(.A1(new_n217), .A2(new_n346), .A3(new_n372), .A4(G179), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n773), .A2(new_n346), .A3(G200), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n784), .B1(new_n786), .B2(new_n592), .C1(new_n787), .C2(new_n325), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n357), .A2(new_n372), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT98), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n790), .A2(new_n217), .A3(G190), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G159), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT99), .B(KEYINPUT32), .Z(new_n794));
  OR3_X1    g0594(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n792), .B2(new_n793), .ZN(new_n796));
  OAI21_X1  g0596(.A(G20), .B1(new_n790), .B2(new_n346), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n795), .B(new_n796), .C1(new_n463), .C2(new_n798), .ZN(new_n799));
  OR3_X1    g0599(.A1(new_n782), .A2(new_n788), .A3(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT100), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n785), .B(KEYINPUT101), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n775), .ZN(new_n805));
  INV_X1    g0605(.A(G326), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n804), .A2(new_n456), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n791), .A2(G329), .ZN(new_n808));
  INV_X1    g0608(.A(G283), .ZN(new_n809));
  INV_X1    g0609(.A(new_n783), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n808), .B(new_n271), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n807), .B(new_n811), .C1(G322), .C2(new_n776), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G294), .A2(new_n797), .B1(new_n779), .B2(G311), .ZN(new_n813));
  XOR2_X1   g0613(.A(KEYINPUT33), .B(G317), .Z(new_n814));
  OAI211_X1 g0614(.A(new_n812), .B(new_n813), .C1(new_n787), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n800), .A2(new_n801), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n802), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n771), .B1(new_n817), .B2(new_n758), .ZN(new_n818));
  INV_X1    g0618(.A(new_n757), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n693), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n754), .B1(new_n820), .B2(new_n752), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT102), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G396));
  INV_X1    g0623(.A(new_n730), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n370), .A2(new_n689), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n373), .B1(new_n355), .B2(new_n690), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(new_n826), .B2(new_n370), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n681), .B2(new_n689), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n374), .A2(new_n690), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n679), .B1(new_n675), .B2(KEYINPUT90), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n665), .A2(new_n648), .A3(new_n669), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n752), .B1(new_n824), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n824), .B2(new_n835), .ZN(new_n837));
  INV_X1    g0637(.A(new_n752), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n758), .A2(new_n755), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(new_n224), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n758), .ZN(new_n841));
  INV_X1    g0641(.A(new_n787), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n803), .A2(G107), .B1(G283), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n456), .B2(new_n805), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n791), .A2(G311), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n304), .B1(new_n783), .B2(G87), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n845), .B(new_n846), .C1(new_n463), .C2(new_n798), .ZN(new_n847));
  INV_X1    g0647(.A(new_n776), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n465), .A2(new_n780), .B1(new_n848), .B2(new_n579), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n844), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n798), .A2(new_n222), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n810), .A2(new_n325), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n271), .B(new_n852), .C1(new_n791), .C2(G132), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n202), .B2(new_n804), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G143), .A2(new_n776), .B1(new_n779), .B2(G159), .ZN(new_n855));
  INV_X1    g0655(.A(G137), .ZN(new_n856));
  INV_X1    g0656(.A(G150), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n855), .B1(new_n856), .B2(new_n805), .C1(new_n857), .C2(new_n787), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT34), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n851), .B(new_n854), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n850), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n840), .B1(new_n841), .B2(new_n862), .C1(new_n827), .C2(new_n756), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n837), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G384));
  OR2_X1    g0665(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n866), .A2(G116), .A3(new_n218), .A4(new_n867), .ZN(new_n868));
  XOR2_X1   g0668(.A(KEYINPUT103), .B(KEYINPUT36), .Z(new_n869));
  XNOR2_X1  g0669(.A(new_n868), .B(new_n869), .ZN(new_n870));
  OR3_X1    g0670(.A1(new_n214), .A2(new_n224), .A3(new_n382), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n202), .A2(G68), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n258), .B(G13), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n422), .A2(new_n428), .A3(new_n423), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n875), .A2(new_n424), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n422), .A2(new_n423), .ZN(new_n878));
  INV_X1    g0678(.A(new_n687), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n384), .B1(new_n419), .B2(new_n420), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n406), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n381), .B1(new_n397), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n430), .B1(new_n884), .B2(new_n687), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n417), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT37), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n884), .A2(new_n687), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n881), .A2(new_n887), .B1(new_n433), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(KEYINPUT106), .A3(KEYINPUT38), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n877), .B1(new_n876), .B2(new_n880), .ZN(new_n892));
  INV_X1    g0692(.A(new_n417), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n878), .A2(new_n893), .ZN(new_n894));
  AND4_X1   g0694(.A1(new_n877), .A2(new_n894), .A3(new_n880), .A4(new_n430), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n880), .B1(new_n640), .B2(new_n644), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n881), .A2(new_n887), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n433), .A2(new_n888), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT38), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT106), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n890), .B(new_n891), .C1(new_n900), .C2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n337), .A2(new_n689), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n901), .A2(new_n902), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(KEYINPUT39), .A3(new_n903), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n906), .A2(new_n907), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n645), .A2(new_n687), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n910), .A2(new_n903), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n336), .A2(new_n689), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n341), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n916), .B1(new_n337), .B2(new_n340), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n661), .B1(new_n544), .B2(new_n545), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n668), .A2(new_n618), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT26), .B1(new_n923), .B2(new_n662), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n630), .B(new_n650), .C1(new_n536), .C2(new_n546), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n668), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n737), .B1(new_n926), .B2(new_n648), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n830), .B1(new_n927), .B2(new_n676), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT104), .B1(new_n928), .B2(new_n825), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT104), .ZN(new_n930));
  INV_X1    g0730(.A(new_n825), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n834), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n920), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n915), .B1(new_n933), .B2(KEYINPUT105), .ZN(new_n934));
  INV_X1    g0734(.A(new_n920), .ZN(new_n935));
  AOI211_X1 g0735(.A(KEYINPUT104), .B(new_n825), .C1(new_n680), .C2(new_n831), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n930), .B1(new_n834), .B2(new_n931), .ZN(new_n937));
  OAI211_X1 g0737(.A(KEYINPUT105), .B(new_n935), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n914), .B1(new_n934), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT107), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT105), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n915), .A3(new_n938), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT107), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n945), .A2(new_n946), .A3(new_n914), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n941), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n745), .A2(new_n434), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n647), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n948), .B(new_n950), .Z(new_n951));
  NAND2_X1  g0751(.A1(new_n547), .A2(new_n635), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT31), .B1(new_n952), .B2(new_n489), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n720), .A2(new_n722), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT92), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT31), .B1(new_n956), .B2(new_n723), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n953), .B1(new_n957), .B2(new_n690), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n956), .A2(KEYINPUT31), .A3(new_n689), .A4(new_n723), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT40), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n903), .A2(new_n904), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT106), .B1(new_n889), .B2(KEYINPUT38), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n909), .B1(new_n896), .B2(new_n898), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n827), .B1(new_n918), .B2(new_n919), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n958), .B2(new_n959), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n961), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT40), .B1(new_n910), .B2(new_n903), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n969), .A2(new_n967), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n434), .B(new_n960), .C1(new_n968), .C2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n964), .A2(new_n904), .A3(new_n903), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(new_n967), .A3(new_n890), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n973), .A2(KEYINPUT40), .B1(new_n967), .B2(new_n969), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n958), .A2(new_n959), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n435), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n971), .A2(new_n976), .A3(G330), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n951), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n258), .B2(new_n749), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n951), .A2(new_n977), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n874), .B1(new_n979), .B2(new_n980), .ZN(G367));
  OAI221_X1 g0781(.A(new_n759), .B1(new_n210), .B2(new_n353), .C1(new_n766), .C2(new_n244), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n792), .A2(new_n856), .B1(new_n222), .B2(new_n786), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(G150), .B2(new_n776), .ZN(new_n984));
  AOI22_X1  g0784(.A1(G143), .A2(new_n775), .B1(new_n842), .B2(G159), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n271), .B1(new_n783), .B2(G77), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT111), .Z(new_n987));
  AOI22_X1  g0787(.A1(G68), .A2(new_n797), .B1(new_n779), .B2(G50), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n984), .A2(new_n985), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT46), .B1(new_n785), .B2(G116), .ZN(new_n990));
  INV_X1    g0790(.A(G317), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n271), .B1(new_n463), .B2(new_n810), .C1(new_n792), .C2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n803), .A2(KEYINPUT46), .A3(G116), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n809), .B2(new_n780), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n798), .A2(new_n363), .B1(new_n579), .B2(new_n787), .ZN(new_n995));
  OR4_X1    g0795(.A1(new_n990), .A2(new_n992), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G303), .A2(new_n776), .B1(new_n775), .B2(G311), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT110), .Z(new_n998));
  OAI21_X1  g0798(.A(new_n989), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT47), .Z(new_n1000));
  OAI211_X1 g0800(.A(new_n752), .B(new_n982), .C1(new_n1000), .C2(new_n841), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n653), .A2(new_n689), .ZN(new_n1002));
  OR3_X1    g0802(.A1(new_n668), .A2(KEYINPUT108), .A3(new_n1002), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n660), .A2(new_n1002), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT108), .B1(new_n668), .B2(new_n1002), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1006), .A2(new_n757), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1001), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n547), .B1(new_n525), .B2(new_n690), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n544), .A2(new_n545), .A3(new_n689), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n703), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT42), .Z(new_n1013));
  INV_X1    g0813(.A(new_n1011), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1014), .A2(new_n586), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n1015), .A2(new_n673), .A3(new_n672), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1013), .B1(new_n689), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT43), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1006), .A2(new_n1018), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1006), .A2(new_n1018), .ZN(new_n1020));
  AND3_X1   g0820(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1019), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n701), .A2(new_n1014), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1025), .A2(KEYINPUT109), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT109), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n700), .B1(new_n683), .B2(new_n690), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1031), .A2(new_n703), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(new_n694), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n705), .A2(new_n1011), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT44), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n705), .A2(new_n1011), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT45), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1036), .A2(new_n701), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n701), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n747), .A2(new_n1034), .A3(new_n1040), .A4(new_n1043), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1044), .A2(new_n747), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n707), .B(KEYINPUT41), .Z(new_n1046));
  OAI21_X1  g0846(.A(new_n750), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1008), .B1(new_n1030), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(G387));
  NAND2_X1  g0849(.A1(new_n747), .A2(new_n1034), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n746), .A2(new_n1033), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n707), .B(KEYINPUT114), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n700), .A2(new_n819), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n709), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n769), .A2(new_n1055), .B1(new_n363), .B2(new_n209), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n351), .A2(new_n202), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT50), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n601), .B1(new_n325), .B2(new_n224), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n1058), .A2(new_n1055), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n765), .B1(new_n241), .B2(new_n601), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1056), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n760), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n838), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT112), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n785), .A2(G77), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n271), .B1(new_n783), .B2(G97), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(new_n792), .C2(new_n857), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT113), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G50), .A2(new_n776), .B1(new_n779), .B2(G68), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n842), .A2(new_n287), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n622), .A2(new_n797), .B1(new_n775), .B2(G159), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n304), .B1(new_n783), .B2(G116), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n798), .A2(new_n809), .B1(new_n579), .B2(new_n786), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G322), .A2(new_n775), .B1(new_n842), .B2(G311), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(new_n456), .B2(new_n780), .C1(new_n991), .C2(new_n848), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT48), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT49), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1074), .B1(new_n806), .B2(new_n792), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1073), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1065), .B1(new_n1084), .B2(new_n758), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1034), .A2(new_n751), .B1(new_n1054), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1053), .A2(new_n1086), .ZN(G393));
  NAND3_X1  g0887(.A1(new_n1043), .A2(new_n751), .A3(new_n1040), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n766), .A2(new_n248), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n759), .B1(new_n210), .B2(new_n463), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n752), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G311), .A2(new_n776), .B1(new_n775), .B2(G317), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT52), .Z(new_n1093));
  OAI221_X1 g0893(.A(new_n271), .B1(new_n810), .B2(new_n363), .C1(new_n786), .C2(new_n809), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G322), .B2(new_n791), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n798), .A2(new_n465), .B1(new_n456), .B2(new_n787), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G294), .B2(new_n779), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1093), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n791), .A2(G143), .B1(G68), .B2(new_n785), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT115), .Z(new_n1100));
  OAI21_X1  g0900(.A(new_n304), .B1(new_n810), .B2(new_n592), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n797), .B2(G77), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n351), .A2(new_n779), .B1(new_n842), .B2(G50), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G150), .A2(new_n775), .B1(new_n776), .B2(G159), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT51), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1098), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1091), .B1(new_n1107), .B2(new_n758), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n1011), .B2(new_n819), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1088), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1043), .A2(new_n1040), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n746), .B2(new_n1033), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1112), .A2(new_n1044), .A3(new_n1052), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT116), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1112), .A2(new_n1044), .A3(KEYINPUT116), .A4(new_n1052), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1110), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(G390));
  INV_X1    g0918(.A(new_n966), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n960), .A2(G330), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT117), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n960), .A2(new_n1119), .A3(KEYINPUT117), .A4(G330), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n907), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n942), .A2(new_n1125), .B1(new_n911), .B2(new_n906), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n826), .A2(new_n370), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n825), .B1(new_n744), .B2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n965), .B(new_n1125), .C1(new_n1128), .C2(new_n920), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1124), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n906), .A2(new_n911), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n933), .B2(new_n907), .ZN(new_n1133));
  OAI211_X1 g0933(.A(G330), .B(new_n827), .C1(new_n727), .C2(new_n728), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1134), .A2(new_n920), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1133), .A2(new_n1129), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1131), .A2(new_n751), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1132), .A2(new_n755), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n304), .B1(new_n810), .B2(new_n202), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n785), .A2(G150), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT53), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1139), .B(new_n1141), .C1(G125), .C2(new_n791), .ZN(new_n1142));
  INV_X1    g0942(.A(G132), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT54), .B(G143), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT119), .Z(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1142), .B1(new_n1143), .B2(new_n848), .C1(new_n780), .C2(new_n1146), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(G159), .A2(new_n797), .B1(new_n842), .B2(G137), .ZN(new_n1148));
  INV_X1    g0948(.A(G128), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1148), .B1(new_n1149), .B2(new_n805), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n803), .A2(G87), .B1(G107), .B2(new_n842), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n463), .B2(new_n780), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n304), .B(new_n852), .C1(new_n791), .C2(G294), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G116), .A2(new_n776), .B1(new_n775), .B2(G283), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1153), .B(new_n1154), .C1(new_n224), .C2(new_n798), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1147), .A2(new_n1150), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n758), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n839), .A2(new_n284), .A3(new_n286), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1138), .A2(new_n752), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1137), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(G330), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n975), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n434), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n949), .A2(new_n1164), .A3(new_n647), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1134), .A2(new_n920), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1122), .A2(new_n1166), .A3(new_n1123), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n929), .A2(new_n932), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n960), .A2(G330), .A3(new_n827), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n920), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1135), .A2(new_n1128), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1165), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1131), .A2(new_n1173), .A3(new_n1136), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1174), .A2(KEYINPUT118), .A3(new_n1052), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1173), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT118), .B1(new_n1174), .B2(new_n1052), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1161), .B1(new_n1179), .B2(new_n1180), .ZN(G378));
  INV_X1    g0981(.A(KEYINPUT57), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1165), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1182), .B1(new_n1174), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n912), .A2(new_n913), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n942), .A2(new_n943), .B1(new_n903), .B2(new_n910), .ZN(new_n1186));
  AOI211_X1 g0986(.A(KEYINPUT107), .B(new_n1185), .C1(new_n1186), .C2(new_n938), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n946), .B1(new_n945), .B2(new_n914), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n348), .A2(new_n302), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n299), .A2(new_n687), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT122), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n974), .B2(new_n1162), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1197), .B(G330), .C1(new_n968), .C2(new_n970), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1187), .A2(new_n1188), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n941), .B2(new_n947), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1184), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n1052), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1199), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n941), .A2(new_n947), .A3(new_n1201), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1174), .A2(new_n1183), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1204), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1193), .A2(new_n755), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n304), .A2(G41), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G50), .B(new_n1212), .C1(new_n267), .C2(new_n442), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G116), .A2(new_n775), .B1(new_n779), .B2(new_n622), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n463), .B2(new_n787), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n325), .A2(new_n798), .B1(new_n848), .B2(new_n363), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n792), .A2(new_n809), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1066), .B(new_n1212), .C1(new_n222), .C2(new_n810), .ZN(new_n1218));
  NOR4_X1   g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT120), .Z(new_n1220));
  INV_X1    g1020(.A(KEYINPUT58), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n776), .A2(G128), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n775), .A2(G125), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n1143), .B2(new_n787), .C1(new_n856), .C2(new_n780), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n786), .A2(new_n1146), .B1(new_n798), .B2(new_n857), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n267), .B(new_n442), .C1(new_n810), .C2(new_n793), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n791), .B2(G124), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT59), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1231), .B1(new_n1227), .B2(new_n1232), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1220), .A2(new_n1221), .B1(new_n1229), .B2(new_n1233), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1213), .B(new_n1234), .C1(new_n1221), .C2(new_n1220), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(new_n841), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT121), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n838), .B(new_n1237), .C1(new_n202), .C2(new_n839), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1207), .A2(new_n751), .B1(new_n1211), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1210), .A2(new_n1239), .ZN(G375));
  INV_X1    g1040(.A(new_n1046), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1169), .A2(new_n1165), .A3(new_n1172), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1177), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n750), .B(KEYINPUT123), .Z(new_n1245));
  NAND2_X1  g1045(.A1(new_n920), .A2(new_n755), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n1143), .A2(new_n805), .B1(new_n780), .B2(new_n857), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n304), .B1(new_n222), .B2(new_n810), .C1(new_n792), .C2(new_n1149), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(G159), .C2(new_n803), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1145), .A2(new_n842), .B1(new_n797), .B2(G50), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(new_n856), .C2(new_n848), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n304), .B1(new_n783), .B2(G77), .ZN(new_n1252));
  XOR2_X1   g1052(.A(new_n1252), .B(KEYINPUT124), .Z(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G97), .B2(new_n803), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G303), .A2(new_n791), .B1(new_n797), .B2(new_n622), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(G294), .A2(new_n775), .B1(new_n842), .B2(G116), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(G107), .A2(new_n779), .B1(new_n776), .B2(G283), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n841), .B1(new_n1251), .B2(new_n1258), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n838), .B(new_n1259), .C1(new_n325), .C2(new_n839), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1244), .A2(new_n1245), .B1(new_n1246), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1243), .A2(new_n1261), .ZN(G381));
  NAND3_X1  g1062(.A1(new_n1053), .A2(new_n822), .A3(new_n1086), .ZN(new_n1263));
  OR3_X1    g1063(.A1(G387), .A2(G384), .A3(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1117), .A2(new_n1261), .A3(new_n1243), .ZN(new_n1265));
  OR4_X1    g1065(.A1(G378), .A2(new_n1264), .A3(G375), .A4(new_n1265), .ZN(G407));
  AND2_X1   g1066(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1180), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1160), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n688), .A2(G213), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G407), .B(G213), .C1(G375), .C2(new_n1272), .ZN(G409));
  NAND2_X1  g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1263), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1117), .A2(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1117), .A2(new_n1275), .ZN(new_n1277));
  OAI21_X1  g1077(.A(G387), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1117), .A2(new_n1275), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1117), .A2(new_n1275), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(new_n1048), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G378), .B(new_n1239), .C1(new_n1204), .C2(new_n1209), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1241), .B(new_n1208), .C1(new_n1200), .C2(new_n1202), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1238), .A2(new_n1211), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1245), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1284), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1269), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1283), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1270), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT60), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1242), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1242), .A2(new_n1291), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1292), .A2(new_n1052), .A3(new_n1177), .A4(new_n1293), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1294), .A2(G384), .A3(new_n1261), .ZN(new_n1295));
  AOI21_X1  g1095(.A(G384), .B1(new_n1294), .B2(new_n1261), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1271), .A2(G2897), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1297), .B(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT61), .B1(new_n1290), .B2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1289), .A2(new_n1270), .A3(new_n1297), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(KEYINPUT62), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1302), .A2(KEYINPUT62), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1282), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT63), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1295), .A2(new_n1296), .A3(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1289), .A2(new_n1270), .A3(new_n1308), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1271), .B1(new_n1283), .B2(new_n1288), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT63), .B1(new_n1312), .B2(new_n1297), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT125), .B1(new_n1314), .B2(new_n1301), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1282), .B1(new_n1312), .B2(new_n1308), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1302), .A2(new_n1307), .ZN(new_n1317));
  AND4_X1   g1117(.A1(KEYINPUT125), .A2(new_n1301), .A3(new_n1316), .A4(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1306), .B1(new_n1315), .B2(new_n1318), .ZN(G405));
  AOI21_X1  g1119(.A(G378), .B1(new_n1210), .B2(new_n1239), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT126), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT127), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1283), .A2(KEYINPUT126), .ZN(new_n1324));
  OAI221_X1 g1124(.A(new_n1322), .B1(new_n1323), .B2(new_n1297), .C1(new_n1320), .C2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1297), .A2(new_n1323), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1282), .B(new_n1326), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1325), .B(new_n1327), .ZN(G402));
endmodule


