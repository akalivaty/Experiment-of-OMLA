//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1293, new_n1294, new_n1295, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT64), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n204), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT65), .B(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n209), .B(new_n214), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT2), .B(G226), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XNOR2_X1  g0034(.A(G50), .B(G68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G58), .B(G77), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  NAND3_X1  g0041(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(new_n212), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT3), .ZN(new_n245));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(new_n204), .A3(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT7), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT75), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n247), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n248), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n253), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT75), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(G107), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G107), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(KEYINPUT6), .A3(G97), .ZN(new_n259));
  INV_X1    g0059(.A(G97), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n258), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G97), .A2(G107), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n259), .B1(new_n263), .B2(KEYINPUT6), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n264), .A2(G20), .B1(G77), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n244), .B1(new_n257), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT67), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n242), .A2(new_n268), .A3(new_n212), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n268), .B1(new_n242), .B2(new_n212), .ZN(new_n270));
  INV_X1    g0070(.A(G13), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n271), .A2(new_n204), .A3(G1), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT81), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n203), .A2(G33), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n243), .A2(KEYINPUT67), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n271), .A2(G1), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G20), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n242), .A2(new_n268), .A3(new_n212), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n277), .A2(new_n279), .A3(new_n280), .A4(new_n275), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT81), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n260), .B1(new_n276), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n279), .A2(G97), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n267), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(G1), .A3(G13), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  AND2_X1   g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NOR2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  OAI211_X1 g0090(.A(G244), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT4), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G283), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n247), .A2(new_n248), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G250), .A2(G1698), .ZN(new_n297));
  NAND2_X1  g0097(.A1(KEYINPUT4), .A2(G244), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n297), .B1(new_n298), .B2(G1698), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n295), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n287), .B1(new_n293), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n203), .A2(G45), .ZN(new_n302));
  OR2_X1    g0102(.A1(KEYINPUT5), .A2(G41), .ZN(new_n303));
  NAND2_X1  g0103(.A1(KEYINPUT5), .A2(G41), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(G274), .A3(new_n287), .ZN(new_n306));
  INV_X1    g0106(.A(G45), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(G1), .ZN(new_n308));
  INV_X1    g0108(.A(new_n304), .ZN(new_n309));
  NOR2_X1   g0109(.A1(KEYINPUT5), .A2(G41), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(G257), .A3(new_n287), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n301), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(G169), .B2(new_n314), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n285), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT83), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n293), .A2(new_n300), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n303), .A2(new_n304), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n321), .B1(new_n308), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G274), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n324), .A2(G257), .B1(new_n326), .B2(new_n305), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G200), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT82), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n314), .B2(G190), .ZN(new_n331));
  INV_X1    g0131(.A(G190), .ZN(new_n332));
  NOR4_X1   g0132(.A1(new_n301), .A2(new_n313), .A3(KEYINPUT82), .A4(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n329), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n283), .A2(new_n284), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n257), .A2(new_n266), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n243), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n319), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G200), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n314), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n322), .A2(G190), .A3(new_n327), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT82), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n314), .A2(new_n330), .A3(G190), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n341), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n345), .A2(KEYINPUT83), .A3(new_n285), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n318), .B1(new_n339), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT80), .ZN(new_n348));
  OR3_X1    g0148(.A1(new_n204), .A2(KEYINPUT68), .A3(G1), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT68), .B1(new_n204), .B2(G1), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT8), .B(G58), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(new_n273), .B1(new_n272), .B2(new_n353), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n254), .A2(G68), .A3(new_n256), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT74), .B1(new_n265), .B2(G159), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n265), .A2(KEYINPUT74), .A3(G159), .ZN(new_n359));
  XNOR2_X1  g0159(.A(G58), .B(G68), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n358), .A2(new_n359), .B1(G20), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT16), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n289), .A2(new_n290), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT7), .B1(new_n363), .B2(new_n204), .ZN(new_n364));
  OAI21_X1  g0164(.A(G68), .B1(new_n364), .B2(new_n255), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(KEYINPUT16), .A3(new_n361), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n243), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n355), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(new_n287), .A3(G274), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n287), .A2(new_n369), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n227), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G87), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n246), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  OR2_X1    g0176(.A1(G223), .A2(G1698), .ZN(new_n377));
  INV_X1    g0177(.A(G226), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G1698), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n376), .B1(new_n380), .B2(new_n363), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT76), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n287), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(G223), .A2(G1698), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n378), .B2(G1698), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n375), .B1(new_n385), .B2(new_n296), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT76), .ZN(new_n387));
  AOI211_X1 g0187(.A(G190), .B(new_n373), .C1(new_n383), .C2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT78), .ZN(new_n389));
  INV_X1    g0189(.A(new_n373), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n321), .B1(new_n386), .B2(KEYINPUT76), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n381), .A2(new_n382), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n388), .A2(new_n389), .B1(new_n340), .B2(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n332), .B(new_n390), .C1(new_n391), .C2(new_n392), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT78), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n368), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n348), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n393), .A2(new_n340), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n383), .A2(new_n387), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n401), .A2(new_n389), .A3(new_n332), .A4(new_n390), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n396), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n355), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n356), .A2(new_n361), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n216), .B1(new_n251), .B2(new_n253), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n360), .A2(G20), .ZN(new_n409));
  INV_X1    g0209(.A(new_n359), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(new_n357), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n244), .B1(new_n412), .B2(KEYINPUT16), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n404), .B1(new_n407), .B2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n403), .A2(new_n414), .A3(new_n348), .A4(new_n398), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT79), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n403), .A2(new_n414), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n417), .B1(new_n418), .B2(KEYINPUT17), .ZN(new_n419));
  AOI211_X1 g0219(.A(KEYINPUT79), .B(new_n398), .C1(new_n403), .C2(new_n414), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n399), .A2(new_n416), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT77), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n401), .A2(new_n422), .A3(new_n315), .A4(new_n390), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n315), .B(new_n390), .C1(new_n391), .C2(new_n392), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT77), .ZN(new_n425));
  AOI21_X1  g0225(.A(G169), .B1(new_n401), .B2(new_n390), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n368), .ZN(new_n428));
  XOR2_X1   g0228(.A(new_n428), .B(KEYINPUT18), .Z(new_n429));
  NAND2_X1  g0229(.A1(new_n421), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT69), .ZN(new_n431));
  INV_X1    g0231(.A(new_n265), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n353), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n431), .B2(new_n432), .ZN(new_n434));
  INV_X1    g0234(.A(G77), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n434), .B1(new_n204), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT70), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n246), .A2(G20), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  XOR2_X1   g0239(.A(KEYINPUT15), .B(G87), .Z(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n436), .A2(new_n437), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n436), .A2(new_n437), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n243), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n352), .A2(new_n435), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n272), .A2(new_n243), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n445), .A2(new_n446), .B1(new_n435), .B2(new_n272), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n363), .A2(G1698), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n450), .A2(G232), .B1(G107), .B2(new_n363), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n363), .A2(new_n288), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n451), .B1(new_n215), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n321), .ZN(new_n455));
  INV_X1    g0255(.A(new_n371), .ZN(new_n456));
  INV_X1    g0256(.A(new_n372), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(G244), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G169), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(G179), .B2(new_n459), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n449), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n272), .A2(new_n216), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n464), .B(KEYINPUT12), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n277), .A2(new_n280), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n265), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n439), .B2(new_n435), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT11), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n446), .A2(new_n351), .A3(G68), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n465), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT11), .B1(new_n466), .B2(new_n468), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT14), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n227), .A2(G1698), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n296), .B(new_n476), .C1(G226), .C2(G1698), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G97), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT73), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n479), .B(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n321), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n456), .B1(G238), .B2(new_n457), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT13), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n482), .B2(new_n483), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n475), .B(G169), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n487), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(G179), .A3(new_n485), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n485), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n475), .B1(new_n492), .B2(G169), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n474), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(G200), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n495), .B(new_n473), .C1(new_n332), .C2(new_n492), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n455), .A2(G190), .A3(new_n458), .ZN(new_n497));
  XOR2_X1   g0297(.A(KEYINPUT71), .B(G200), .Z(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n459), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n444), .A2(new_n447), .A3(new_n497), .A4(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n463), .A2(new_n494), .A3(new_n496), .A4(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n456), .B1(G226), .B2(new_n457), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n450), .A2(G222), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n505), .B(KEYINPUT66), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n452), .A2(G223), .B1(G77), .B2(new_n363), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n504), .B1(new_n508), .B2(new_n321), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n499), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n273), .A2(G50), .A3(new_n351), .ZN(new_n512));
  INV_X1    g0312(.A(G150), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n353), .A2(new_n439), .B1(new_n513), .B2(new_n432), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G58), .A2(G68), .ZN(new_n515));
  INV_X1    g0315(.A(G50), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n204), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n466), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n512), .B(new_n518), .C1(G50), .C2(new_n279), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n519), .A2(KEYINPUT9), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(KEYINPUT9), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n509), .A2(G190), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n511), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT72), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT10), .ZN(new_n525));
  OR2_X1    g0325(.A1(new_n524), .A2(KEYINPUT10), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n511), .A2(new_n522), .A3(new_n524), .A4(KEYINPUT10), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n509), .A2(new_n315), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n529), .B(new_n519), .C1(G169), .C2(new_n509), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n430), .A2(new_n502), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n296), .A2(G257), .A3(G1698), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n296), .A2(G250), .A3(new_n288), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G294), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n321), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n324), .A2(G264), .B1(new_n326), .B2(new_n305), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G169), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n537), .A2(G179), .A3(new_n538), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT92), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT24), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT89), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n204), .B(G87), .C1(new_n289), .C2(new_n290), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT90), .ZN(new_n548));
  OR2_X1    g0348(.A1(new_n546), .A2(KEYINPUT22), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n548), .B1(new_n547), .B2(new_n549), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n546), .B(KEYINPUT22), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n547), .A2(new_n549), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT90), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n546), .A2(KEYINPUT22), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT91), .B1(new_n258), .B2(G20), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT23), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n561), .A2(new_n562), .B1(G116), .B2(new_n438), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n545), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n563), .ZN(new_n565));
  AOI211_X1 g0365(.A(KEYINPUT24), .B(new_n565), .C1(new_n552), .C2(new_n557), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n243), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n272), .A2(new_n258), .ZN(new_n568));
  XNOR2_X1  g0368(.A(new_n568), .B(KEYINPUT25), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n276), .A2(new_n282), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n569), .B1(new_n570), .B2(G107), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n544), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n539), .A2(new_n340), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(G190), .B2(new_n539), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n567), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n570), .A2(new_n440), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n440), .A2(new_n279), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT19), .B1(new_n438), .B2(G97), .ZN(new_n580));
  AOI21_X1  g0380(.A(G20), .B1(new_n247), .B2(new_n248), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n580), .B1(G68), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(G20), .B1(new_n481), .B2(KEYINPUT19), .ZN(new_n583));
  NOR3_X1   g0383(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n579), .B1(new_n585), .B2(new_n243), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n578), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(G250), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n307), .B2(G1), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n203), .A2(new_n325), .A3(G45), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n287), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT84), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n287), .A2(new_n589), .A3(new_n590), .A4(KEYINPUT84), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G116), .ZN(new_n596));
  INV_X1    g0396(.A(G244), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G1698), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(G238), .B2(G1698), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n596), .B1(new_n599), .B2(new_n363), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n321), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT85), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT85), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n595), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n315), .A3(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n595), .A2(new_n601), .A3(new_n604), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n604), .B1(new_n595), .B2(new_n601), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n460), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n587), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n498), .B1(new_n603), .B2(new_n605), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n603), .A2(G190), .A3(new_n605), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT87), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT87), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n603), .A2(new_n614), .A3(G190), .A4(new_n605), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n611), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n585), .A2(new_n243), .ZN(new_n617));
  INV_X1    g0417(.A(new_n579), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n274), .B1(new_n273), .B2(new_n275), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n281), .A2(KEYINPUT81), .ZN(new_n621));
  OAI21_X1  g0421(.A(G87), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT86), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT86), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n570), .A2(new_n624), .A3(G87), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n619), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n610), .B1(new_n616), .B2(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n294), .B(new_n204), .C1(G33), .C2(new_n260), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n204), .A2(G116), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n630), .A3(new_n243), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT20), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(G116), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n203), .B2(G33), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n446), .A2(new_n635), .B1(new_n278), .B2(new_n629), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n324), .A2(G270), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n306), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n637), .A2(G179), .A3(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(G264), .B(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n642));
  OAI211_X1 g0442(.A(G257), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n643));
  INV_X1    g0443(.A(G303), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n296), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n645), .A2(KEYINPUT88), .A3(new_n321), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT88), .B1(new_n645), .B2(new_n321), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT21), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n640), .B1(new_n647), .B2(new_n648), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n460), .B1(new_n633), .B2(new_n636), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n652), .A2(new_n651), .A3(new_n653), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n650), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n637), .B1(new_n652), .B2(G200), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n332), .B2(new_n652), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n627), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  AND4_X1   g0460(.A1(new_n347), .A2(new_n532), .A3(new_n577), .A4(new_n660), .ZN(G372));
  XNOR2_X1  g0461(.A(new_n428), .B(KEYINPUT18), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n449), .A2(new_n462), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n496), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n494), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n662), .B1(new_n665), .B2(new_n421), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n527), .A2(new_n528), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n530), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n602), .A2(new_n499), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n607), .A2(new_n608), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n614), .B1(new_n670), .B2(G190), .ZN(new_n671));
  INV_X1    g0471(.A(new_n615), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n626), .B(new_n669), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT26), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n602), .A2(new_n460), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n587), .A2(new_n606), .A3(new_n675), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n673), .A2(new_n674), .A3(new_n318), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n676), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n674), .B1(new_n627), .B2(new_n318), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n572), .A2(new_n542), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n657), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n673), .A2(new_n676), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n347), .A4(new_n576), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n668), .B1(new_n532), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT93), .ZN(G369));
  AND3_X1   g0487(.A1(new_n652), .A2(new_n653), .A3(new_n651), .ZN(new_n688));
  OAI22_X1  g0488(.A1(new_n688), .A2(new_n654), .B1(new_n649), .B2(new_n641), .ZN(new_n689));
  INV_X1    g0489(.A(new_n278), .ZN(new_n690));
  OR3_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .A3(G20), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT27), .B1(new_n690), .B2(G20), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n689), .A2(new_n637), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT94), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n637), .A2(new_n695), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n657), .A2(new_n659), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(new_n696), .A3(new_n697), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  INV_X1    g0503(.A(new_n695), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n573), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n572), .A2(new_n695), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(new_n577), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n657), .A2(new_n695), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n577), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n681), .B2(new_n695), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n708), .A2(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n207), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n584), .A2(new_n634), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n714), .A2(new_n715), .A3(new_n203), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n211), .B2(new_n714), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n717), .B(KEYINPUT28), .Z(new_n718));
  NAND2_X1  g0518(.A1(new_n685), .A2(new_n704), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT96), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n683), .A2(new_n347), .A3(new_n576), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n689), .B1(new_n572), .B2(new_n544), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n676), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n611), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n626), .B(new_n724), .C1(new_n671), .C2(new_n672), .ZN(new_n725));
  INV_X1    g0525(.A(new_n610), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n725), .A2(new_n318), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(KEYINPUT26), .ZN(new_n728));
  AND4_X1   g0528(.A1(KEYINPUT26), .A2(new_n673), .A3(new_n318), .A4(new_n676), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n704), .B1(new_n723), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n720), .A2(KEYINPUT29), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT96), .B1(new_n685), .B2(new_n704), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n733), .A2(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n577), .A2(new_n660), .A3(new_n347), .A4(new_n704), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n649), .A2(new_n608), .A3(new_n607), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n314), .A2(new_n638), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n541), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  AND4_X1   g0541(.A1(new_n315), .A2(new_n539), .A3(new_n328), .A4(new_n602), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n740), .A2(new_n741), .B1(new_n652), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT95), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n537), .A2(new_n538), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n745), .A2(G179), .A3(new_n314), .A4(new_n638), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n603), .B(new_n605), .C1(new_n648), .C2(new_n647), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n744), .B1(new_n748), .B2(KEYINPUT30), .ZN(new_n749));
  NOR4_X1   g0549(.A1(new_n746), .A2(new_n747), .A3(KEYINPUT95), .A4(new_n741), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n743), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n695), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT31), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n736), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G330), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n735), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n718), .B1(new_n759), .B2(G1), .ZN(G364));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n702), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n271), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n203), .B1(new_n766), .B2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n714), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n713), .A2(new_n296), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n211), .B2(new_n307), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n237), .B2(new_n307), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n713), .A2(new_n363), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n774), .A2(G355), .B1(new_n634), .B2(new_n713), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n212), .B1(G20), .B2(new_n460), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n763), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n769), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(KEYINPUT97), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n332), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n315), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n260), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n204), .A2(new_n315), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n332), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n787), .B(KEYINPUT98), .Z(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n782), .ZN(new_n793));
  INV_X1    g0593(.A(G58), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n296), .B1(new_n516), .B2(new_n790), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n204), .A2(G179), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G190), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G159), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(KEYINPUT99), .B(KEYINPUT32), .Z(new_n802));
  AND2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n788), .A2(G190), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n805), .A2(new_n216), .B1(new_n801), .B2(new_n802), .ZN(new_n806));
  OR4_X1    g0606(.A1(new_n786), .A2(new_n795), .A3(new_n803), .A4(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n499), .A2(new_n332), .A3(new_n796), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n258), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n792), .A2(new_n797), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n809), .B1(new_n811), .B2(G77), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n499), .A2(G190), .A3(new_n796), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n374), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(KEYINPUT33), .B(G317), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n804), .A2(new_n815), .B1(new_n784), .B2(G294), .ZN(new_n816));
  INV_X1    g0616(.A(new_n798), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n296), .B1(new_n817), .B2(G329), .ZN(new_n818));
  INV_X1    g0618(.A(G326), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n816), .B(new_n818), .C1(new_n819), .C2(new_n790), .ZN(new_n820));
  INV_X1    g0620(.A(new_n808), .ZN(new_n821));
  INV_X1    g0621(.A(new_n813), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G283), .A2(new_n821), .B1(new_n822), .B2(G303), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  INV_X1    g0624(.A(G322), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n823), .B1(new_n824), .B2(new_n810), .C1(new_n825), .C2(new_n793), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n807), .A2(new_n814), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n777), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n780), .A2(KEYINPUT97), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n765), .A2(new_n781), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n703), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(new_n769), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n702), .A2(G330), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n831), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G396));
  AOI22_X1  g0637(.A1(new_n811), .A2(G116), .B1(G107), .B2(new_n822), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n821), .A2(G87), .ZN(new_n839));
  INV_X1    g0639(.A(G294), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n838), .B(new_n839), .C1(new_n840), .C2(new_n793), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n363), .B1(new_n798), .B2(new_n824), .ZN(new_n842));
  INV_X1    g0642(.A(G283), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n805), .A2(new_n843), .B1(new_n790), .B2(new_n644), .ZN(new_n844));
  NOR4_X1   g0644(.A1(new_n841), .A2(new_n786), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT100), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n804), .A2(G150), .B1(new_n789), .B2(G137), .ZN(new_n847));
  INV_X1    g0647(.A(G143), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n847), .B1(new_n810), .B2(new_n799), .C1(new_n848), .C2(new_n793), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT34), .ZN(new_n850));
  OR2_X1    g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n808), .A2(new_n216), .ZN(new_n852));
  INV_X1    g0652(.A(G132), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n296), .B1(new_n798), .B2(new_n853), .C1(new_n785), .C2(new_n794), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n852), .B(new_n854), .C1(G50), .C2(new_n822), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n850), .B2(new_n849), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n777), .B1(new_n846), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n769), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n777), .A2(new_n761), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n859), .B1(new_n435), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n501), .B1(new_n449), .B2(new_n704), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n463), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n663), .A2(new_n704), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n858), .B(new_n861), .C1(new_n866), .C2(new_n762), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n463), .A2(new_n501), .A3(new_n704), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n680), .B2(new_n684), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n719), .B2(new_n865), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n769), .B1(new_n871), .B2(new_n757), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n871), .A2(new_n757), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n867), .B1(new_n873), .B2(new_n874), .ZN(G384));
  OR2_X1    g0675(.A1(new_n264), .A2(KEYINPUT35), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n264), .A2(KEYINPUT35), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n876), .A2(G116), .A3(new_n213), .A4(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT36), .ZN(new_n879));
  INV_X1    g0679(.A(new_n211), .ZN(new_n880));
  OAI21_X1  g0680(.A(G77), .B1(new_n794), .B2(new_n216), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n880), .A2(new_n881), .B1(G50), .B2(new_n216), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(G1), .A3(new_n271), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT101), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT103), .ZN(new_n886));
  XNOR2_X1  g0686(.A(KEYINPUT102), .B(KEYINPUT37), .ZN(new_n887));
  INV_X1    g0687(.A(new_n693), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n368), .A2(new_n888), .ZN(new_n889));
  AND4_X1   g0689(.A1(new_n428), .A2(new_n418), .A3(new_n887), .A4(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT37), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n406), .B1(new_n408), .B2(new_n411), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(new_n366), .A3(new_n466), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n693), .B1(new_n893), .B2(new_n355), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n403), .B2(new_n414), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n355), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n427), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n891), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n886), .B1(new_n890), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n894), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n897), .A2(new_n418), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n428), .A2(new_n418), .A3(new_n887), .A4(new_n889), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(KEYINPUT103), .A3(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n900), .B1(new_n421), .B2(new_n429), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n885), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT79), .B1(new_n397), .B2(new_n398), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n418), .A2(new_n417), .A3(KEYINPUT17), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT80), .B1(new_n418), .B2(KEYINPUT17), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n908), .A2(new_n909), .B1(new_n910), .B2(new_n415), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n894), .B1(new_n911), .B2(new_n662), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n899), .A2(new_n904), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(KEYINPUT38), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n907), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n494), .A2(new_n496), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n473), .A2(new_n704), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n917), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n494), .B2(new_n496), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n868), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n676), .B(new_n677), .C1(new_n727), .C2(new_n674), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n689), .B1(new_n572), .B2(new_n542), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n576), .A2(new_n673), .A3(new_n676), .ZN(new_n925));
  INV_X1    g0725(.A(new_n318), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n334), .A2(new_n338), .A3(new_n319), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT83), .B1(new_n345), .B2(new_n285), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n924), .A2(new_n925), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n922), .B1(new_n923), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n921), .B1(new_n931), .B2(new_n864), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n915), .A2(new_n932), .B1(new_n662), .B2(new_n693), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n912), .A2(KEYINPUT38), .A3(new_n913), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT38), .B1(new_n912), .B2(new_n913), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT39), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT104), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n915), .A2(KEYINPUT104), .A3(KEYINPUT39), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n889), .B1(new_n421), .B2(new_n429), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n428), .A2(new_n418), .A3(new_n889), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(new_n887), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n885), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n943), .A2(new_n914), .ZN(new_n944));
  XNOR2_X1  g0744(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n938), .A2(new_n939), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n491), .A2(new_n493), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(new_n474), .A3(new_n704), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n933), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n735), .A2(new_n532), .ZN(new_n950));
  INV_X1    g0750(.A(new_n668), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n949), .B(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(G330), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n752), .A2(KEYINPUT106), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT106), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n751), .A2(new_n956), .A3(KEYINPUT31), .A4(new_n695), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n736), .A2(new_n955), .A3(new_n957), .A4(new_n755), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n921), .A2(new_n865), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(KEYINPUT40), .B1(new_n944), .B2(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n958), .A2(new_n959), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT40), .B1(new_n907), .B2(new_n914), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n958), .A2(new_n532), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n954), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n966), .B2(new_n965), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n953), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n203), .B2(new_n766), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n953), .A2(new_n968), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n879), .B(new_n884), .C1(new_n970), .C2(new_n971), .ZN(G367));
  OAI21_X1  g0772(.A(new_n347), .B1(new_n285), .B2(new_n704), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n318), .A2(new_n695), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n975), .A2(new_n710), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT42), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n927), .A2(new_n928), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n926), .B1(new_n979), .B2(new_n573), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n977), .A2(KEYINPUT42), .B1(new_n704), .B2(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n626), .A2(new_n704), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n683), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n676), .B2(new_n982), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n978), .A2(new_n981), .B1(KEYINPUT43), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n985), .B(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n708), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n988), .A2(new_n975), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n987), .B(new_n989), .Z(new_n990));
  XOR2_X1   g0790(.A(new_n714), .B(KEYINPUT41), .Z(new_n991));
  INV_X1    g0791(.A(new_n709), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n707), .A2(KEYINPUT108), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n710), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT108), .B1(new_n707), .B2(new_n992), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(new_n703), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n759), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT109), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(KEYINPUT109), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n711), .A2(new_n975), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT44), .Z(new_n1003));
  NOR2_X1   g0803(.A1(new_n711), .A2(new_n975), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n708), .A2(KEYINPUT107), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1001), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n991), .B1(new_n1009), .B2(new_n759), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n990), .B1(new_n1010), .B2(new_n768), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n770), .A2(new_n233), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1012), .B(new_n778), .C1(new_n207), .C2(new_n441), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT110), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n859), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n1014), .B2(new_n1013), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n785), .A2(new_n216), .ZN(new_n1017));
  INV_X1    g0817(.A(G137), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n296), .B1(new_n798), .B2(new_n1018), .C1(new_n805), .C2(new_n799), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1017), .B(new_n1019), .C1(G143), .C2(new_n789), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G58), .A2(new_n822), .B1(new_n821), .B2(G77), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n793), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n811), .A2(G50), .B1(new_n1022), .B2(G150), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n811), .A2(G283), .B1(G97), .B2(new_n821), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n644), .B2(new_n793), .ZN(new_n1026));
  INV_X1    g0826(.A(G317), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n363), .B1(new_n798), .B2(new_n1027), .C1(new_n790), .C2(new_n824), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n805), .A2(new_n840), .B1(new_n785), .B2(new_n258), .ZN(new_n1029));
  OR3_X1    g0829(.A1(new_n1026), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n813), .A2(new_n634), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT46), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1024), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT47), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1016), .B1(new_n1034), .B2(new_n777), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n764), .B2(new_n984), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1011), .A2(new_n1036), .ZN(G387));
  NAND2_X1  g0837(.A1(new_n999), .A2(new_n1000), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n759), .A2(new_n997), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n714), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n777), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n644), .A2(new_n810), .B1(new_n793), .B2(new_n1027), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT111), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n804), .A2(G311), .B1(new_n789), .B2(G322), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  OR3_X1    g0849(.A1(new_n1046), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1049), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n822), .A2(G294), .B1(G283), .B2(new_n784), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT49), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n363), .B1(new_n819), .B2(new_n798), .C1(new_n808), .C2(new_n634), .ZN(new_n1057));
  OR3_X1    g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n785), .A2(new_n441), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n296), .B1(new_n798), .B2(new_n513), .C1(new_n790), .C2(new_n799), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n353), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1059), .B(new_n1060), .C1(new_n1061), .C2(new_n804), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1022), .A2(G50), .B1(G97), .B2(new_n821), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n811), .A2(G68), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n822), .A2(G77), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1043), .B1(new_n1058), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n353), .A2(G50), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT50), .ZN(new_n1069));
  AOI211_X1 g0869(.A(G45), .B(new_n715), .C1(G68), .C2(G77), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n771), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n307), .B2(new_n230), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n774), .A2(new_n715), .B1(new_n258), .B2(new_n713), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n769), .B1(new_n1075), .B2(new_n779), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n1067), .A2(KEYINPUT112), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n707), .B2(new_n763), .ZN(new_n1078));
  OAI21_X1  g0878(.A(KEYINPUT112), .B1(new_n1067), .B2(new_n1076), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1078), .A2(new_n1079), .B1(new_n768), .B2(new_n997), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1042), .A2(new_n1080), .ZN(G393));
  INV_X1    g0881(.A(new_n1006), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT113), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n1082), .A2(new_n1083), .A3(new_n988), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT113), .B1(new_n1006), .B2(new_n708), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1006), .A2(new_n708), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1009), .B(new_n714), .C1(new_n1001), .C2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n975), .A2(new_n763), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n778), .B1(new_n260), .B2(new_n207), .C1(new_n771), .C2(new_n240), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n769), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n793), .A2(new_n799), .B1(new_n513), .B2(new_n790), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT51), .Z(new_n1093));
  NOR2_X1   g0893(.A1(new_n785), .A2(new_n435), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n296), .B1(new_n798), .B2(new_n848), .C1(new_n805), .C2(new_n516), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n811), .A2(new_n1061), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n822), .A2(G68), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n839), .A3(new_n1097), .ZN(new_n1098));
  NOR4_X1   g0898(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1100), .A2(KEYINPUT114), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n793), .A2(new_n824), .B1(new_n1027), .B2(new_n790), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT52), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n813), .A2(new_n843), .B1(new_n825), .B2(new_n798), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT115), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n363), .B1(new_n785), .B2(new_n634), .C1(new_n805), .C2(new_n644), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n809), .B(new_n1108), .C1(new_n811), .C2(G294), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1103), .A2(new_n1106), .A3(new_n1107), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1100), .A2(KEYINPUT114), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1101), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1091), .B1(new_n1112), .B2(new_n777), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1087), .A2(new_n768), .B1(new_n1089), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1088), .A2(new_n1114), .ZN(G390));
  INV_X1    g0915(.A(new_n948), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n944), .A2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n704), .B(new_n863), .C1(new_n723), .C2(new_n730), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n864), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n921), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n944), .A2(new_n945), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT104), .B1(new_n915), .B2(KEYINPUT39), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT39), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n937), .B(new_n1125), .C1(new_n907), .C2(new_n914), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1123), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT116), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n932), .B2(new_n1116), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n864), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1120), .B1(new_n869), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(KEYINPUT116), .A3(new_n948), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1122), .B1(new_n1127), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n958), .A2(new_n959), .A3(G330), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n932), .A2(new_n1128), .A3(new_n1116), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT116), .B1(new_n1131), .B2(new_n948), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n938), .A2(new_n939), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n1140), .A3(new_n1123), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n756), .A2(G330), .A3(new_n866), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1142), .A2(new_n921), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1134), .A2(new_n1136), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n958), .A2(G330), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n532), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n950), .A2(new_n951), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1143), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1119), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1146), .A2(new_n866), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1149), .B(new_n1150), .C1(new_n1151), .C2(new_n1120), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n869), .A2(new_n1130), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1142), .A2(new_n921), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1153), .B1(new_n1154), .B2(new_n1135), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT117), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI211_X1 g0957(.A(KEYINPUT117), .B(new_n1153), .C1(new_n1154), .C2(new_n1135), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1152), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1145), .A2(new_n1148), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1144), .B1(new_n1127), .B2(new_n1133), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n946), .A2(new_n1139), .B1(new_n1121), .B2(new_n1117), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1161), .B1(new_n1162), .B2(new_n1135), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1159), .A2(new_n1148), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1160), .A2(new_n1165), .A3(new_n714), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT121), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1161), .A2(new_n768), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1135), .B1(new_n1141), .B2(new_n1122), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT118), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n767), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT118), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n859), .B1(new_n353), .B2(new_n860), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n852), .B1(G87), .B2(new_n822), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n634), .B2(new_n793), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n790), .A2(new_n843), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n363), .B1(new_n798), .B2(new_n840), .ZN(new_n1180));
  NOR4_X1   g0980(.A1(new_n1178), .A2(new_n1094), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n810), .A2(new_n260), .B1(new_n258), .B2(new_n805), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT120), .Z(new_n1183));
  NAND2_X1  g0983(.A1(new_n822), .A2(G150), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT53), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n785), .A2(new_n799), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT54), .B(G143), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n810), .A2(new_n1187), .B1(new_n516), .B2(new_n808), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n363), .B1(new_n817), .B2(G125), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n805), .B2(new_n1018), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .A4(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(G128), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n793), .A2(new_n853), .B1(new_n1192), .B2(new_n790), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT119), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1181), .A2(new_n1183), .B1(new_n1191), .B2(new_n1194), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1176), .B1(new_n1043), .B2(new_n1195), .C1(new_n1127), .C2(new_n762), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1167), .B1(new_n1175), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1196), .ZN(new_n1198));
  AOI211_X1 g0998(.A(KEYINPUT121), .B(new_n1198), .C1(new_n1170), .C2(new_n1174), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1166), .B1(new_n1197), .B2(new_n1199), .ZN(G378));
  NAND2_X1  g1000(.A1(new_n943), .A2(new_n914), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n958), .A3(new_n959), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1202), .A2(KEYINPUT40), .B1(new_n962), .B2(new_n963), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n519), .A2(new_n888), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n531), .B(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1203), .A2(new_n1209), .A3(new_n954), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1209), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n965), .B2(G330), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n949), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1209), .B1(new_n1203), .B2(new_n954), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n965), .A2(G330), .A3(new_n1211), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1127), .A2(new_n1116), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n933), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1213), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1209), .A2(new_n761), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n810), .A2(new_n1018), .B1(new_n853), .B2(new_n805), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT122), .Z(new_n1221));
  AOI22_X1  g1021(.A1(new_n789), .A2(G125), .B1(new_n784), .B2(G150), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n813), .B2(new_n1187), .C1(new_n793), .C2(new_n1192), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  OR2_X1    g1024(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n821), .A2(G159), .ZN(new_n1227));
  AOI211_X1 g1027(.A(G33), .B(G41), .C1(new_n817), .C2(G124), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(G41), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G50), .B1(new_n246), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n296), .B2(G41), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n811), .A2(new_n440), .B1(new_n1022), .B2(G107), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n821), .A2(G58), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n1065), .A3(new_n1234), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1230), .B(new_n363), .C1(new_n798), .C2(new_n843), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n805), .A2(new_n260), .B1(new_n790), .B2(new_n634), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(new_n1235), .A2(new_n1017), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1232), .B1(new_n1238), .B2(KEYINPUT58), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(KEYINPUT58), .B2(new_n1238), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1043), .B1(new_n1229), .B2(new_n1240), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT123), .Z(new_n1242));
  AOI211_X1 g1042(.A(new_n859), .B(new_n1242), .C1(new_n516), .C2(new_n860), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1218), .A2(new_n768), .B1(new_n1219), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1218), .A2(KEYINPUT57), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1148), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1145), .B2(new_n1159), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n714), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1148), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT57), .B1(new_n1249), .B2(new_n1218), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1244), .B1(new_n1248), .B2(new_n1250), .ZN(G375));
  OR2_X1    g1051(.A1(new_n1159), .A2(new_n1148), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n991), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(new_n1253), .A3(new_n1164), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1159), .A2(new_n768), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n296), .B1(new_n798), .B2(new_n1192), .C1(new_n785), .C2(new_n516), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n1018), .A2(new_n793), .B1(new_n810), .B2(new_n513), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1234), .B1(new_n799), .B2(new_n813), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n853), .A2(new_n790), .B1(new_n805), .B2(new_n1187), .ZN(new_n1259));
  OR4_X1    g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n363), .B1(new_n798), .B2(new_n644), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1261), .B(new_n1059), .C1(G294), .C2(new_n789), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G77), .A2(new_n821), .B1(new_n822), .B2(G97), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1262), .B(new_n1263), .C1(new_n843), .C2(new_n793), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n810), .A2(new_n258), .B1(new_n634), .B2(new_n805), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(KEYINPUT124), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1260), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n777), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n859), .B1(new_n216), .B2(new_n860), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(new_n1120), .C2(new_n762), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1255), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1254), .A2(new_n1272), .ZN(G381));
  INV_X1    g1073(.A(G390), .ZN(new_n1274));
  INV_X1    g1074(.A(G384), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1042), .A2(new_n836), .A3(new_n1080), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1277), .A2(G387), .A3(G381), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1243), .A2(new_n1219), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1218), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(new_n767), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT57), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n1280), .B2(new_n1247), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1282), .B1(new_n1213), .B2(new_n1217), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1040), .B1(new_n1249), .B2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1281), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1160), .A2(new_n714), .A3(new_n1165), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1173), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1196), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1278), .A2(new_n1286), .A3(new_n1291), .ZN(G407));
  NAND2_X1  g1092(.A1(new_n694), .A2(G213), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1286), .A2(new_n1291), .A3(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(G407), .A2(G213), .A3(new_n1295), .ZN(G409));
  AOI21_X1  g1096(.A(new_n836), .B1(new_n1042), .B2(new_n1080), .ZN(new_n1297));
  OAI21_X1  g1097(.A(KEYINPUT125), .B1(new_n1276), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G393), .A2(G396), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT125), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1042), .A2(new_n836), .A3(new_n1080), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1298), .A2(new_n1302), .A3(G390), .ZN(new_n1303));
  AOI21_X1  g1103(.A(G390), .B1(new_n1302), .B2(new_n1298), .ZN(new_n1304));
  OAI21_X1  g1104(.A(G387), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1298), .A2(new_n1302), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1274), .ZN(new_n1307));
  INV_X1    g1107(.A(G387), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1298), .A2(new_n1302), .A3(G390), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1307), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1305), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1249), .A2(new_n1253), .A3(new_n1218), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1244), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(G378), .A2(new_n1286), .B1(new_n1291), .B2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(KEYINPUT126), .B1(new_n1314), .B2(new_n1294), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1291), .A2(new_n1313), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1290), .A2(KEYINPUT121), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1175), .A2(new_n1167), .A3(new_n1196), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1287), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1316), .B1(new_n1319), .B2(G375), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT126), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n1321), .A3(new_n1293), .ZN(new_n1322));
  AND2_X1   g1122(.A1(new_n1164), .A2(KEYINPUT60), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1252), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1040), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1164), .A2(KEYINPUT60), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1252), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(G384), .B1(new_n1328), .B2(new_n1272), .ZN(new_n1329));
  AOI211_X1 g1129(.A(new_n1275), .B(new_n1271), .C1(new_n1325), .C2(new_n1327), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT62), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(new_n1329), .A2(new_n1330), .A3(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1315), .A2(new_n1322), .A3(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1320), .A2(new_n1293), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1331), .B1(new_n1334), .B2(new_n1336), .ZN(new_n1337));
  AND2_X1   g1137(.A1(new_n1333), .A2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1328), .A2(new_n1272), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1275), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1328), .A2(G384), .A3(new_n1272), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1340), .A2(G2897), .A3(new_n1294), .A4(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1294), .A2(G2897), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1343), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1342), .A2(new_n1344), .ZN(new_n1345));
  NOR3_X1   g1145(.A1(new_n1314), .A2(KEYINPUT126), .A3(new_n1294), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1321), .B1(new_n1320), .B2(new_n1293), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1345), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT61), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1311), .B1(new_n1338), .B2(new_n1350), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1311), .A2(KEYINPUT61), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1315), .A2(new_n1322), .A3(KEYINPUT63), .A4(new_n1335), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT63), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1354), .B1(new_n1334), .B2(new_n1336), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1345), .A2(new_n1334), .ZN(new_n1356));
  NAND4_X1  g1156(.A1(new_n1352), .A2(new_n1353), .A3(new_n1355), .A4(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1351), .A2(new_n1357), .ZN(G405));
  AND2_X1   g1158(.A1(new_n1305), .A2(new_n1310), .ZN(new_n1359));
  OR2_X1    g1159(.A1(new_n1335), .A2(KEYINPUT127), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1335), .A2(KEYINPUT127), .ZN(new_n1361));
  NOR2_X1   g1161(.A1(new_n1319), .A2(G375), .ZN(new_n1362));
  AND2_X1   g1162(.A1(G375), .A2(new_n1291), .ZN(new_n1363));
  OAI211_X1 g1163(.A(new_n1360), .B(new_n1361), .C1(new_n1362), .C2(new_n1363), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1363), .A2(new_n1362), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1365), .A2(KEYINPUT127), .A3(new_n1335), .ZN(new_n1366));
  AND3_X1   g1166(.A1(new_n1359), .A2(new_n1364), .A3(new_n1366), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1359), .B1(new_n1364), .B2(new_n1366), .ZN(new_n1368));
  NOR2_X1   g1168(.A1(new_n1367), .A2(new_n1368), .ZN(G402));
endmodule


