//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1292, new_n1293,
    new_n1294;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n215));
  XOR2_X1   g0015(.A(new_n214), .B(new_n215), .Z(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n202), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n206), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n212), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n203), .A2(G50), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR3_X1   g0033(.A1(new_n216), .A2(new_n228), .A3(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT65), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G200), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n255));
  NOR3_X1   g0055(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n255), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n256), .B1(G226), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT3), .B(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G222), .A2(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G223), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n264), .B(new_n253), .C1(G77), .C2(new_n260), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n252), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n259), .A2(new_n265), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n266), .B1(new_n268), .B2(G190), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n229), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT66), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT66), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n270), .A2(new_n273), .A3(new_n229), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G150), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT8), .B(G58), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n210), .A2(G33), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G58), .A2(G68), .ZN(new_n281));
  INV_X1    g0081(.A(G50), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n210), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n275), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n282), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n275), .A2(new_n286), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n209), .A2(G20), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(G50), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(KEYINPUT9), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT9), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n288), .B2(new_n291), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n269), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n269), .B(new_n298), .C1(new_n293), .C2(new_n295), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n268), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n267), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(new_n292), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT67), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n301), .A2(new_n292), .A3(KEYINPUT67), .A4(new_n303), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n297), .A2(new_n299), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n260), .A2(G232), .A3(new_n262), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(new_n206), .B2(new_n260), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G33), .ZN(new_n312));
  INV_X1    g0112(.A(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT3), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n315), .A2(new_n218), .A3(new_n262), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n253), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT68), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n256), .B1(G244), .B2(new_n258), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n318), .B1(new_n317), .B2(new_n319), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n300), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n322), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(new_n302), .A3(new_n320), .ZN(new_n325));
  INV_X1    g0125(.A(new_n271), .ZN(new_n326));
  INV_X1    g0126(.A(new_n278), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(new_n276), .B1(G20), .B2(G77), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT15), .B(G87), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n329), .A2(new_n279), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n326), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n286), .A2(new_n271), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(G77), .A3(new_n290), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(G77), .B2(new_n285), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n323), .A2(new_n325), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(G190), .B1(new_n321), .B2(new_n322), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n324), .A2(G200), .A3(new_n320), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n339), .A3(new_n335), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n337), .A2(new_n340), .A3(KEYINPUT69), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT69), .B1(new_n337), .B2(new_n340), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n308), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n276), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(new_n223), .B2(new_n279), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n275), .A2(new_n345), .ZN(new_n346));
  XOR2_X1   g0146(.A(new_n346), .B(KEYINPUT11), .Z(new_n347));
  INV_X1    g0147(.A(KEYINPUT72), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT73), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n285), .A2(G68), .B1(new_n350), .B2(KEYINPUT12), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT12), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(KEYINPUT73), .B2(new_n352), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n350), .B(KEYINPUT12), .C1(new_n285), .C2(G68), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n202), .B1(new_n209), .B2(G20), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n353), .A2(new_n354), .B1(new_n332), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n347), .B2(new_n348), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G41), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n230), .B1(new_n313), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G226), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(G1698), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(new_n312), .A3(new_n314), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT70), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n260), .A2(KEYINPUT70), .A3(new_n362), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n312), .A2(new_n314), .A3(G232), .A4(G1698), .ZN(new_n368));
  AND3_X1   g0168(.A1(KEYINPUT71), .A2(G33), .A3(G97), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT71), .B1(G33), .B2(G97), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n360), .B1(new_n367), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n360), .A2(G274), .A3(new_n257), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n360), .A2(new_n255), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(new_n218), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT13), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n377), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT13), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n372), .B1(new_n365), .B2(new_n366), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n379), .B(new_n380), .C1(new_n360), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT14), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n384), .A3(G169), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n378), .A2(new_n382), .A3(G179), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT74), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n384), .B1(new_n383), .B2(G169), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n385), .A2(new_n386), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT74), .B1(new_n392), .B2(new_n389), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n358), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n367), .A2(new_n373), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n253), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n380), .B1(new_n396), .B2(new_n379), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n374), .A2(KEYINPUT13), .A3(new_n377), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G190), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n358), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n399), .A2(new_n252), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n343), .A2(new_n394), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n278), .B1(new_n209), .B2(G20), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n289), .A2(new_n405), .B1(new_n286), .B2(new_n278), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n361), .A2(G1698), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n260), .B(new_n407), .C1(G223), .C2(G1698), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G87), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n253), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n256), .B1(G232), .B2(new_n258), .ZN(new_n412));
  INV_X1    g0212(.A(G190), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n360), .B1(new_n408), .B2(new_n409), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n375), .B1(new_n376), .B2(new_n236), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n252), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT75), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n313), .B2(KEYINPUT3), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n311), .A2(KEYINPUT75), .A3(G33), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(new_n421), .A3(new_n314), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT7), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(G20), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(KEYINPUT76), .A3(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n423), .B1(new_n260), .B2(G20), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT76), .B1(new_n422), .B2(new_n424), .ZN(new_n428));
  OAI21_X1  g0228(.A(G68), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n201), .A2(new_n202), .ZN(new_n430));
  OAI21_X1  g0230(.A(G20), .B1(new_n430), .B2(new_n281), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n276), .A2(G159), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT16), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n315), .A2(new_n210), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n436), .A2(new_n423), .B1(new_n424), .B2(new_n315), .ZN(new_n437));
  OAI211_X1 g0237(.A(KEYINPUT16), .B(new_n434), .C1(new_n437), .C2(new_n202), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n271), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n406), .B(new_n418), .C1(new_n435), .C2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT17), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n315), .A2(new_n424), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n426), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n433), .B1(new_n444), .B2(G68), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n326), .B1(new_n445), .B2(KEYINPUT16), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n422), .A2(new_n424), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT76), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(new_n426), .A3(new_n425), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n433), .B1(new_n450), .B2(G68), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n446), .B1(new_n451), .B2(KEYINPUT16), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n452), .A2(KEYINPUT17), .A3(new_n406), .A4(new_n418), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n442), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT77), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n406), .B1(new_n435), .B2(new_n439), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT18), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n411), .A2(new_n412), .A3(G179), .ZN(new_n459));
  OAI21_X1  g0259(.A(G169), .B1(new_n415), .B2(new_n416), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n457), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n458), .B1(new_n457), .B2(new_n461), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n442), .A2(new_n453), .A3(KEYINPUT77), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n456), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT78), .ZN(new_n467));
  OR2_X1    g0267(.A1(new_n466), .A2(KEYINPUT78), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n404), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G303), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n315), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(G257), .A2(G1698), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(new_n225), .B2(G1698), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n471), .B(new_n253), .C1(new_n315), .C2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G45), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G1), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT5), .B(G41), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n360), .A2(G274), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n476), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(G270), .A3(new_n360), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n474), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT84), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n474), .A2(KEYINPUT84), .A3(new_n478), .A4(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G190), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(G200), .A3(new_n484), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n488), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n489));
  INV_X1    g0289(.A(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G20), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n271), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT20), .ZN(new_n493));
  XNOR2_X1  g0293(.A(new_n492), .B(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT85), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n285), .B2(G116), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n286), .A2(KEYINPUT85), .A3(new_n490), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n490), .B1(new_n209), .B2(G33), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n496), .A2(new_n497), .B1(new_n332), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n486), .A2(new_n487), .A3(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n312), .A2(new_n314), .A3(new_n210), .A4(G87), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT22), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT22), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n260), .A2(new_n505), .A3(new_n210), .A4(G87), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n279), .A2(new_n490), .ZN(new_n508));
  OAI21_X1  g0308(.A(KEYINPUT87), .B1(new_n210), .B2(G107), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT23), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT23), .ZN(new_n511));
  OAI211_X1 g0311(.A(KEYINPUT87), .B(new_n511), .C1(new_n210), .C2(G107), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n508), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(KEYINPUT24), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT24), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n507), .B2(new_n513), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n271), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n286), .A2(new_n206), .ZN(new_n519));
  XNOR2_X1  g0319(.A(new_n519), .B(KEYINPUT25), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n209), .A2(G33), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n272), .A2(new_n285), .A3(new_n274), .A4(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n520), .B1(new_n523), .B2(G107), .ZN(new_n524));
  MUX2_X1   g0324(.A(G250), .B(G257), .S(G1698), .Z(new_n525));
  XNOR2_X1  g0325(.A(KEYINPUT88), .B(G294), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n525), .A2(new_n260), .B1(new_n526), .B2(G33), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n253), .B1(new_n476), .B2(new_n477), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n528), .A2(new_n253), .B1(G264), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(G190), .A3(new_n478), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(G264), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n532), .B(new_n478), .C1(new_n360), .C2(new_n527), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G200), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n518), .A2(new_n524), .A3(new_n531), .A4(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n260), .A2(new_n210), .A3(G68), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT19), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n279), .B2(new_n205), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n207), .A2(G87), .ZN(new_n540));
  OAI21_X1  g0340(.A(KEYINPUT19), .B1(new_n369), .B2(new_n370), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(new_n210), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n271), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n329), .A2(new_n286), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n543), .B(new_n544), .C1(new_n329), .C2(new_n522), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n360), .A2(G274), .A3(new_n476), .ZN(new_n546));
  NOR2_X1   g0346(.A1(G238), .A2(G1698), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n224), .B2(G1698), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(new_n260), .B1(G33), .B2(G116), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n546), .B1(new_n549), .B2(new_n360), .ZN(new_n550));
  NOR4_X1   g0350(.A1(new_n253), .A2(KEYINPUT83), .A3(new_n476), .A4(new_n220), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT83), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n476), .A2(new_n220), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n360), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n302), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g0356(.A1(new_n549), .A2(new_n360), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n360), .A2(new_n553), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT83), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n360), .A2(new_n553), .A3(new_n552), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n557), .A2(new_n561), .A3(new_n300), .A4(new_n546), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n545), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n543), .A2(new_n544), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n557), .A2(new_n561), .A3(G190), .A4(new_n546), .ZN(new_n565));
  OAI21_X1  g0365(.A(G200), .B1(new_n550), .B2(new_n555), .ZN(new_n566));
  OR2_X1    g0366(.A1(new_n522), .A2(new_n219), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n564), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n502), .A2(new_n535), .A3(new_n563), .A4(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n479), .A2(G257), .A3(new_n360), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n478), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT81), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT4), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n262), .A2(G244), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n573), .B1(new_n315), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n260), .A2(KEYINPUT4), .A3(G244), .A4(new_n262), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n260), .A2(G250), .A3(G1698), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n488), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n253), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT81), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n570), .A2(new_n580), .A3(new_n478), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n572), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n302), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n572), .A2(new_n579), .A3(new_n581), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n300), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT79), .ZN(new_n586));
  INV_X1    g0386(.A(new_n276), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT6), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n588), .A2(new_n205), .A3(G107), .ZN(new_n589));
  XNOR2_X1  g0389(.A(G97), .B(G107), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  OAI221_X1 g0391(.A(new_n586), .B1(new_n223), .B2(new_n587), .C1(new_n591), .C2(new_n210), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n588), .ZN(new_n593));
  INV_X1    g0393(.A(new_n589), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n210), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n587), .A2(new_n223), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT79), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n450), .A2(G107), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n326), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n522), .A2(G97), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n285), .A2(new_n205), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n603), .B(KEYINPUT80), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n583), .B(new_n585), .C1(new_n600), .C2(new_n604), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n450), .A2(G107), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n592), .A2(new_n597), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n271), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT80), .ZN(new_n609));
  XNOR2_X1  g0409(.A(new_n603), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n582), .A2(G200), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n572), .A2(new_n579), .A3(G190), .A4(new_n581), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n608), .A2(new_n610), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT82), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n569), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n605), .A2(new_n613), .A3(KEYINPUT82), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n483), .A2(new_n500), .A3(G169), .A4(new_n484), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT21), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n474), .A2(G179), .A3(new_n478), .A4(new_n480), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n618), .A2(new_n619), .B1(new_n500), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n483), .A2(new_n484), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT86), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n302), .B1(new_n494), .B2(new_n499), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT21), .A4(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT86), .B1(new_n618), .B2(new_n619), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n622), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT89), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n533), .A2(new_n629), .A3(G169), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n530), .A2(G179), .A3(new_n478), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n533), .A2(G169), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(KEYINPUT89), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n632), .A2(new_n634), .B1(new_n518), .B2(new_n524), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n628), .A2(new_n635), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n469), .A2(new_n616), .A3(new_n617), .A4(new_n636), .ZN(G372));
  AND2_X1   g0437(.A1(new_n622), .A2(new_n626), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT90), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n632), .A2(new_n634), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n518), .A2(new_n524), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n638), .A2(new_n639), .A3(new_n642), .A4(new_n627), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n568), .A2(new_n563), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n605), .A2(new_n645), .A3(new_n613), .A4(new_n535), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT90), .B1(new_n628), .B2(new_n635), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n643), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n563), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n605), .B2(new_n644), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n585), .A2(new_n583), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n608), .A2(new_n610), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n645), .A2(new_n652), .A3(KEYINPUT26), .A4(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n649), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n648), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n469), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n306), .A2(new_n307), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n297), .A2(new_n299), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT91), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n297), .A2(KEYINPUT91), .A3(new_n299), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n456), .A2(new_n465), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n403), .A2(new_n337), .ZN(new_n665));
  INV_X1    g0465(.A(new_n358), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n388), .B1(new_n387), .B2(new_n390), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n392), .A2(new_n389), .A3(KEYINPUT74), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n664), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n464), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n663), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n657), .A2(new_n658), .A3(new_n672), .ZN(G369));
  INV_X1    g0473(.A(G13), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n674), .A2(G1), .A3(G20), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT92), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT27), .ZN(new_n677));
  OAI21_X1  g0477(.A(G213), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT93), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT93), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G343), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n641), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n642), .A2(new_n685), .A3(new_n535), .ZN(new_n686));
  XOR2_X1   g0486(.A(new_n686), .B(KEYINPUT94), .Z(new_n687));
  NAND2_X1  g0487(.A1(new_n635), .A2(new_n684), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n502), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n683), .A2(new_n501), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n628), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n628), .A2(new_n691), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n690), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G330), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n628), .A2(new_n683), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n687), .A2(new_n697), .B1(new_n642), .B2(new_n684), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n696), .A2(new_n698), .ZN(G399));
  NAND2_X1  g0499(.A1(new_n213), .A2(new_n359), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n540), .A2(new_n490), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n232), .B2(new_n700), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT97), .ZN(new_n706));
  OAI211_X1 g0506(.A(new_n706), .B(new_n650), .C1(new_n605), .C2(new_n644), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n563), .B(KEYINPUT96), .Z(new_n708));
  NAND4_X1  g0508(.A1(new_n605), .A2(new_n645), .A3(new_n613), .A4(new_n535), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n707), .B(new_n708), .C1(new_n636), .C2(new_n709), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n651), .A2(new_n654), .A3(KEYINPUT97), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n683), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n616), .A2(new_n617), .A3(new_n636), .A4(new_n683), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n550), .A2(new_n555), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n621), .A2(new_n715), .A3(new_n530), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(KEYINPUT30), .A3(new_n584), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n716), .B2(new_n582), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n715), .A2(G179), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n623), .A2(new_n582), .A3(new_n533), .A4(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n718), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT31), .B1(new_n723), .B2(new_n684), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n720), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT95), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n722), .A2(new_n720), .A3(KEYINPUT95), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n718), .A3(new_n728), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n684), .A2(KEYINPUT31), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n724), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n714), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G330), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n684), .B1(new_n648), .B2(new_n655), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT29), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n713), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n705), .B1(new_n737), .B2(G1), .ZN(G364));
  NOR2_X1   g0538(.A1(new_n674), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n209), .B1(new_n739), .B2(G45), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n700), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n213), .A2(new_n260), .ZN(new_n743));
  INV_X1    g0543(.A(G355), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n743), .A2(new_n744), .B1(G116), .B2(new_n213), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n213), .A2(new_n315), .ZN(new_n746));
  INV_X1    g0546(.A(new_n232), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n746), .B1(new_n475), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n250), .A2(G45), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n745), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT98), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n229), .B1(G20), .B2(new_n302), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n742), .B1(new_n750), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n210), .A2(new_n300), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(KEYINPUT33), .B(G317), .Z(new_n762));
  NOR4_X1   g0562(.A1(new_n210), .A2(new_n413), .A3(new_n252), .A4(G179), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n761), .A2(new_n762), .B1(new_n470), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n759), .A2(new_n413), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G326), .ZN(new_n768));
  INV_X1    g0568(.A(G283), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n210), .A2(new_n252), .A3(G179), .A4(G190), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n767), .A2(new_n768), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n765), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n252), .A2(G190), .ZN(new_n774));
  OAI21_X1  g0574(.A(G20), .B1(new_n774), .B2(G179), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT101), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n526), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G190), .A2(G200), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n782), .A2(G20), .A3(new_n300), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT100), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G329), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n774), .A2(new_n210), .A3(new_n300), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G322), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n315), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n758), .A2(new_n782), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n793), .B1(G311), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n773), .A2(new_n781), .A3(new_n789), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n771), .A2(new_n206), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n761), .A2(new_n202), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(G50), .C2(new_n766), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n791), .A2(new_n201), .B1(new_n794), .B2(new_n223), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT99), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n260), .B1(new_n764), .B2(new_n219), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n802), .B2(new_n801), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n780), .A2(G97), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n800), .A2(new_n803), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n788), .A2(G159), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT32), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n797), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n757), .B1(new_n810), .B2(new_n754), .ZN(new_n811));
  INV_X1    g0611(.A(new_n753), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n694), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT102), .Z(new_n814));
  NOR2_X1   g0614(.A1(new_n694), .A2(G330), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n695), .A2(new_n741), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(G396));
  NOR2_X1   g0617(.A1(new_n771), .A2(new_n219), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n761), .A2(new_n769), .B1(new_n206), .B2(new_n764), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(G303), .C2(new_n766), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n788), .A2(G311), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n315), .B1(new_n794), .B2(new_n490), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G294), .B2(new_n790), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n820), .A2(new_n806), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n795), .A2(G159), .B1(new_n790), .B2(G143), .ZN(new_n825));
  INV_X1    g0625(.A(G150), .ZN(new_n826));
  INV_X1    g0626(.A(G137), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n761), .B2(new_n826), .C1(new_n827), .C2(new_n767), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT34), .Z(new_n829));
  NOR2_X1   g0629(.A1(new_n771), .A2(new_n202), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n315), .B(new_n830), .C1(G50), .C2(new_n763), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n201), .B2(new_n779), .C1(new_n832), .C2(new_n787), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n824), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n754), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n754), .A2(new_n751), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n741), .B1(new_n223), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n340), .B1(new_n335), .B2(new_n683), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n337), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n337), .A2(new_n684), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n835), .B(new_n837), .C1(new_n842), .C2(new_n752), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n734), .B(new_n841), .ZN(new_n844));
  INV_X1    g0644(.A(new_n733), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n741), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n846), .B1(new_n848), .B2(KEYINPUT103), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n848), .A2(KEYINPUT103), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n843), .B1(new_n850), .B2(new_n851), .ZN(G384));
  NOR2_X1   g0652(.A1(new_n739), .A2(new_n209), .ZN(new_n853));
  INV_X1    g0653(.A(new_n682), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n671), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n403), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n666), .A2(new_n684), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n669), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n391), .A2(new_n393), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n666), .B(new_n684), .C1(new_n859), .C2(new_n403), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n656), .A2(new_n683), .A3(new_n842), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n840), .B(KEYINPUT105), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT38), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n457), .A2(new_n461), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n457), .A2(new_n682), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n866), .A2(new_n867), .A3(new_n868), .A4(new_n440), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n438), .A2(new_n275), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n445), .A2(KEYINPUT16), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n406), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n682), .B2(new_n461), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n440), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT37), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n872), .A2(new_n682), .ZN(new_n876));
  AOI221_X4 g0676(.A(new_n865), .B1(new_n869), .B2(new_n875), .C1(new_n466), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n466), .A2(new_n876), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n875), .A2(new_n869), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT38), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n855), .B1(new_n864), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT39), .B1(new_n877), .B2(new_n880), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT106), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n878), .A2(KEYINPUT107), .A3(KEYINPUT38), .A4(new_n879), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT107), .ZN(new_n886));
  INV_X1    g0686(.A(new_n867), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n866), .A2(KEYINPUT18), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n457), .A2(new_n458), .A3(new_n461), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n442), .A4(new_n453), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n866), .A2(new_n867), .A3(new_n440), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n887), .A2(new_n890), .B1(new_n892), .B2(new_n869), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n886), .B1(new_n893), .B2(KEYINPUT38), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n885), .B1(new_n877), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT39), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT106), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n898), .B(KEYINPUT39), .C1(new_n877), .C2(new_n880), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n884), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n394), .A2(new_n683), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n882), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n404), .A2(new_n467), .A3(new_n468), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n736), .B2(new_n713), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n672), .A2(new_n658), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n903), .B(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(G330), .ZN(new_n909));
  INV_X1    g0709(.A(new_n895), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(new_n724), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n841), .B1(new_n714), .B2(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n861), .A2(new_n913), .A3(KEYINPUT40), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n861), .B(new_n913), .C1(new_n877), .C2(new_n880), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT40), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n910), .A2(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n714), .A2(new_n912), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n404), .A2(new_n919), .A3(new_n467), .A4(new_n468), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n909), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n920), .B2(new_n918), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n853), .B1(new_n908), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n908), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g0724(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n232), .A2(new_n925), .B1(G50), .B2(new_n202), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(G1), .A3(new_n674), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT104), .ZN(new_n928));
  INV_X1    g0728(.A(new_n591), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n490), .B(new_n231), .C1(new_n929), .C2(KEYINPUT35), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(KEYINPUT35), .B2(new_n929), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT36), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n932), .B2(new_n931), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n924), .A2(new_n934), .ZN(G367));
  NAND2_X1  g0735(.A1(new_n684), .A2(new_n653), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(new_n605), .A3(new_n613), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n937), .A2(new_n642), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n684), .B1(new_n938), .B2(new_n605), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n687), .A2(new_n697), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n652), .A2(new_n653), .A3(new_n684), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n939), .B1(new_n944), .B2(KEYINPUT42), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(KEYINPUT42), .B2(new_n944), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n683), .B1(new_n564), .B2(new_n567), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n649), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n644), .B2(new_n947), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT108), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n946), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n696), .A2(new_n942), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n954), .B(new_n955), .Z(new_n956));
  XNOR2_X1  g0756(.A(new_n700), .B(KEYINPUT41), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n698), .A2(new_n943), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT45), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n698), .A2(new_n943), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT44), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n960), .A2(new_n961), .B1(new_n696), .B2(KEYINPUT110), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n959), .B(new_n962), .C1(new_n961), .C2(new_n960), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n696), .A2(KEYINPUT110), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n689), .A2(new_n697), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n940), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(new_n695), .Z(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n737), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT109), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n968), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n957), .B1(new_n974), .B2(new_n737), .ZN(new_n975));
  INV_X1    g0775(.A(new_n740), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n956), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n755), .B1(new_n213), .B2(new_n329), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n242), .A2(new_n746), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n742), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n771), .A2(new_n223), .ZN(new_n981));
  INV_X1    g0781(.A(G159), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n761), .A2(new_n982), .B1(new_n201), .B2(new_n764), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n981), .B(new_n983), .C1(G143), .C2(new_n766), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n780), .A2(G68), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n788), .A2(G137), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n260), .B1(new_n794), .B2(new_n282), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G150), .B2(new_n790), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n984), .A2(new_n985), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n788), .A2(G317), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n315), .B1(new_n794), .B2(new_n769), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G303), .B2(new_n790), .ZN(new_n992));
  NOR2_X1   g0792(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n993));
  AND2_X1   g0793(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n764), .A2(new_n490), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n763), .A2(KEYINPUT46), .A3(G116), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n990), .A2(new_n992), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n766), .A2(G311), .B1(G97), .B2(new_n770), .ZN(new_n998));
  INV_X1    g0798(.A(new_n526), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n998), .B1(new_n999), .B2(new_n761), .C1(new_n779), .C2(new_n206), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n989), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT47), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n980), .B1(new_n1002), .B2(new_n754), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n812), .B2(new_n949), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n977), .A2(new_n1004), .ZN(G387));
  NAND2_X1  g0805(.A1(new_n689), .A2(new_n753), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n743), .A2(new_n702), .B1(G107), .B2(new_n213), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n239), .A2(new_n475), .ZN(new_n1008));
  AOI211_X1 g0808(.A(G45), .B(new_n701), .C1(G68), .C2(G77), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n278), .A2(G50), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT50), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n746), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1007), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n742), .B1(new_n1013), .B2(new_n756), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n795), .A2(G303), .B1(new_n790), .B2(G317), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n792), .B2(new_n767), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G311), .B2(new_n760), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT114), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT48), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n779), .A2(new_n769), .B1(new_n999), .B2(new_n764), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(KEYINPUT49), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n260), .B1(new_n770), .B2(G116), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(new_n768), .C2(new_n787), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1023), .A2(KEYINPUT49), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n779), .A2(new_n329), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n282), .B2(new_n791), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT113), .Z(new_n1030));
  OAI221_X1 g0830(.A(new_n260), .B1(new_n202), .B2(new_n794), .C1(new_n771), .C2(new_n205), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(KEYINPUT112), .B(G150), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1031), .B1(new_n788), .B2(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n760), .A2(new_n327), .B1(G77), .B2(new_n763), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(new_n982), .C2(new_n767), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n1026), .A2(new_n1027), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1014), .B1(new_n1036), .B2(new_n754), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n971), .A2(new_n976), .B1(new_n1006), .B2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n700), .B(KEYINPUT115), .Z(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n971), .B2(new_n737), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1038), .B1(new_n973), .B2(new_n1040), .ZN(G393));
  INV_X1    g0841(.A(new_n973), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n967), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1043), .A2(new_n974), .A3(new_n1039), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n968), .A2(new_n976), .ZN(new_n1045));
  AND3_X1   g0845(.A1(new_n247), .A2(new_n213), .A3(new_n315), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n755), .B1(new_n205), .B2(new_n213), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n742), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n260), .B(new_n798), .C1(G294), .C2(new_n795), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n760), .A2(G303), .B1(G283), .B2(new_n763), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n490), .B2(new_n779), .C1(new_n792), .C2(new_n787), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n766), .A2(G317), .B1(G311), .B2(new_n790), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT52), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n315), .B(new_n818), .C1(G68), .C2(new_n763), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n780), .A2(G77), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n788), .A2(G143), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n766), .A2(G150), .B1(G159), .B2(new_n790), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT51), .Z(new_n1060));
  AOI22_X1  g0860(.A1(new_n760), .A2(G50), .B1(new_n795), .B2(new_n327), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT116), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n1052), .A2(new_n1054), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1048), .B1(new_n1064), .B2(new_n754), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n942), .B2(new_n812), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1044), .A2(new_n1045), .A3(new_n1066), .ZN(G390));
  NAND4_X1  g0867(.A1(new_n469), .A2(KEYINPUT117), .A3(G330), .A4(new_n919), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT117), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n920), .B2(new_n909), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n907), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n858), .A2(new_n860), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n841), .A2(new_n909), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n919), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n861), .A2(new_n732), .A3(new_n1074), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n683), .B(new_n839), .C1(new_n710), .C2(new_n711), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1078), .A2(new_n840), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n863), .B1(new_n734), .B2(new_n842), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n732), .A2(new_n1074), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1073), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n861), .A2(new_n919), .A3(new_n1074), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1072), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n901), .B1(new_n1081), .B2(new_n1073), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n884), .A2(new_n897), .A3(new_n899), .A4(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n910), .B(new_n901), .C1(new_n1073), .C2(new_n1079), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1090), .A2(new_n1077), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1084), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1088), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1084), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1090), .A2(new_n1077), .A3(new_n1091), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(new_n1087), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1094), .A2(new_n1099), .A3(new_n1039), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n836), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n742), .B1(new_n327), .B2(new_n1101), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n206), .A2(new_n761), .B1(new_n767), .B2(new_n769), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n830), .B(new_n1103), .C1(G87), .C2(new_n763), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n788), .A2(G294), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n315), .B1(new_n791), .B2(new_n490), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G97), .B2(new_n795), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1104), .A2(new_n1056), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n761), .A2(new_n827), .B1(new_n282), .B2(new_n771), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G128), .B2(new_n766), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n788), .A2(G125), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n790), .A2(G132), .ZN(new_n1112));
  XOR2_X1   g0912(.A(KEYINPUT54), .B(G143), .Z(new_n1113));
  AOI21_X1  g0913(.A(new_n315), .B1(new_n795), .B2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n763), .A2(new_n1032), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1117));
  XNOR2_X1  g0917(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n982), .B2(new_n779), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1108), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1102), .B1(new_n1120), .B2(new_n754), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n900), .B2(new_n752), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n1123), .A2(KEYINPUT118), .A3(new_n976), .ZN(new_n1124));
  AOI21_X1  g0924(.A(KEYINPUT118), .B1(new_n1123), .B2(new_n976), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1100), .B(new_n1122), .C1(new_n1124), .C2(new_n1125), .ZN(G378));
  INV_X1    g0926(.A(KEYINPUT122), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n878), .A2(KEYINPUT38), .A3(new_n879), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1128), .B(new_n886), .C1(KEYINPUT38), .C2(new_n893), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n914), .A2(new_n1129), .A3(new_n885), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n915), .A2(new_n916), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n1131), .A3(G330), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n661), .A2(new_n304), .A3(new_n662), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n682), .A2(new_n292), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT55), .Z(new_n1135));
  OR2_X1    g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g0938(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1136), .A2(new_n1139), .A3(new_n1137), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1132), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n917), .A2(G330), .A3(new_n1143), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n903), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n900), .A2(new_n902), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n882), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1145), .A2(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(KEYINPUT57), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1072), .B1(new_n1123), .B2(new_n1087), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1127), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT57), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1154), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1071), .A2(new_n907), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1099), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n903), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n903), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1158), .A2(new_n1163), .A3(KEYINPUT122), .A4(KEYINPUT57), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1153), .A2(new_n1156), .A3(new_n1039), .A4(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n742), .B1(G50), .B2(new_n1101), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1143), .A2(new_n752), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n790), .A2(G128), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n827), .B2(new_n794), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G132), .B2(new_n760), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n766), .A2(G125), .B1(new_n763), .B2(new_n1113), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(new_n826), .C2(new_n779), .ZN(new_n1172));
  OR2_X1    g0972(.A1(new_n1172), .A2(KEYINPUT59), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(KEYINPUT59), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n313), .A2(new_n359), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n771), .A2(new_n982), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n788), .C2(G124), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1173), .A2(new_n1174), .A3(new_n1177), .ZN(new_n1178));
  AOI211_X1 g0978(.A(G41), .B(new_n260), .C1(new_n790), .C2(G107), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n329), .B2(new_n794), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G283), .B2(new_n788), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n760), .A2(G97), .B1(G77), .B2(new_n763), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n771), .A2(new_n201), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G116), .B2(new_n766), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1181), .A2(new_n985), .A3(new_n1182), .A4(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT58), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n282), .B(new_n1175), .C1(new_n260), .C2(G41), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT120), .Z(new_n1190));
  NAND4_X1  g0990(.A1(new_n1178), .A2(new_n1187), .A3(new_n1188), .A4(new_n1190), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1166), .B(new_n1167), .C1(new_n754), .C2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1163), .B2(new_n976), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1165), .A2(new_n1193), .ZN(G375));
  OR2_X1    g0994(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1073), .A2(new_n751), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n742), .B1(G68), .B2(new_n1101), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n766), .A2(G294), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n205), .B2(new_n764), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n981), .B(new_n1199), .C1(G116), .C2(new_n760), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n788), .A2(G303), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n315), .B1(new_n794), .B2(new_n206), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G283), .B2(new_n790), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1200), .A2(new_n1028), .A3(new_n1201), .A4(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n260), .B1(new_n791), .B2(new_n827), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G150), .B2(new_n795), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n788), .A2(G128), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1183), .B1(new_n760), .B2(new_n1113), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n766), .A2(G132), .B1(G159), .B2(new_n763), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n779), .A2(new_n282), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1204), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1197), .B1(new_n1212), .B2(new_n754), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1195), .A2(new_n976), .B1(new_n1196), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n957), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1088), .A2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1157), .A2(new_n1195), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1214), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT123), .Z(G381));
  OR4_X1    g1019(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1220));
  INV_X1    g1020(.A(G378), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1165), .A2(new_n1221), .A3(new_n1193), .ZN(new_n1222));
  OR4_X1    g1022(.A1(G387), .A2(new_n1220), .A3(G381), .A4(new_n1222), .ZN(G407));
  OAI211_X1 g1023(.A(G407), .B(G213), .C1(G343), .C2(new_n1222), .ZN(G409));
  NAND3_X1  g1024(.A1(new_n1165), .A2(G378), .A3(new_n1193), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1158), .A2(new_n1215), .A3(new_n1163), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1193), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1221), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(G213), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(G343), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT125), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT125), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1229), .A2(new_n1235), .A3(new_n1232), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1217), .A2(KEYINPUT60), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1217), .A2(KEYINPUT60), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1237), .A2(new_n1039), .A3(new_n1088), .A4(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1214), .ZN(new_n1240));
  INV_X1    g1040(.A(G384), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1239), .A2(G384), .A3(new_n1214), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT62), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1234), .A2(KEYINPUT126), .A3(new_n1236), .A4(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1231), .A2(G2897), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1232), .A2(KEYINPUT124), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1248), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1248), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1244), .A2(new_n1253), .A3(new_n1250), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1235), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1256));
  AOI211_X1 g1056(.A(KEYINPUT125), .B(new_n1231), .C1(new_n1225), .C2(new_n1228), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1255), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1247), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1246), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1256), .A2(new_n1257), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT126), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1231), .B(new_n1244), .C1(new_n1225), .C2(new_n1228), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1264), .B2(KEYINPUT62), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(KEYINPUT127), .B1(new_n1260), .B2(new_n1266), .ZN(new_n1267));
  XOR2_X1   g1067(.A(G393), .B(G396), .Z(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n977), .A2(G390), .A3(new_n1004), .ZN(new_n1270));
  AOI21_X1  g1070(.A(G390), .B1(new_n977), .B2(new_n1004), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(G390), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G387), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n977), .A2(G390), .A3(new_n1004), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1268), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1272), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT61), .B1(new_n1278), .B2(new_n1255), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1234), .A2(new_n1236), .A3(new_n1246), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1229), .A2(new_n1232), .A3(new_n1249), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT126), .B1(new_n1281), .B2(new_n1245), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT127), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1279), .A2(new_n1283), .A3(new_n1284), .A4(new_n1247), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1267), .A2(new_n1277), .A3(new_n1285), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1255), .A2(new_n1233), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1277), .A2(new_n1287), .A3(KEYINPUT61), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1234), .A2(KEYINPUT63), .A3(new_n1236), .A4(new_n1249), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1288), .B(new_n1289), .C1(KEYINPUT63), .C2(new_n1264), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1286), .A2(new_n1290), .ZN(G405));
  NAND2_X1  g1091(.A1(G375), .A2(new_n1221), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1225), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1293), .B(new_n1249), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n1277), .B(new_n1294), .ZN(G402));
endmodule


