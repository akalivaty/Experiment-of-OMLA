//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n827, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936;
  XOR2_X1   g000(.A(G141gat), .B(G148gat), .Z(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(KEYINPUT2), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n202), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G141gat), .B(G148gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n206), .B(new_n205), .C1(new_n210), .C2(KEYINPUT2), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n213));
  XNOR2_X1  g012(.A(G197gat), .B(G204gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(G211gat), .A2(G218gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT79), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT22), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n216), .B1(new_n215), .B2(new_n217), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n214), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G211gat), .B(G218gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n221), .B(new_n214), .C1(new_n218), .C2(new_n219), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT29), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n213), .B1(new_n225), .B2(KEYINPUT86), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT86), .ZN(new_n227));
  AOI211_X1 g026(.A(new_n227), .B(KEYINPUT29), .C1(new_n223), .C2(new_n224), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n212), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G228gat), .A2(G233gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n223), .A2(new_n224), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT80), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n223), .A2(new_n224), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT80), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n212), .A2(KEYINPUT3), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n233), .B(new_n236), .C1(KEYINPUT29), .C2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n229), .A2(new_n231), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G22gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n212), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n223), .A2(KEYINPUT85), .A3(new_n224), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT29), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT85), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n220), .A2(new_n244), .A3(new_n222), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n241), .B1(new_n246), .B2(new_n213), .ZN(new_n247));
  INV_X1    g046(.A(new_n237), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n234), .B1(new_n248), .B2(new_n243), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n230), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n239), .A2(new_n240), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT87), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G78gat), .B(G106gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT31), .B(G50gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT88), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n250), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G22gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n251), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT88), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n253), .A2(new_n263), .A3(new_n256), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n258), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n263), .B1(new_n253), .B2(new_n256), .ZN(new_n266));
  INV_X1    g065(.A(new_n256), .ZN(new_n267));
  AOI211_X1 g066(.A(KEYINPUT88), .B(new_n267), .C1(new_n251), .C2(new_n252), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n261), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT24), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(G183gat), .A3(G190gat), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n274));
  AND2_X1   g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT64), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT23), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(G169gat), .B2(G176gat), .ZN(new_n279));
  INV_X1    g078(.A(G169gat), .ZN(new_n280));
  INV_X1    g079(.A(G176gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT23), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n273), .B(new_n283), .C1(new_n274), .C2(new_n275), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n277), .A2(new_n279), .A3(new_n282), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n271), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT24), .B1(new_n289), .B2(KEYINPUT67), .ZN(new_n290));
  NAND2_X1  g089(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n291), .A2(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n292));
  OAI22_X1  g091(.A1(new_n290), .A2(new_n292), .B1(G183gat), .B2(G190gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n286), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n296));
  AND4_X1   g095(.A1(new_n279), .A2(new_n282), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n293), .A2(new_n297), .A3(KEYINPUT25), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT68), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n293), .A2(new_n297), .A3(KEYINPUT68), .A4(KEYINPUT25), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n288), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G134gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G127gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G127gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G134gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n303), .A2(KEYINPUT72), .A3(G127gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G113gat), .B(G120gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(KEYINPUT1), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n313));
  INV_X1    g112(.A(G113gat), .ZN(new_n314));
  INV_X1    g113(.A(G120gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT73), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G120gat), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n314), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n314), .A2(KEYINPUT74), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G113gat), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n315), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n313), .B(new_n308), .C1(new_n319), .C2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n304), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n312), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT26), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n286), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT71), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n328), .A2(new_n329), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n275), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT70), .ZN(new_n334));
  OR2_X1    g133(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G190gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT28), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n334), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT69), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n342), .A3(new_n340), .ZN(new_n343));
  AOI21_X1  g142(.A(G190gat), .B1(new_n335), .B2(new_n336), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT69), .B1(new_n344), .B2(KEYINPUT28), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n341), .A2(new_n343), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n333), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n302), .A2(new_n327), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT75), .ZN(new_n350));
  INV_X1    g149(.A(new_n285), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT25), .B1(new_n351), .B2(new_n286), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n300), .A2(new_n301), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n326), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n302), .A2(new_n356), .A3(new_n327), .A4(new_n348), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n350), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G227gat), .A2(G233gat), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT33), .ZN(new_n362));
  XNOR2_X1  g161(.A(G15gat), .B(G43gat), .ZN(new_n363));
  INV_X1    g162(.A(G99gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT76), .B(G71gat), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n365), .B(new_n366), .Z(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n361), .B(KEYINPUT32), .C1(new_n362), .C2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n362), .A2(KEYINPUT32), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n361), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT77), .B1(new_n372), .B2(new_n367), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n370), .B1(new_n358), .B2(new_n360), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n374), .A2(new_n375), .A3(new_n368), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n369), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n358), .A2(new_n360), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT34), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n379), .A2(KEYINPUT78), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(KEYINPUT78), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  OAI211_X1 g181(.A(KEYINPUT78), .B(new_n379), .C1(new_n358), .C2(new_n360), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n377), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n372), .A2(KEYINPUT77), .A3(new_n367), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n375), .B1(new_n374), .B2(new_n368), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n389), .A2(new_n384), .A3(new_n369), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n270), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT35), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n233), .A2(new_n236), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G226gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(new_n354), .B2(new_n243), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n302), .B2(new_n348), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n354), .A2(new_n396), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT29), .B1(new_n302), .B2(new_n348), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n404), .B(new_n234), .C1(new_n396), .C2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n399), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT30), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n354), .A2(new_n243), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n395), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n393), .B1(new_n411), .B2(new_n404), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n397), .A2(new_n398), .A3(new_n232), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n402), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n399), .A2(KEYINPUT30), .A3(new_n406), .A4(new_n403), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n409), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(KEYINPUT83), .B(KEYINPUT5), .Z(new_n417));
  AOI21_X1  g216(.A(new_n213), .B1(new_n209), .B2(new_n211), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n237), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n420), .B(new_n312), .C1(new_n324), .C2(new_n325), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(KEYINPUT73), .B(G120gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT74), .B(G113gat), .ZN(new_n424));
  OAI22_X1  g223(.A1(new_n314), .A2(new_n423), .B1(new_n424), .B2(new_n315), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n425), .A2(new_n313), .A3(new_n308), .A4(new_n304), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n420), .B1(new_n426), .B2(new_n312), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n419), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT4), .B1(new_n326), .B2(new_n212), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n241), .A2(new_n426), .A3(new_n430), .A4(new_n312), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G225gat), .A2(G233gat), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n433), .B(KEYINPUT82), .Z(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n428), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n212), .B1(new_n422), .B2(new_n427), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n326), .A2(new_n212), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n435), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n417), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n428), .A2(new_n432), .A3(new_n435), .ZN(new_n442));
  INV_X1    g241(.A(new_n417), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G1gat), .B(G29gat), .ZN(new_n445));
  INV_X1    g244(.A(G85gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT0), .B(G57gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  NAND3_X1  g248(.A1(new_n441), .A2(new_n444), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n326), .A2(KEYINPUT81), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n241), .B1(new_n452), .B2(new_n421), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n434), .B1(new_n453), .B2(new_n438), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n443), .B1(new_n454), .B2(new_n442), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(new_n421), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n456), .A2(new_n419), .B1(new_n429), .B2(new_n431), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n417), .B1(new_n457), .B2(new_n435), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n451), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n450), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT89), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT89), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n450), .A2(new_n459), .A3(new_n463), .A4(new_n460), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n441), .A2(KEYINPUT6), .A3(new_n444), .A4(new_n449), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT84), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n455), .A2(new_n458), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT6), .A4(new_n449), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT92), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n467), .A2(new_n470), .A3(KEYINPUT92), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n465), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n391), .A2(new_n392), .A3(new_n416), .A4(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n467), .A3(new_n470), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n477), .A2(new_n416), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n265), .A2(new_n269), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n389), .A2(new_n369), .A3(new_n384), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n384), .B1(new_n389), .B2(new_n369), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n478), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n416), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n437), .A2(new_n435), .A3(new_n439), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n486), .B(KEYINPUT39), .C1(new_n457), .C2(new_n435), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n457), .A2(new_n435), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n487), .B(new_n451), .C1(new_n488), .C2(KEYINPUT39), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT40), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n485), .A2(new_n450), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT91), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n397), .A2(new_n398), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(new_n493), .B2(new_n234), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(KEYINPUT90), .A3(new_n393), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n404), .B(new_n393), .C1(new_n396), .C2(new_n405), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(KEYINPUT91), .B(new_n232), .C1(new_n397), .C2(new_n398), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n494), .A2(new_n495), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT37), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT38), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT37), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n399), .A2(new_n503), .A3(new_n406), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n504), .A2(new_n402), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n407), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT37), .B1(new_n412), .B2(new_n413), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(new_n402), .A3(new_n504), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n507), .B1(new_n509), .B2(KEYINPUT38), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n491), .B(new_n479), .C1(new_n475), .C2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n386), .A2(KEYINPUT36), .A3(new_n390), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n480), .B2(new_n481), .ZN(new_n515));
  INV_X1    g314(.A(new_n477), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n270), .B1(new_n516), .B2(new_n485), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n512), .A2(new_n513), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n484), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G15gat), .B(G22gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT16), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n521), .B2(G1gat), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(G1gat), .B2(new_n520), .ZN(new_n523));
  INV_X1    g322(.A(G8gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(G57gat), .B(G64gat), .Z(new_n527));
  INV_X1    g326(.A(KEYINPUT9), .ZN(new_n528));
  INV_X1    g327(.A(G71gat), .ZN(new_n529));
  INV_X1    g328(.A(G78gat), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G71gat), .B(G78gat), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n527), .A2(new_n533), .A3(new_n531), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n537), .B(KEYINPUT100), .Z(new_n538));
  AOI21_X1  g337(.A(new_n526), .B1(new_n538), .B2(KEYINPUT21), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(G183gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT21), .B1(new_n535), .B2(new_n536), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(G211gat), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n542), .B(new_n544), .Z(new_n545));
  XNOR2_X1  g344(.A(G127gat), .B(G155gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n542), .B(new_n544), .ZN(new_n550));
  INV_X1    g349(.A(new_n548), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(G29gat), .A2(G36gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT14), .ZN(new_n555));
  XOR2_X1   g354(.A(KEYINPUT94), .B(G29gat), .Z(new_n556));
  XOR2_X1   g355(.A(KEYINPUT95), .B(G36gat), .Z(new_n557));
  AOI21_X1  g356(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G43gat), .B(G50gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT15), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT96), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n559), .A2(KEYINPUT15), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n558), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT97), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n566), .A2(KEYINPUT97), .A3(new_n567), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G85gat), .A2(G92gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT7), .ZN(new_n574));
  INV_X1    g373(.A(G106gat), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT8), .B1(new_n364), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n574), .B(new_n576), .C1(G85gat), .C2(G92gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(G99gat), .B(G106gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT101), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n572), .B(new_n581), .C1(new_n567), .C2(new_n566), .ZN(new_n582));
  AND2_X1   g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n566), .A2(new_n580), .B1(KEYINPUT41), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G134gat), .B(G162gat), .Z(new_n588));
  NOR2_X1   g387(.A1(new_n583), .A2(KEYINPUT41), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n586), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n582), .A2(new_n584), .A3(new_n591), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n587), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n590), .B1(new_n587), .B2(new_n592), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n553), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G169gat), .B(G197gat), .Z(new_n597));
  XNOR2_X1  g396(.A(G113gat), .B(G141gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n601), .B(KEYINPUT12), .Z(new_n602));
  INV_X1    g401(.A(new_n566), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n526), .B1(new_n603), .B2(KEYINPUT17), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n572), .A2(new_n604), .B1(new_n566), .B2(new_n526), .ZN(new_n605));
  NAND2_X1  g404(.A1(G229gat), .A2(G233gat), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n605), .A2(KEYINPUT98), .A3(KEYINPUT18), .A4(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n571), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT97), .B1(new_n566), .B2(new_n567), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n604), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n566), .A2(new_n526), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n610), .A2(KEYINPUT18), .A3(new_n606), .A4(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT98), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  OR3_X1    g414(.A1(new_n566), .A2(KEYINPUT99), .A3(new_n526), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT99), .B1(new_n566), .B2(new_n526), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n611), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n606), .B(KEYINPUT13), .Z(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n610), .A2(new_n606), .A3(new_n611), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n620), .B1(new_n621), .B2(KEYINPUT18), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n602), .B1(new_n615), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n620), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n606), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT18), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n602), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n627), .A2(new_n614), .A3(new_n607), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n580), .A2(KEYINPUT10), .A3(new_n538), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n579), .B(new_n537), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT102), .ZN(new_n636));
  NAND2_X1  g435(.A1(G230gat), .A2(G233gat), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n631), .A2(new_n638), .A3(new_n634), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G176gat), .B(G204gat), .Z(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n644), .B1(new_n632), .B2(new_n637), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n644), .B(KEYINPUT103), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n635), .A2(new_n637), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n632), .A2(new_n637), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n519), .A2(new_n596), .A3(new_n630), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT104), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n516), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g456(.A1(new_n655), .A2(new_n485), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT16), .B(G8gat), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT42), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n658), .A2(new_n524), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(G1325gat));
  NAND2_X1  g462(.A1(new_n386), .A2(new_n390), .ZN(new_n664));
  AOI21_X1  g463(.A(G15gat), .B1(new_n655), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n515), .A2(new_n513), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n655), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n665), .B1(G15gat), .B2(new_n667), .ZN(G1326gat));
  NAND2_X1  g467(.A1(new_n655), .A2(new_n270), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT43), .B(G22gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  AND3_X1   g470(.A1(new_n515), .A2(new_n513), .A3(new_n517), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n672), .A2(new_n512), .B1(new_n476), .B2(new_n483), .ZN(new_n673));
  INV_X1    g472(.A(new_n595), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT44), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n519), .A2(new_n676), .A3(new_n595), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n630), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n652), .B(KEYINPUT106), .Z(new_n682));
  NAND2_X1  g481(.A1(new_n553), .A2(KEYINPUT105), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n549), .A2(new_n552), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n682), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n556), .B1(new_n688), .B2(new_n477), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n553), .A2(new_n630), .A3(new_n653), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n673), .A2(new_n690), .A3(new_n674), .ZN(new_n691));
  INV_X1    g490(.A(new_n556), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n516), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n689), .A2(new_n694), .ZN(G1328gat));
  OAI21_X1  g494(.A(new_n557), .B1(new_n688), .B2(new_n416), .ZN(new_n696));
  INV_X1    g495(.A(new_n557), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n691), .A2(new_n485), .A3(new_n697), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT46), .Z(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(G1329gat));
  NAND4_X1  g499(.A1(new_n681), .A2(G43gat), .A3(new_n666), .A4(new_n687), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n691), .A2(new_n664), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n702), .A2(G43gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n701), .A2(new_n703), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT47), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n705), .A2(new_n706), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(G1330gat));
  NAND3_X1  g510(.A1(new_n681), .A2(new_n270), .A3(new_n687), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G50gat), .ZN(new_n713));
  INV_X1    g512(.A(G50gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n691), .A2(new_n714), .A3(new_n270), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT111), .Z(new_n716));
  NAND3_X1  g515(.A1(new_n713), .A2(KEYINPUT48), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n715), .B(KEYINPUT110), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(G50gat), .B2(new_n712), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n717), .B1(new_n719), .B2(new_n720), .ZN(G1331gat));
  INV_X1    g520(.A(new_n682), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n673), .A2(new_n722), .A3(new_n630), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n596), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n516), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g526(.A(new_n416), .B(KEYINPUT112), .Z(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  AOI211_X1 g528(.A(new_n729), .B(new_n724), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT113), .B(KEYINPUT114), .Z(new_n731));
  NOR2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n730), .B(new_n733), .ZN(G1333gat));
  NAND3_X1  g533(.A1(new_n725), .A2(new_n529), .A3(new_n664), .ZN(new_n735));
  INV_X1    g534(.A(new_n666), .ZN(new_n736));
  OAI21_X1  g535(.A(G71gat), .B1(new_n724), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n479), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(new_n530), .ZN(G1335gat));
  INV_X1    g540(.A(KEYINPUT116), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n673), .B2(new_n674), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n519), .A2(KEYINPUT116), .A3(new_n595), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n684), .A2(new_n630), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n743), .A2(new_n744), .A3(KEYINPUT51), .A4(new_n745), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n750), .A2(new_n446), .A3(new_n516), .A4(new_n652), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT115), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n745), .A2(new_n652), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n752), .B1(new_n678), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  AOI211_X1 g555(.A(KEYINPUT115), .B(new_n753), .C1(new_n675), .C2(new_n677), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n477), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n751), .B1(new_n759), .B2(new_n446), .ZN(G1336gat));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n485), .B1(new_n755), .B2(new_n757), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G92gat), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n722), .B1(new_n748), .B2(new_n749), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n729), .A2(G92gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n761), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n678), .A2(new_n728), .A3(new_n754), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT52), .B1(new_n768), .B2(G92gat), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT117), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n766), .A2(new_n769), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n762), .A2(G92gat), .B1(new_n764), .B2(new_n765), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n772), .B(new_n773), .C1(new_n774), .C2(new_n761), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n771), .A2(new_n775), .ZN(G1337gat));
  NAND4_X1  g575(.A1(new_n750), .A2(new_n364), .A3(new_n664), .A4(new_n652), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n736), .B1(new_n756), .B2(new_n758), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n364), .ZN(G1338gat));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n575), .A3(new_n270), .ZN(new_n780));
  XOR2_X1   g579(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n781));
  NOR3_X1   g580(.A1(new_n679), .A2(new_n479), .A3(new_n753), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n780), .B(new_n781), .C1(new_n782), .C2(new_n575), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n270), .B1(new_n755), .B2(new_n757), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G106gat), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(new_n780), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(G1339gat));
  INV_X1    g587(.A(new_n391), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n683), .A2(new_n686), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n640), .B(KEYINPUT54), .C1(new_n637), .C2(new_n635), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n644), .B1(new_n649), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT55), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n646), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n791), .A2(KEYINPUT55), .A3(new_n793), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT119), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n791), .A2(new_n793), .A3(new_n798), .A4(KEYINPUT55), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n630), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n605), .A2(new_n606), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n618), .A2(new_n619), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n601), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n629), .A2(new_n652), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n595), .B1(new_n801), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n629), .A2(new_n804), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(new_n595), .A3(new_n795), .A4(new_n800), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n790), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n684), .A2(new_n674), .A3(new_n653), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n630), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n789), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(new_n516), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n729), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n630), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G113gat), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n819), .B1(new_n818), .B2(new_n424), .ZN(G1340gat));
  NAND4_X1  g619(.A1(new_n814), .A2(new_n516), .A3(new_n682), .A4(new_n729), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G120gat), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n653), .A2(new_n423), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n816), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n824), .B(new_n825), .ZN(G1341gat));
  NOR3_X1   g625(.A1(new_n816), .A2(new_n307), .A3(new_n790), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n817), .A2(new_n684), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n827), .B1(new_n307), .B2(new_n828), .ZN(G1342gat));
  NOR2_X1   g628(.A1(new_n674), .A2(new_n485), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n303), .A3(new_n830), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n831), .A2(KEYINPUT56), .ZN(new_n832));
  OAI21_X1  g631(.A(G134gat), .B1(new_n816), .B2(new_n674), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(KEYINPUT56), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(G1343gat));
  NAND2_X1  g634(.A1(new_n801), .A2(new_n805), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n674), .ZN(new_n837));
  AOI22_X1  g636(.A1(new_n837), .A2(new_n808), .B1(new_n683), .B2(new_n686), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n270), .B1(new_n838), .B2(new_n812), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n736), .A2(new_n516), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n839), .A2(new_n728), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(G141gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n842), .A3(new_n630), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n553), .B1(new_n806), .B2(new_n809), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g646(.A(KEYINPUT121), .B(new_n553), .C1(new_n806), .C2(new_n809), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n847), .A2(new_n813), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n844), .B1(new_n849), .B2(new_n270), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n736), .A2(new_n516), .A3(new_n729), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n839), .B2(KEYINPUT57), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n850), .A2(new_n853), .A3(new_n680), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n843), .B1(new_n854), .B2(new_n842), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT58), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n843), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  OAI221_X1 g658(.A(new_n843), .B1(new_n857), .B2(new_n856), .C1(new_n854), .C2(new_n842), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1344gat));
  AOI21_X1  g660(.A(new_n479), .B1(new_n810), .B2(new_n813), .ZN(new_n862));
  INV_X1    g661(.A(G148gat), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n851), .A2(new_n653), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n839), .A2(KEYINPUT57), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n845), .A2(new_n813), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n844), .A3(new_n270), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n864), .A3(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n863), .B1(new_n870), .B2(new_n871), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n866), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n851), .B1(new_n862), .B2(new_n844), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n848), .A2(new_n813), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n479), .B1(new_n876), .B2(new_n847), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n875), .B(new_n652), .C1(new_n877), .C2(new_n844), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n878), .A2(new_n866), .A3(G148gat), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n865), .B1(new_n874), .B2(new_n879), .ZN(G1345gat));
  OAI21_X1  g679(.A(new_n875), .B1(new_n877), .B2(new_n844), .ZN(new_n881));
  OAI21_X1  g680(.A(G155gat), .B1(new_n881), .B2(new_n790), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n841), .A2(new_n203), .A3(new_n684), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1346gat));
  OAI21_X1  g683(.A(G162gat), .B1(new_n881), .B2(new_n674), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n839), .A2(new_n840), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n204), .A3(new_n830), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(G1347gat));
  NOR2_X1   g687(.A1(new_n729), .A2(new_n516), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n814), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n280), .A3(new_n630), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n516), .A2(new_n416), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n814), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G169gat), .B1(new_n893), .B2(new_n680), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n894), .ZN(G1348gat));
  AOI21_X1  g694(.A(G176gat), .B1(new_n890), .B2(new_n652), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n893), .A2(new_n281), .A3(new_n722), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(G1349gat));
  NOR2_X1   g697(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n890), .A2(new_n337), .A3(new_n684), .ZN(new_n900));
  OAI21_X1  g699(.A(G183gat), .B1(new_n893), .B2(new_n790), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AND2_X1   g701(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n902), .B(new_n903), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n893), .B2(new_n674), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT61), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n338), .A3(new_n595), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1351gat));
  NOR3_X1   g707(.A1(new_n666), .A2(new_n729), .A3(new_n516), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n862), .A2(new_n909), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n910), .A2(G197gat), .A3(new_n680), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n666), .A2(new_n516), .A3(new_n416), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n912), .A2(KEYINPUT125), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(KEYINPUT125), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n867), .A2(new_n630), .A3(new_n869), .A4(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n911), .B1(G197gat), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT126), .ZN(G1352gat));
  NOR3_X1   g718(.A1(new_n910), .A2(G204gat), .A3(new_n653), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT62), .ZN(new_n921));
  INV_X1    g720(.A(G204gat), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n867), .A2(new_n869), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n923), .A2(new_n722), .A3(new_n915), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n922), .B2(new_n924), .ZN(G1353gat));
  NAND4_X1  g724(.A1(new_n867), .A2(new_n684), .A3(new_n869), .A4(new_n912), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n926), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT63), .B1(new_n926), .B2(G211gat), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n553), .A2(G211gat), .ZN(new_n929));
  OAI22_X1  g728(.A1(new_n927), .A2(new_n928), .B1(new_n910), .B2(new_n929), .ZN(G1354gat));
  OAI21_X1  g729(.A(KEYINPUT127), .B1(new_n923), .B2(new_n915), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n867), .A2(new_n932), .A3(new_n869), .A4(new_n916), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n931), .A2(new_n933), .A3(new_n595), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G218gat), .ZN(new_n935));
  OR3_X1    g734(.A1(new_n910), .A2(G218gat), .A3(new_n674), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1355gat));
endmodule


