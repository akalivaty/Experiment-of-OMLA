

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n652, n653, n654, n655, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772;

  INV_X1 U373 ( .A(n743), .ZN(n352) );
  INV_X1 U374 ( .A(n743), .ZN(n356) );
  INV_X1 U375 ( .A(n743), .ZN(n360) );
  XNOR2_X1 U376 ( .A(n449), .B(n370), .ZN(n641) );
  XNOR2_X1 U377 ( .A(n757), .B(n536), .ZN(n424) );
  INV_X1 U378 ( .A(n351), .ZN(n736) );
  NAND2_X1 U379 ( .A1(n353), .A2(n352), .ZN(n351) );
  XNOR2_X1 U380 ( .A(n733), .B(n354), .ZN(n353) );
  INV_X1 U381 ( .A(n734), .ZN(n354) );
  INV_X1 U382 ( .A(n355), .ZN(n658) );
  NAND2_X1 U383 ( .A1(n357), .A2(n356), .ZN(n355) );
  XNOR2_X1 U384 ( .A(n654), .B(n358), .ZN(n357) );
  INV_X1 U385 ( .A(n655), .ZN(n358) );
  INV_X1 U386 ( .A(n359), .ZN(n652) );
  NAND2_X1 U387 ( .A1(n361), .A2(n360), .ZN(n359) );
  XNOR2_X1 U388 ( .A(n650), .B(n362), .ZN(n361) );
  INV_X1 U389 ( .A(n489), .ZN(n362) );
  XNOR2_X2 U390 ( .A(n564), .B(n493), .ZN(n757) );
  XOR2_X1 U391 ( .A(KEYINPUT77), .B(KEYINPUT18), .Z(n372) );
  XNOR2_X1 U392 ( .A(G137), .B(G128), .ZN(n517) );
  XNOR2_X1 U393 ( .A(n415), .B(n414), .ZN(n772) );
  XNOR2_X2 U394 ( .A(n578), .B(KEYINPUT22), .ZN(n582) );
  XNOR2_X2 U395 ( .A(n437), .B(KEYINPUT33), .ZN(n721) );
  INV_X4 U396 ( .A(G953), .ZN(n761) );
  AND2_X1 U397 ( .A1(n410), .A2(n409), .ZN(n408) );
  XNOR2_X1 U398 ( .A(n527), .B(n445), .ZN(n609) );
  AND2_X1 U399 ( .A1(n769), .A2(n584), .ZN(n444) );
  NOR2_X1 U400 ( .A1(n455), .A2(n452), .ZN(n451) );
  NOR2_X1 U401 ( .A1(n582), .A2(n456), .ZN(n455) );
  NAND2_X1 U402 ( .A1(n435), .A2(n431), .ZN(n437) );
  XNOR2_X1 U403 ( .A(n366), .B(n388), .ZN(n692) );
  AND2_X1 U404 ( .A1(n433), .A2(n432), .ZN(n431) );
  NAND2_X1 U405 ( .A1(n408), .A2(n406), .ZN(n390) );
  OR2_X2 U406 ( .A1(n609), .A2(n607), .ZN(n705) );
  NAND2_X1 U407 ( .A1(n407), .A2(n373), .ZN(n406) );
  NOR2_X1 U408 ( .A1(n588), .A2(n576), .ZN(n694) );
  BUF_X1 U409 ( .A(n590), .Z(n619) );
  NOR2_X1 U410 ( .A1(n739), .A2(G902), .ZN(n527) );
  XOR2_X1 U411 ( .A(n732), .B(KEYINPUT121), .Z(n734) );
  OR2_X1 U412 ( .A1(n660), .A2(G902), .ZN(n481) );
  XNOR2_X1 U413 ( .A(n523), .B(n522), .ZN(n739) );
  XNOR2_X1 U414 ( .A(n515), .B(n486), .ZN(n516) );
  XNOR2_X1 U415 ( .A(KEYINPUT67), .B(n494), .ZN(n758) );
  XOR2_X1 U416 ( .A(KEYINPUT75), .B(KEYINPUT23), .Z(n514) );
  BUF_X1 U417 ( .A(n769), .Z(n363) );
  BUF_X1 U418 ( .A(n725), .Z(n364) );
  XNOR2_X1 U419 ( .A(n443), .B(n442), .ZN(n769) );
  BUF_X1 U420 ( .A(n579), .Z(n365) );
  INV_X1 U421 ( .A(n407), .ZN(n366) );
  BUF_X1 U422 ( .A(n647), .Z(n367) );
  AND2_X2 U423 ( .A1(n725), .A2(n646), .ZN(n426) );
  XNOR2_X2 U424 ( .A(n532), .B(G134), .ZN(n564) );
  NAND2_X1 U425 ( .A1(n623), .A2(n381), .ZN(n380) );
  XNOR2_X1 U426 ( .A(n389), .B(KEYINPUT47), .ZN(n381) );
  NAND2_X1 U427 ( .A1(n772), .A2(KEYINPUT46), .ZN(n382) );
  NAND2_X1 U428 ( .A1(n387), .A2(n385), .ZN(n384) );
  AND2_X1 U429 ( .A1(n392), .A2(n386), .ZN(n385) );
  XNOR2_X1 U430 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U431 ( .A(KEYINPUT3), .B(KEYINPUT69), .ZN(n490) );
  XOR2_X1 U432 ( .A(G116), .B(G119), .Z(n491) );
  XNOR2_X1 U433 ( .A(n463), .B(G107), .ZN(n567) );
  INV_X1 U434 ( .A(G122), .ZN(n463) );
  XNOR2_X1 U435 ( .A(G137), .B(G131), .ZN(n493) );
  XNOR2_X1 U436 ( .A(G101), .B(n758), .ZN(n536) );
  XNOR2_X1 U437 ( .A(n418), .B(n417), .ZN(n423) );
  INV_X1 U438 ( .A(KEYINPUT48), .ZN(n417) );
  NAND2_X1 U439 ( .A1(n394), .A2(n395), .ZN(n418) );
  AND2_X1 U440 ( .A1(n624), .A2(n636), .ZN(n395) );
  XOR2_X1 U441 ( .A(KEYINPUT86), .B(n530), .Z(n691) );
  INV_X1 U442 ( .A(n637), .ZN(n457) );
  AND2_X1 U443 ( .A1(n694), .A2(n699), .ZN(n577) );
  XNOR2_X1 U444 ( .A(n400), .B(n478), .ZN(n643) );
  NOR2_X1 U445 ( .A1(n635), .A2(n692), .ZN(n400) );
  NOR2_X1 U446 ( .A1(n383), .A2(n379), .ZN(n394) );
  NAND2_X1 U447 ( .A1(n382), .A2(n380), .ZN(n379) );
  XNOR2_X1 U448 ( .A(n465), .B(G104), .ZN(n557) );
  INV_X1 U449 ( .A(G113), .ZN(n465) );
  INV_X1 U450 ( .A(KEYINPUT16), .ZN(n462) );
  NOR2_X1 U451 ( .A1(n692), .A2(n691), .ZN(n689) );
  XNOR2_X1 U452 ( .A(n500), .B(n540), .ZN(n482) );
  XOR2_X1 U453 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n569) );
  XNOR2_X1 U454 ( .A(G116), .B(KEYINPUT102), .ZN(n565) );
  XOR2_X1 U455 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n566) );
  NAND2_X1 U456 ( .A1(n391), .A2(n375), .ZN(n377) );
  XNOR2_X1 U457 ( .A(n466), .B(G110), .ZN(n538) );
  INV_X1 U458 ( .A(KEYINPUT72), .ZN(n466) );
  XNOR2_X1 U459 ( .A(G104), .B(G107), .ZN(n501) );
  NOR2_X1 U460 ( .A1(n620), .A2(n619), .ZN(n633) );
  XNOR2_X1 U461 ( .A(n632), .B(KEYINPUT41), .ZN(n720) );
  NAND2_X1 U462 ( .A1(n689), .A2(n694), .ZN(n632) );
  INV_X1 U463 ( .A(KEYINPUT34), .ZN(n471) );
  NAND2_X1 U464 ( .A1(n402), .A2(n401), .ZN(n635) );
  AND2_X1 U465 ( .A1(n626), .A2(n479), .ZN(n401) );
  XNOR2_X1 U466 ( .A(n516), .B(n556), .ZN(n523) );
  XNOR2_X1 U467 ( .A(G119), .B(G110), .ZN(n520) );
  NOR2_X1 U468 ( .A1(G952), .A2(n761), .ZN(n743) );
  XNOR2_X1 U469 ( .A(n413), .B(KEYINPUT32), .ZN(n584) );
  INV_X1 U470 ( .A(KEYINPUT107), .ZN(n434) );
  INV_X1 U471 ( .A(KEYINPUT44), .ZN(n469) );
  NAND2_X1 U472 ( .A1(n705), .A2(n434), .ZN(n432) );
  OR2_X1 U473 ( .A1(G237), .A2(G902), .ZN(n542) );
  INV_X1 U474 ( .A(KEYINPUT0), .ZN(n422) );
  XNOR2_X1 U475 ( .A(G113), .B(KEYINPUT93), .ZN(n497) );
  XNOR2_X1 U476 ( .A(n448), .B(n447), .ZN(n759) );
  INV_X1 U477 ( .A(G140), .ZN(n447) );
  XNOR2_X1 U478 ( .A(KEYINPUT10), .B(G125), .ZN(n448) );
  NOR2_X1 U479 ( .A1(G953), .A2(G237), .ZN(n495) );
  XNOR2_X1 U480 ( .A(G131), .B(KEYINPUT97), .ZN(n552) );
  XOR2_X1 U481 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n553) );
  XNOR2_X1 U482 ( .A(G143), .B(G122), .ZN(n550) );
  XOR2_X1 U483 ( .A(KEYINPUT99), .B(KEYINPUT12), .Z(n551) );
  XOR2_X1 U484 ( .A(KEYINPUT15), .B(G902), .Z(n644) );
  INV_X1 U485 ( .A(G125), .ZN(n534) );
  NAND2_X1 U486 ( .A1(G234), .A2(G237), .ZN(n544) );
  INV_X1 U487 ( .A(KEYINPUT38), .ZN(n388) );
  INV_X1 U488 ( .A(n627), .ZN(n479) );
  NAND2_X1 U489 ( .A1(n691), .A2(n411), .ZN(n409) );
  XNOR2_X1 U490 ( .A(KEYINPUT1), .B(KEYINPUT66), .ZN(n473) );
  XNOR2_X1 U491 ( .A(n464), .B(n461), .ZN(n539) );
  XNOR2_X1 U492 ( .A(n567), .B(n462), .ZN(n461) );
  XNOR2_X1 U493 ( .A(n538), .B(n557), .ZN(n464) );
  XNOR2_X1 U494 ( .A(G146), .B(n759), .ZN(n556) );
  NAND2_X1 U495 ( .A1(n457), .A2(n459), .ZN(n456) );
  NAND2_X1 U496 ( .A1(n454), .A2(n453), .ZN(n452) );
  NAND2_X1 U497 ( .A1(n637), .A2(KEYINPUT106), .ZN(n454) );
  XNOR2_X1 U498 ( .A(n702), .B(n438), .ZN(n610) );
  INV_X1 U499 ( .A(KEYINPUT6), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n574), .B(n439), .ZN(n732) );
  XNOR2_X1 U501 ( .A(n564), .B(n573), .ZN(n439) );
  XOR2_X1 U502 ( .A(n653), .B(KEYINPUT59), .Z(n655) );
  XNOR2_X1 U503 ( .A(n424), .B(n506), .ZN(n731) );
  NOR2_X1 U504 ( .A1(n727), .A2(n376), .ZN(n728) );
  INV_X1 U505 ( .A(KEYINPUT42), .ZN(n414) );
  INV_X1 U506 ( .A(KEYINPUT40), .ZN(n477) );
  INV_X1 U507 ( .A(KEYINPUT35), .ZN(n442) );
  INV_X1 U508 ( .A(n635), .ZN(n634) );
  INV_X1 U509 ( .A(n389), .ZN(n675) );
  XNOR2_X1 U510 ( .A(n526), .B(n446), .ZN(n445) );
  INV_X1 U511 ( .A(KEYINPUT25), .ZN(n446) );
  NAND2_X1 U512 ( .A1(n398), .A2(n397), .ZN(n396) );
  INV_X1 U513 ( .A(n743), .ZN(n397) );
  XNOR2_X1 U514 ( .A(n399), .B(n661), .ZN(n398) );
  XNOR2_X1 U515 ( .A(n484), .B(n483), .ZN(G75) );
  XNOR2_X1 U516 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n483) );
  OR2_X1 U517 ( .A1(n728), .A2(n485), .ZN(n484) );
  NAND2_X1 U518 ( .A1(n729), .A2(n761), .ZN(n485) );
  INV_X1 U519 ( .A(n584), .ZN(n770) );
  AND2_X2 U520 ( .A1(n378), .A2(n377), .ZN(n737) );
  INV_X1 U521 ( .A(n458), .ZN(n453) );
  INV_X1 U522 ( .A(n702), .ZN(n458) );
  OR2_X1 U523 ( .A1(n548), .A2(n422), .ZN(n368) );
  AND2_X1 U524 ( .A1(n423), .A2(n687), .ZN(n369) );
  XOR2_X1 U525 ( .A(n543), .B(KEYINPUT85), .Z(n370) );
  XOR2_X1 U526 ( .A(n535), .B(n534), .Z(n371) );
  NOR2_X1 U527 ( .A1(n691), .A2(n411), .ZN(n373) );
  AND2_X1 U528 ( .A1(n687), .A2(n686), .ZN(n374) );
  NAND2_X1 U529 ( .A1(n644), .A2(KEYINPUT2), .ZN(n375) );
  INV_X1 U530 ( .A(G472), .ZN(n480) );
  AND2_X1 U531 ( .A1(n378), .A2(G472), .ZN(n659) );
  INV_X1 U532 ( .A(n378), .ZN(n376) );
  XNOR2_X2 U533 ( .A(n425), .B(KEYINPUT74), .ZN(n378) );
  AND2_X1 U534 ( .A1(n659), .A2(n377), .ZN(n399) );
  NAND2_X1 U535 ( .A1(n384), .A2(n393), .ZN(n383) );
  INV_X1 U536 ( .A(KEYINPUT46), .ZN(n386) );
  INV_X1 U537 ( .A(n772), .ZN(n387) );
  NOR2_X1 U538 ( .A1(n390), .A2(n368), .ZN(n419) );
  NAND2_X1 U539 ( .A1(n390), .A2(n422), .ZN(n412) );
  OR2_X1 U540 ( .A1(n621), .A2(n390), .ZN(n389) );
  NAND2_X1 U541 ( .A1(n428), .A2(n427), .ZN(n391) );
  NAND2_X1 U542 ( .A1(n771), .A2(KEYINPUT46), .ZN(n393) );
  INV_X1 U543 ( .A(n771), .ZN(n392) );
  XNOR2_X1 U544 ( .A(n396), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U545 ( .A(n625), .B(KEYINPUT30), .ZN(n402) );
  OR2_X1 U546 ( .A1(n420), .A2(n419), .ZN(n403) );
  OR2_X2 U547 ( .A1(n420), .A2(n419), .ZN(n596) );
  NAND2_X1 U548 ( .A1(n470), .A2(n488), .ZN(n443) );
  INV_X1 U549 ( .A(n724), .ZN(n427) );
  BUF_X1 U550 ( .A(n721), .Z(n404) );
  NAND2_X1 U551 ( .A1(n365), .A2(n609), .ZN(n405) );
  NAND2_X1 U552 ( .A1(n579), .A2(n609), .ZN(n669) );
  XNOR2_X1 U553 ( .A(n424), .B(n482), .ZN(n660) );
  NAND2_X1 U554 ( .A1(n548), .A2(n422), .ZN(n421) );
  INV_X1 U555 ( .A(n641), .ZN(n407) );
  NAND2_X1 U556 ( .A1(n641), .A2(n411), .ZN(n410) );
  INV_X1 U557 ( .A(KEYINPUT19), .ZN(n411) );
  NAND2_X1 U558 ( .A1(n412), .A2(n421), .ZN(n420) );
  NOR2_X1 U559 ( .A1(n436), .A2(n610), .ZN(n435) );
  NAND2_X1 U560 ( .A1(n583), .A2(n610), .ZN(n413) );
  NAND2_X1 U561 ( .A1(n633), .A2(n720), .ZN(n415) );
  XNOR2_X1 U562 ( .A(n602), .B(KEYINPUT83), .ZN(n428) );
  XNOR2_X2 U563 ( .A(n416), .B(n477), .ZN(n771) );
  NAND2_X1 U564 ( .A1(n643), .A2(n678), .ZN(n416) );
  NAND2_X2 U565 ( .A1(n596), .A2(n577), .ZN(n578) );
  NAND2_X1 U566 ( .A1(n423), .A2(n374), .ZN(n724) );
  NAND2_X1 U567 ( .A1(n426), .A2(n369), .ZN(n425) );
  INV_X1 U568 ( .A(n705), .ZN(n430) );
  NOR2_X1 U569 ( .A1(n706), .A2(n429), .ZN(n436) );
  NAND2_X1 U570 ( .A1(n430), .A2(KEYINPUT107), .ZN(n429) );
  NAND2_X1 U571 ( .A1(n706), .A2(n434), .ZN(n433) );
  NOR2_X1 U572 ( .A1(n457), .A2(n705), .ZN(n594) );
  XNOR2_X2 U573 ( .A(n481), .B(n480), .ZN(n702) );
  XNOR2_X1 U574 ( .A(n472), .B(n471), .ZN(n470) );
  XNOR2_X1 U575 ( .A(n568), .B(n569), .ZN(n570) );
  XNOR2_X1 U576 ( .A(n440), .B(n371), .ZN(n537) );
  XNOR2_X1 U577 ( .A(n532), .B(n533), .ZN(n440) );
  XNOR2_X2 U578 ( .A(n441), .B(KEYINPUT65), .ZN(n579) );
  NAND2_X1 U579 ( .A1(n451), .A2(n450), .ZN(n441) );
  XNOR2_X1 U580 ( .A(n460), .B(n469), .ZN(n468) );
  NAND2_X1 U581 ( .A1(n444), .A2(n669), .ZN(n460) );
  OR2_X2 U582 ( .A1(n647), .A2(n644), .ZN(n449) );
  XNOR2_X1 U583 ( .A(n541), .B(n751), .ZN(n647) );
  NOR2_X1 U584 ( .A1(n582), .A2(n637), .ZN(n585) );
  NAND2_X1 U585 ( .A1(n582), .A2(KEYINPUT106), .ZN(n450) );
  INV_X1 U586 ( .A(KEYINPUT106), .ZN(n459) );
  NAND2_X1 U587 ( .A1(n468), .A2(n601), .ZN(n467) );
  XNOR2_X2 U588 ( .A(n467), .B(KEYINPUT45), .ZN(n725) );
  NAND2_X1 U589 ( .A1(n721), .A2(n403), .ZN(n472) );
  XNOR2_X2 U590 ( .A(n590), .B(n473), .ZN(n706) );
  NOR2_X1 U591 ( .A1(n474), .A2(n743), .ZN(G54) );
  XNOR2_X1 U592 ( .A(n476), .B(n475), .ZN(n474) );
  XNOR2_X1 U593 ( .A(n731), .B(n730), .ZN(n475) );
  NAND2_X1 U594 ( .A1(n737), .A2(G469), .ZN(n476) );
  INV_X1 U595 ( .A(KEYINPUT39), .ZN(n478) );
  XOR2_X1 U596 ( .A(n514), .B(n513), .Z(n486) );
  XNOR2_X1 U597 ( .A(KEYINPUT62), .B(KEYINPUT110), .ZN(n487) );
  AND2_X1 U598 ( .A1(n588), .A2(n576), .ZN(n488) );
  XOR2_X1 U599 ( .A(n649), .B(n648), .Z(n489) );
  INV_X1 U600 ( .A(KEYINPUT5), .ZN(n496) );
  XNOR2_X1 U601 ( .A(n497), .B(n496), .ZN(n498) );
  INV_X1 U602 ( .A(KEYINPUT68), .ZN(n507) );
  XNOR2_X1 U603 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U604 ( .A(n660), .B(n487), .ZN(n661) );
  INV_X1 U605 ( .A(KEYINPUT123), .ZN(n738) );
  XNOR2_X1 U606 ( .A(KEYINPUT120), .B(KEYINPUT60), .ZN(n657) );
  XNOR2_X1 U607 ( .A(n491), .B(n490), .ZN(n540) );
  XNOR2_X2 U608 ( .A(G128), .B(KEYINPUT64), .ZN(n492) );
  XNOR2_X2 U609 ( .A(n492), .B(G143), .ZN(n532) );
  XOR2_X1 U610 ( .A(G146), .B(KEYINPUT4), .Z(n494) );
  XOR2_X1 U611 ( .A(KEYINPUT73), .B(n495), .Z(n549) );
  NAND2_X1 U612 ( .A1(n549), .A2(G210), .ZN(n499) );
  XOR2_X1 U613 ( .A(KEYINPUT88), .B(G140), .Z(n502) );
  XNOR2_X1 U614 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U615 ( .A(n538), .B(n503), .Z(n505) );
  NAND2_X1 U616 ( .A1(G227), .A2(n761), .ZN(n504) );
  XNOR2_X1 U617 ( .A(n505), .B(n504), .ZN(n506) );
  NOR2_X2 U618 ( .A1(G902), .A2(n731), .ZN(n510) );
  INV_X1 U619 ( .A(G469), .ZN(n508) );
  XNOR2_X2 U620 ( .A(n510), .B(n509), .ZN(n590) );
  XOR2_X1 U621 ( .A(KEYINPUT82), .B(KEYINPUT8), .Z(n512) );
  NAND2_X1 U622 ( .A1(G234), .A2(n761), .ZN(n511) );
  XNOR2_X1 U623 ( .A(n512), .B(n511), .ZN(n572) );
  NAND2_X1 U624 ( .A1(G221), .A2(n572), .ZN(n515) );
  XNOR2_X1 U625 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n513) );
  XOR2_X1 U626 ( .A(KEYINPUT24), .B(KEYINPUT70), .Z(n518) );
  XNOR2_X1 U627 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U628 ( .A(n519), .B(KEYINPUT91), .Z(n521) );
  XNOR2_X1 U629 ( .A(n521), .B(n520), .ZN(n522) );
  INV_X1 U630 ( .A(n644), .ZN(n524) );
  NAND2_X1 U631 ( .A1(n524), .A2(G234), .ZN(n525) );
  XNOR2_X1 U632 ( .A(n525), .B(KEYINPUT20), .ZN(n528) );
  NAND2_X1 U633 ( .A1(G217), .A2(n528), .ZN(n526) );
  NAND2_X1 U634 ( .A1(G221), .A2(n528), .ZN(n529) );
  XNOR2_X1 U635 ( .A(KEYINPUT21), .B(n529), .ZN(n607) );
  NAND2_X1 U636 ( .A1(n542), .A2(G214), .ZN(n530) );
  XNOR2_X1 U637 ( .A(KEYINPUT17), .B(KEYINPUT76), .ZN(n531) );
  XNOR2_X1 U638 ( .A(n372), .B(n531), .ZN(n533) );
  NAND2_X1 U639 ( .A1(G224), .A2(n761), .ZN(n535) );
  XNOR2_X1 U640 ( .A(n537), .B(n536), .ZN(n541) );
  XNOR2_X1 U641 ( .A(n540), .B(n539), .ZN(n751) );
  NAND2_X1 U642 ( .A1(G210), .A2(n542), .ZN(n543) );
  XOR2_X1 U643 ( .A(KEYINPUT71), .B(KEYINPUT14), .Z(n545) );
  XNOR2_X1 U644 ( .A(n545), .B(n544), .ZN(n546) );
  NAND2_X1 U645 ( .A1(G952), .A2(n546), .ZN(n719) );
  NOR2_X1 U646 ( .A1(G953), .A2(n719), .ZN(n606) );
  NAND2_X1 U647 ( .A1(G902), .A2(n546), .ZN(n603) );
  XNOR2_X1 U648 ( .A(G898), .B(KEYINPUT87), .ZN(n746) );
  NAND2_X1 U649 ( .A1(G953), .A2(n746), .ZN(n753) );
  NOR2_X1 U650 ( .A1(n603), .A2(n753), .ZN(n547) );
  NOR2_X1 U651 ( .A1(n606), .A2(n547), .ZN(n548) );
  XNOR2_X1 U652 ( .A(KEYINPUT13), .B(G475), .ZN(n563) );
  NAND2_X1 U653 ( .A1(G214), .A2(n549), .ZN(n561) );
  XNOR2_X1 U654 ( .A(n551), .B(n550), .ZN(n555) );
  XNOR2_X1 U655 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U656 ( .A(n555), .B(n554), .Z(n559) );
  XNOR2_X1 U657 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U658 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U659 ( .A(n561), .B(n560), .ZN(n653) );
  NOR2_X1 U660 ( .A1(G902), .A2(n653), .ZN(n562) );
  XNOR2_X1 U661 ( .A(n563), .B(n562), .ZN(n588) );
  XNOR2_X1 U662 ( .A(n566), .B(n565), .ZN(n571) );
  XNOR2_X1 U663 ( .A(n567), .B(KEYINPUT103), .ZN(n568) );
  XOR2_X1 U664 ( .A(n571), .B(n570), .Z(n574) );
  NAND2_X1 U665 ( .A1(G217), .A2(n572), .ZN(n573) );
  NOR2_X1 U666 ( .A1(n732), .A2(G902), .ZN(n575) );
  XNOR2_X1 U667 ( .A(n575), .B(G478), .ZN(n589) );
  INV_X1 U668 ( .A(n589), .ZN(n576) );
  INV_X1 U669 ( .A(n607), .ZN(n699) );
  INV_X1 U670 ( .A(n706), .ZN(n637) );
  XOR2_X1 U671 ( .A(KEYINPUT104), .B(n609), .Z(n700) );
  NOR2_X1 U672 ( .A1(n457), .A2(n700), .ZN(n580) );
  XNOR2_X1 U673 ( .A(n580), .B(KEYINPUT105), .ZN(n581) );
  NOR2_X1 U674 ( .A1(n582), .A2(n581), .ZN(n583) );
  INV_X1 U675 ( .A(n610), .ZN(n587) );
  NAND2_X1 U676 ( .A1(n700), .A2(n585), .ZN(n586) );
  NOR2_X1 U677 ( .A1(n587), .A2(n586), .ZN(n662) );
  NOR2_X1 U678 ( .A1(n588), .A2(n589), .ZN(n680) );
  NAND2_X1 U679 ( .A1(n589), .A2(n588), .ZN(n612) );
  INV_X1 U680 ( .A(n612), .ZN(n678) );
  NOR2_X1 U681 ( .A1(n680), .A2(n678), .ZN(n688) );
  XOR2_X1 U682 ( .A(n688), .B(KEYINPUT81), .Z(n622) );
  NOR2_X2 U683 ( .A1(n619), .A2(n705), .ZN(n626) );
  NAND2_X1 U684 ( .A1(n626), .A2(n403), .ZN(n591) );
  XNOR2_X1 U685 ( .A(KEYINPUT92), .B(n591), .ZN(n592) );
  NOR2_X1 U686 ( .A1(n592), .A2(n458), .ZN(n593) );
  XNOR2_X1 U687 ( .A(n593), .B(KEYINPUT94), .ZN(n664) );
  NAND2_X1 U688 ( .A1(n594), .A2(n458), .ZN(n595) );
  XNOR2_X1 U689 ( .A(n595), .B(KEYINPUT95), .ZN(n711) );
  NAND2_X1 U690 ( .A1(n403), .A2(n711), .ZN(n598) );
  XNOR2_X1 U691 ( .A(KEYINPUT96), .B(KEYINPUT31), .ZN(n597) );
  XNOR2_X1 U692 ( .A(n598), .B(n597), .ZN(n681) );
  NOR2_X1 U693 ( .A1(n664), .A2(n681), .ZN(n599) );
  NOR2_X1 U694 ( .A1(n622), .A2(n599), .ZN(n600) );
  NOR2_X1 U695 ( .A1(n662), .A2(n600), .ZN(n601) );
  NAND2_X1 U696 ( .A1(n725), .A2(n644), .ZN(n602) );
  INV_X1 U697 ( .A(n691), .ZN(n614) );
  OR2_X1 U698 ( .A1(n761), .A2(n603), .ZN(n604) );
  NOR2_X1 U699 ( .A1(G900), .A2(n604), .ZN(n605) );
  NOR2_X1 U700 ( .A1(n606), .A2(n605), .ZN(n627) );
  NOR2_X1 U701 ( .A1(n627), .A2(n607), .ZN(n608) );
  NAND2_X1 U702 ( .A1(n609), .A2(n608), .ZN(n617) );
  OR2_X1 U703 ( .A1(n617), .A2(n610), .ZN(n611) );
  NOR2_X1 U704 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U705 ( .A1(n614), .A2(n613), .ZN(n638) );
  NOR2_X1 U706 ( .A1(n366), .A2(n638), .ZN(n615) );
  XNOR2_X1 U707 ( .A(n615), .B(KEYINPUT36), .ZN(n616) );
  NAND2_X1 U708 ( .A1(n616), .A2(n637), .ZN(n683) );
  XNOR2_X1 U709 ( .A(KEYINPUT84), .B(n683), .ZN(n624) );
  NOR2_X1 U710 ( .A1(n453), .A2(n617), .ZN(n618) );
  XOR2_X1 U711 ( .A(n618), .B(KEYINPUT28), .Z(n620) );
  INV_X1 U712 ( .A(n633), .ZN(n621) );
  NAND2_X1 U713 ( .A1(n675), .A2(n622), .ZN(n623) );
  NAND2_X1 U714 ( .A1(KEYINPUT47), .A2(n688), .ZN(n630) );
  NOR2_X1 U715 ( .A1(n691), .A2(n702), .ZN(n625) );
  NAND2_X1 U716 ( .A1(n407), .A2(n634), .ZN(n628) );
  XNOR2_X1 U717 ( .A(KEYINPUT109), .B(n628), .ZN(n629) );
  NAND2_X1 U718 ( .A1(n629), .A2(n488), .ZN(n674) );
  NAND2_X1 U719 ( .A1(n630), .A2(n674), .ZN(n631) );
  XNOR2_X1 U720 ( .A(n631), .B(KEYINPUT79), .ZN(n636) );
  OR2_X1 U721 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U722 ( .A(n639), .B(KEYINPUT108), .ZN(n640) );
  XNOR2_X1 U723 ( .A(n640), .B(KEYINPUT43), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n642), .A2(n366), .ZN(n687) );
  NAND2_X1 U725 ( .A1(n643), .A2(n680), .ZN(n686) );
  NAND2_X1 U726 ( .A1(KEYINPUT2), .A2(n686), .ZN(n645) );
  XOR2_X1 U727 ( .A(KEYINPUT78), .B(n645), .Z(n646) );
  NAND2_X1 U728 ( .A1(n737), .A2(G210), .ZN(n650) );
  XNOR2_X1 U729 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n367), .B(KEYINPUT80), .ZN(n648) );
  XNOR2_X1 U731 ( .A(n652), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U732 ( .A1(n737), .A2(G475), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n658), .B(n657), .ZN(G60) );
  XOR2_X1 U734 ( .A(G101), .B(n662), .Z(G3) );
  NAND2_X1 U735 ( .A1(n664), .A2(n678), .ZN(n663) );
  XNOR2_X1 U736 ( .A(n663), .B(G104), .ZN(G6) );
  XOR2_X1 U737 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n666) );
  NAND2_X1 U738 ( .A1(n680), .A2(n664), .ZN(n665) );
  XNOR2_X1 U739 ( .A(n666), .B(n665), .ZN(n668) );
  XOR2_X1 U740 ( .A(G107), .B(KEYINPUT111), .Z(n667) );
  XNOR2_X1 U741 ( .A(n668), .B(n667), .ZN(G9) );
  XNOR2_X1 U742 ( .A(n405), .B(G110), .ZN(G12) );
  XOR2_X1 U743 ( .A(KEYINPUT29), .B(KEYINPUT112), .Z(n671) );
  NAND2_X1 U744 ( .A1(n675), .A2(n680), .ZN(n670) );
  XNOR2_X1 U745 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U746 ( .A(G128), .B(n672), .ZN(G30) );
  XOR2_X1 U747 ( .A(G143), .B(KEYINPUT113), .Z(n673) );
  XNOR2_X1 U748 ( .A(n674), .B(n673), .ZN(G45) );
  NAND2_X1 U749 ( .A1(n675), .A2(n678), .ZN(n676) );
  XNOR2_X1 U750 ( .A(n676), .B(KEYINPUT114), .ZN(n677) );
  XNOR2_X1 U751 ( .A(G146), .B(n677), .ZN(G48) );
  NAND2_X1 U752 ( .A1(n681), .A2(n678), .ZN(n679) );
  XNOR2_X1 U753 ( .A(n679), .B(G113), .ZN(G15) );
  NAND2_X1 U754 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U755 ( .A(n682), .B(G116), .ZN(G18) );
  XNOR2_X1 U756 ( .A(KEYINPUT37), .B(KEYINPUT115), .ZN(n684) );
  XNOR2_X1 U757 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U758 ( .A(G125), .B(n685), .ZN(G27) );
  XNOR2_X1 U759 ( .A(G134), .B(n686), .ZN(G36) );
  XNOR2_X1 U760 ( .A(G140), .B(n687), .ZN(G42) );
  INV_X1 U761 ( .A(n688), .ZN(n690) );
  NAND2_X1 U762 ( .A1(n690), .A2(n689), .ZN(n697) );
  NAND2_X1 U763 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U764 ( .A(KEYINPUT118), .B(n693), .ZN(n695) );
  NAND2_X1 U765 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U766 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U767 ( .A1(n698), .A2(n404), .ZN(n716) );
  XNOR2_X1 U768 ( .A(KEYINPUT51), .B(KEYINPUT117), .ZN(n713) );
  NOR2_X1 U769 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U770 ( .A(n701), .B(KEYINPUT49), .ZN(n703) );
  NAND2_X1 U771 ( .A1(n703), .A2(n453), .ZN(n704) );
  XNOR2_X1 U772 ( .A(KEYINPUT116), .B(n704), .ZN(n709) );
  NAND2_X1 U773 ( .A1(n457), .A2(n705), .ZN(n707) );
  XOR2_X1 U774 ( .A(KEYINPUT50), .B(n707), .Z(n708) );
  NOR2_X1 U775 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U776 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U777 ( .A(n713), .B(n712), .Z(n714) );
  NAND2_X1 U778 ( .A1(n720), .A2(n714), .ZN(n715) );
  NAND2_X1 U779 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U780 ( .A(KEYINPUT52), .B(n717), .Z(n718) );
  NOR2_X1 U781 ( .A1(n719), .A2(n718), .ZN(n723) );
  AND2_X1 U782 ( .A1(n404), .A2(n720), .ZN(n722) );
  NOR2_X1 U783 ( .A1(n723), .A2(n722), .ZN(n729) );
  INV_X1 U784 ( .A(n364), .ZN(n747) );
  NOR2_X1 U785 ( .A1(n724), .A2(n747), .ZN(n726) );
  NOR2_X1 U786 ( .A1(KEYINPUT2), .A2(n726), .ZN(n727) );
  XOR2_X1 U787 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n730) );
  NAND2_X1 U788 ( .A1(n737), .A2(G478), .ZN(n733) );
  XNOR2_X1 U789 ( .A(n736), .B(KEYINPUT122), .ZN(G63) );
  NAND2_X1 U790 ( .A1(n737), .A2(G217), .ZN(n741) );
  XNOR2_X1 U791 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U792 ( .A(n741), .B(n740), .ZN(n742) );
  NOR2_X1 U793 ( .A1(n743), .A2(n742), .ZN(G66) );
  NAND2_X1 U794 ( .A1(G953), .A2(G224), .ZN(n744) );
  XOR2_X1 U795 ( .A(KEYINPUT61), .B(n744), .Z(n745) );
  NOR2_X1 U796 ( .A1(n746), .A2(n745), .ZN(n750) );
  NOR2_X1 U797 ( .A1(G953), .A2(n747), .ZN(n748) );
  XNOR2_X1 U798 ( .A(n748), .B(KEYINPUT124), .ZN(n749) );
  NOR2_X1 U799 ( .A1(n750), .A2(n749), .ZN(n756) );
  XOR2_X1 U800 ( .A(G101), .B(n751), .Z(n752) );
  NAND2_X1 U801 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U802 ( .A(KEYINPUT125), .B(n754), .Z(n755) );
  XNOR2_X1 U803 ( .A(n756), .B(n755), .ZN(G69) );
  XNOR2_X1 U804 ( .A(n757), .B(n758), .ZN(n760) );
  XNOR2_X1 U805 ( .A(n760), .B(n759), .ZN(n763) );
  XNOR2_X1 U806 ( .A(n763), .B(n724), .ZN(n762) );
  NAND2_X1 U807 ( .A1(n762), .A2(n761), .ZN(n768) );
  XNOR2_X1 U808 ( .A(G227), .B(n763), .ZN(n764) );
  NAND2_X1 U809 ( .A1(n764), .A2(G900), .ZN(n765) );
  XNOR2_X1 U810 ( .A(KEYINPUT126), .B(n765), .ZN(n766) );
  NAND2_X1 U811 ( .A1(n766), .A2(G953), .ZN(n767) );
  NAND2_X1 U812 ( .A1(n768), .A2(n767), .ZN(G72) );
  XNOR2_X1 U813 ( .A(n363), .B(G122), .ZN(G24) );
  XOR2_X1 U814 ( .A(G119), .B(n770), .Z(G21) );
  XOR2_X1 U815 ( .A(n771), .B(G131), .Z(G33) );
  XOR2_X1 U816 ( .A(G137), .B(n772), .Z(G39) );
endmodule

