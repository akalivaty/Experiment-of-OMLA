

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587;

  XOR2_X2 U322 ( .A(n454), .B(n368), .Z(n458) );
  XNOR2_X1 U323 ( .A(KEYINPUT54), .B(KEYINPUT123), .ZN(n417) );
  XNOR2_X1 U324 ( .A(KEYINPUT55), .B(n290), .ZN(n464) );
  AND2_X1 U325 ( .A1(n463), .A2(n480), .ZN(n290) );
  XNOR2_X1 U326 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U327 ( .A(KEYINPUT125), .B(n457), .ZN(n584) );
  XNOR2_X1 U328 ( .A(KEYINPUT116), .B(KEYINPUT47), .ZN(n392) );
  INV_X1 U329 ( .A(G204GAT), .ZN(n459) );
  XOR2_X1 U330 ( .A(n437), .B(n436), .Z(n543) );
  XNOR2_X1 U331 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U332 ( .A(n462), .B(n461), .ZN(G1353GAT) );
  XOR2_X1 U333 ( .A(G155GAT), .B(G148GAT), .Z(n292) );
  XNOR2_X1 U334 ( .A(G1GAT), .B(G120GAT), .ZN(n291) );
  XNOR2_X1 U335 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U336 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n294) );
  XNOR2_X1 U337 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U339 ( .A(n296), .B(n295), .Z(n303) );
  XOR2_X1 U340 ( .A(G85GAT), .B(G162GAT), .Z(n300) );
  XOR2_X1 U341 ( .A(KEYINPUT2), .B(KEYINPUT85), .Z(n298) );
  XNOR2_X1 U342 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n441) );
  XNOR2_X1 U344 ( .A(G29GAT), .B(n441), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U346 ( .A(G127GAT), .B(n301), .ZN(n302) );
  XNOR2_X1 U347 ( .A(n303), .B(n302), .ZN(n313) );
  XOR2_X1 U348 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n305) );
  XNOR2_X1 U349 ( .A(KEYINPUT4), .B(KEYINPUT89), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n311) );
  XOR2_X1 U351 ( .A(KEYINPUT0), .B(KEYINPUT80), .Z(n307) );
  XNOR2_X1 U352 ( .A(G113GAT), .B(G134GAT), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n426) );
  XOR2_X1 U354 ( .A(n426), .B(KEYINPUT90), .Z(n309) );
  NAND2_X1 U355 ( .A1(G225GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U357 ( .A(n311), .B(n310), .Z(n312) );
  XOR2_X1 U358 ( .A(n313), .B(n312), .Z(n476) );
  INV_X1 U359 ( .A(n476), .ZN(n529) );
  XOR2_X1 U360 ( .A(G92GAT), .B(G218GAT), .Z(n315) );
  XNOR2_X1 U361 ( .A(G134GAT), .B(G106GAT), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U363 ( .A(KEYINPUT9), .B(KEYINPUT75), .Z(n317) );
  XNOR2_X1 U364 ( .A(KEYINPUT10), .B(KEYINPUT64), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U366 ( .A(n319), .B(n318), .Z(n324) );
  XOR2_X1 U367 ( .A(KEYINPUT65), .B(KEYINPUT11), .Z(n321) );
  NAND2_X1 U368 ( .A1(G232GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U370 ( .A(KEYINPUT76), .B(n322), .ZN(n323) );
  XNOR2_X1 U371 ( .A(n324), .B(n323), .ZN(n332) );
  XNOR2_X1 U372 ( .A(G99GAT), .B(G85GAT), .ZN(n325) );
  XNOR2_X1 U373 ( .A(n325), .B(KEYINPUT72), .ZN(n365) );
  XOR2_X1 U374 ( .A(G36GAT), .B(G190GAT), .Z(n412) );
  XOR2_X1 U375 ( .A(n365), .B(n412), .Z(n330) );
  XOR2_X1 U376 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n327) );
  XNOR2_X1 U377 ( .A(G43GAT), .B(G29GAT), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U379 ( .A(KEYINPUT7), .B(n328), .Z(n345) );
  XOR2_X1 U380 ( .A(G50GAT), .B(G162GAT), .Z(n450) );
  XNOR2_X1 U381 ( .A(n345), .B(n450), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U383 ( .A(n332), .B(n331), .Z(n567) );
  XOR2_X1 U384 ( .A(G113GAT), .B(G15GAT), .Z(n334) );
  XOR2_X1 U385 ( .A(KEYINPUT69), .B(G1GAT), .Z(n378) );
  XOR2_X1 U386 ( .A(G169GAT), .B(G8GAT), .Z(n413) );
  XNOR2_X1 U387 ( .A(n378), .B(n413), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U389 ( .A(n335), .B(G50GAT), .Z(n340) );
  XOR2_X1 U390 ( .A(KEYINPUT66), .B(G141GAT), .Z(n337) );
  XNOR2_X1 U391 ( .A(G197GAT), .B(G22GAT), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n338), .B(G36GAT), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U395 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n342) );
  NAND2_X1 U396 ( .A1(G229GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U398 ( .A(n344), .B(n343), .Z(n347) );
  XNOR2_X1 U399 ( .A(n345), .B(KEYINPUT67), .ZN(n346) );
  XOR2_X1 U400 ( .A(n347), .B(n346), .Z(n515) );
  INV_X1 U401 ( .A(n515), .ZN(n577) );
  XOR2_X1 U402 ( .A(G148GAT), .B(G106GAT), .Z(n349) );
  XNOR2_X1 U403 ( .A(KEYINPUT71), .B(G78GAT), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U405 ( .A(KEYINPUT70), .B(n350), .Z(n454) );
  XOR2_X1 U406 ( .A(G64GAT), .B(KEYINPUT74), .Z(n352) );
  XNOR2_X1 U407 ( .A(G176GAT), .B(G92GAT), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U409 ( .A(G204GAT), .B(n353), .Z(n411) );
  INV_X1 U410 ( .A(n411), .ZN(n357) );
  XOR2_X1 U411 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n355) );
  XOR2_X1 U412 ( .A(G120GAT), .B(G71GAT), .Z(n422) );
  XOR2_X1 U413 ( .A(KEYINPUT13), .B(G57GAT), .Z(n371) );
  XNOR2_X1 U414 ( .A(n422), .B(n371), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n358) );
  INV_X1 U416 ( .A(n358), .ZN(n356) );
  NAND2_X1 U417 ( .A1(n357), .A2(n356), .ZN(n360) );
  NAND2_X1 U418 ( .A1(n411), .A2(n358), .ZN(n359) );
  NAND2_X1 U419 ( .A1(n360), .A2(n359), .ZN(n364) );
  AND2_X1 U420 ( .A1(G230GAT), .A2(G233GAT), .ZN(n362) );
  INV_X1 U421 ( .A(KEYINPUT33), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n365), .B(KEYINPUT73), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U425 ( .A(KEYINPUT41), .B(n458), .Z(n514) );
  AND2_X1 U426 ( .A1(n577), .A2(n514), .ZN(n370) );
  INV_X1 U427 ( .A(KEYINPUT46), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n389) );
  XOR2_X1 U429 ( .A(G22GAT), .B(G155GAT), .Z(n449) );
  XOR2_X1 U430 ( .A(n371), .B(n449), .Z(n373) );
  XNOR2_X1 U431 ( .A(G183GAT), .B(G71GAT), .ZN(n372) );
  XNOR2_X1 U432 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U433 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n375) );
  NAND2_X1 U434 ( .A1(G231GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U436 ( .A(n377), .B(n376), .Z(n380) );
  XOR2_X1 U437 ( .A(G15GAT), .B(G127GAT), .Z(n423) );
  XNOR2_X1 U438 ( .A(n378), .B(n423), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n388) );
  XOR2_X1 U440 ( .A(G64GAT), .B(G211GAT), .Z(n382) );
  XNOR2_X1 U441 ( .A(G8GAT), .B(G78GAT), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U443 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n384) );
  XNOR2_X1 U444 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U446 ( .A(n386), .B(n385), .Z(n387) );
  XOR2_X1 U447 ( .A(n388), .B(n387), .Z(n485) );
  AND2_X1 U448 ( .A1(n389), .A2(n485), .ZN(n390) );
  XNOR2_X1 U449 ( .A(n390), .B(KEYINPUT115), .ZN(n391) );
  NOR2_X1 U450 ( .A1(n567), .A2(n391), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n399) );
  INV_X1 U452 ( .A(n458), .ZN(n470) );
  XOR2_X1 U453 ( .A(KEYINPUT45), .B(KEYINPUT117), .Z(n395) );
  INV_X1 U454 ( .A(n485), .ZN(n582) );
  XNOR2_X1 U455 ( .A(KEYINPUT36), .B(n567), .ZN(n585) );
  NAND2_X1 U456 ( .A1(n582), .A2(n585), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n395), .B(n394), .ZN(n396) );
  NOR2_X1 U458 ( .A1(n396), .A2(n577), .ZN(n397) );
  NAND2_X1 U459 ( .A1(n470), .A2(n397), .ZN(n398) );
  NAND2_X1 U460 ( .A1(n399), .A2(n398), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n400), .B(KEYINPUT48), .ZN(n559) );
  INV_X1 U462 ( .A(n559), .ZN(n545) );
  XOR2_X1 U463 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n402) );
  NAND2_X1 U464 ( .A1(G226GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U465 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U466 ( .A(n403), .B(KEYINPUT93), .Z(n409) );
  XOR2_X1 U467 ( .A(G183GAT), .B(KEYINPUT17), .Z(n405) );
  XNOR2_X1 U468 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n427) );
  XOR2_X1 U470 ( .A(G211GAT), .B(KEYINPUT21), .Z(n407) );
  XNOR2_X1 U471 ( .A(G197GAT), .B(G218GAT), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n442) );
  XNOR2_X1 U473 ( .A(n427), .B(n442), .ZN(n408) );
  XNOR2_X1 U474 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U475 ( .A(n411), .B(n410), .Z(n415) );
  XNOR2_X1 U476 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U477 ( .A(n415), .B(n414), .Z(n532) );
  XOR2_X1 U478 ( .A(n532), .B(KEYINPUT122), .Z(n416) );
  NOR2_X1 U479 ( .A1(n545), .A2(n416), .ZN(n418) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  NOR2_X1 U481 ( .A1(n529), .A2(n419), .ZN(n463) );
  XOR2_X1 U482 ( .A(KEYINPUT84), .B(KEYINPUT82), .Z(n421) );
  XNOR2_X1 U483 ( .A(G169GAT), .B(G43GAT), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n437) );
  XOR2_X1 U485 ( .A(G99GAT), .B(G190GAT), .Z(n425) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U489 ( .A(KEYINPUT20), .B(KEYINPUT81), .Z(n429) );
  XNOR2_X1 U490 ( .A(KEYINPUT83), .B(G176GAT), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U493 ( .A(n433), .B(n432), .Z(n435) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U495 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U496 ( .A(KEYINPUT24), .B(KEYINPUT86), .Z(n439) );
  NAND2_X1 U497 ( .A1(G228GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U499 ( .A(n440), .B(KEYINPUT87), .Z(n444) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U502 ( .A(G204GAT), .B(KEYINPUT88), .Z(n446) );
  XNOR2_X1 U503 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U505 ( .A(n448), .B(n447), .Z(n452) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n454), .B(n453), .ZN(n480) );
  NOR2_X1 U509 ( .A1(n543), .A2(n480), .ZN(n456) );
  XNOR2_X1 U510 ( .A(KEYINPUT26), .B(KEYINPUT98), .ZN(n455) );
  XNOR2_X1 U511 ( .A(n456), .B(n455), .ZN(n558) );
  NAND2_X1 U512 ( .A1(n463), .A2(n558), .ZN(n457) );
  NAND2_X1 U513 ( .A1(n584), .A2(n458), .ZN(n462) );
  XOR2_X1 U514 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n460) );
  INV_X1 U515 ( .A(G190GAT), .ZN(n469) );
  INV_X1 U516 ( .A(n543), .ZN(n465) );
  NOR2_X2 U517 ( .A1(n465), .A2(n464), .ZN(n575) );
  NAND2_X1 U518 ( .A1(n575), .A2(n567), .ZN(n467) );
  XOR2_X1 U519 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n466) );
  XNOR2_X1 U520 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U521 ( .A(n469), .B(n468), .ZN(G1351GAT) );
  XOR2_X1 U522 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n490) );
  NAND2_X1 U523 ( .A1(n577), .A2(n470), .ZN(n503) );
  NAND2_X1 U524 ( .A1(n532), .A2(n543), .ZN(n471) );
  NAND2_X1 U525 ( .A1(n471), .A2(n480), .ZN(n472) );
  XNOR2_X1 U526 ( .A(n472), .B(KEYINPUT99), .ZN(n473) );
  XNOR2_X1 U527 ( .A(n473), .B(KEYINPUT25), .ZN(n475) );
  XNOR2_X1 U528 ( .A(n532), .B(KEYINPUT27), .ZN(n479) );
  NAND2_X1 U529 ( .A1(n558), .A2(n479), .ZN(n474) );
  NAND2_X1 U530 ( .A1(n475), .A2(n474), .ZN(n477) );
  NAND2_X1 U531 ( .A1(n477), .A2(n476), .ZN(n478) );
  XOR2_X1 U532 ( .A(KEYINPUT100), .B(n478), .Z(n484) );
  NAND2_X1 U533 ( .A1(n479), .A2(n529), .ZN(n561) );
  XOR2_X1 U534 ( .A(KEYINPUT28), .B(n480), .Z(n536) );
  NOR2_X1 U535 ( .A1(n561), .A2(n536), .ZN(n542) );
  XOR2_X1 U536 ( .A(n542), .B(KEYINPUT96), .Z(n481) );
  NOR2_X1 U537 ( .A1(n543), .A2(n481), .ZN(n482) );
  XOR2_X1 U538 ( .A(KEYINPUT97), .B(n482), .Z(n483) );
  NOR2_X1 U539 ( .A1(n484), .A2(n483), .ZN(n499) );
  NOR2_X1 U540 ( .A1(n567), .A2(n485), .ZN(n486) );
  XOR2_X1 U541 ( .A(KEYINPUT16), .B(n486), .Z(n487) );
  NOR2_X1 U542 ( .A1(n499), .A2(n487), .ZN(n488) );
  XNOR2_X1 U543 ( .A(KEYINPUT101), .B(n488), .ZN(n517) );
  NOR2_X1 U544 ( .A1(n503), .A2(n517), .ZN(n496) );
  NAND2_X1 U545 ( .A1(n496), .A2(n529), .ZN(n489) );
  XNOR2_X1 U546 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U547 ( .A(G1GAT), .B(n491), .Z(G1324GAT) );
  XOR2_X1 U548 ( .A(G8GAT), .B(KEYINPUT103), .Z(n493) );
  NAND2_X1 U549 ( .A1(n496), .A2(n532), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n493), .B(n492), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(G15GAT), .B(KEYINPUT35), .Z(n495) );
  NAND2_X1 U552 ( .A1(n496), .A2(n543), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NAND2_X1 U554 ( .A1(n536), .A2(n496), .ZN(n497) );
  XNOR2_X1 U555 ( .A(n497), .B(KEYINPUT104), .ZN(n498) );
  XNOR2_X1 U556 ( .A(G22GAT), .B(n498), .ZN(G1327GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT37), .B(KEYINPUT106), .Z(n502) );
  NOR2_X1 U558 ( .A1(n499), .A2(n582), .ZN(n500) );
  NAND2_X1 U559 ( .A1(n500), .A2(n585), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n502), .B(n501), .ZN(n528) );
  NOR2_X1 U561 ( .A1(n503), .A2(n528), .ZN(n504) );
  XNOR2_X1 U562 ( .A(n504), .B(KEYINPUT38), .ZN(n512) );
  NAND2_X1 U563 ( .A1(n512), .A2(n529), .ZN(n507) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n505), .B(KEYINPUT39), .ZN(n506) );
  XNOR2_X1 U566 ( .A(n507), .B(n506), .ZN(G1328GAT) );
  NAND2_X1 U567 ( .A1(n512), .A2(n532), .ZN(n508) );
  XNOR2_X1 U568 ( .A(n508), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n510) );
  NAND2_X1 U570 ( .A1(n543), .A2(n512), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n511), .ZN(G1330GAT) );
  NAND2_X1 U573 ( .A1(n512), .A2(n536), .ZN(n513) );
  XNOR2_X1 U574 ( .A(n513), .B(G50GAT), .ZN(G1331GAT) );
  BUF_X1 U575 ( .A(n514), .Z(n571) );
  NAND2_X1 U576 ( .A1(n515), .A2(n571), .ZN(n516) );
  XNOR2_X1 U577 ( .A(n516), .B(KEYINPUT108), .ZN(n527) );
  NOR2_X1 U578 ( .A1(n527), .A2(n517), .ZN(n523) );
  NAND2_X1 U579 ( .A1(n529), .A2(n523), .ZN(n518) );
  XNOR2_X1 U580 ( .A(n518), .B(KEYINPUT42), .ZN(n519) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(n519), .ZN(G1332GAT) );
  NAND2_X1 U582 ( .A1(n532), .A2(n523), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n520), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U584 ( .A(G71GAT), .B(KEYINPUT109), .Z(n522) );
  NAND2_X1 U585 ( .A1(n523), .A2(n543), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(G1334GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n525) );
  NAND2_X1 U588 ( .A1(n523), .A2(n536), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(G78GAT), .B(n526), .ZN(G1335GAT) );
  XOR2_X1 U591 ( .A(G85GAT), .B(KEYINPUT111), .Z(n531) );
  NOR2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n537), .A2(n529), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n531), .B(n530), .ZN(G1336GAT) );
  NAND2_X1 U595 ( .A1(n532), .A2(n537), .ZN(n533) );
  XNOR2_X1 U596 ( .A(n533), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U597 ( .A1(n537), .A2(n543), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n534), .B(KEYINPUT112), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G99GAT), .B(n535), .ZN(G1338GAT) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(KEYINPUT113), .ZN(n541) );
  XOR2_X1 U601 ( .A(KEYINPUT114), .B(KEYINPUT44), .Z(n539) );
  NAND2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n541), .B(n540), .ZN(G1339GAT) );
  NAND2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U607 ( .A(KEYINPUT118), .B(n546), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n554), .A2(n577), .ZN(n547) );
  XNOR2_X1 U609 ( .A(n547), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT49), .B(KEYINPUT120), .Z(n549) );
  NAND2_X1 U611 ( .A1(n571), .A2(n554), .ZN(n548) );
  XNOR2_X1 U612 ( .A(n549), .B(n548), .ZN(n551) );
  XOR2_X1 U613 ( .A(G120GAT), .B(KEYINPUT119), .Z(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(G1341GAT) );
  NAND2_X1 U615 ( .A1(n554), .A2(n582), .ZN(n552) );
  XNOR2_X1 U616 ( .A(n552), .B(KEYINPUT50), .ZN(n553) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n553), .ZN(G1342GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT51), .B(KEYINPUT121), .Z(n556) );
  NAND2_X1 U619 ( .A1(n567), .A2(n554), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U621 ( .A(G134GAT), .B(n557), .Z(G1343GAT) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U623 ( .A1(n561), .A2(n560), .ZN(n568) );
  NAND2_X1 U624 ( .A1(n577), .A2(n568), .ZN(n562) );
  XNOR2_X1 U625 ( .A(G141GAT), .B(n562), .ZN(G1344GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n564) );
  NAND2_X1 U627 ( .A1(n568), .A2(n571), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(n565), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n582), .A2(n568), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U633 ( .A(n569), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U634 ( .A1(n577), .A2(n575), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G169GAT), .B(n570), .ZN(G1348GAT) );
  NAND2_X1 U636 ( .A1(n575), .A2(n571), .ZN(n573) );
  XOR2_X1 U637 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G176GAT), .ZN(G1349GAT) );
  NAND2_X1 U640 ( .A1(n582), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U642 ( .A1(n584), .A2(n577), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  NAND2_X1 U647 ( .A1(n582), .A2(n584), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(n586), .B(KEYINPUT62), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

