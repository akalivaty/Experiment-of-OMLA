//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(G148gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G141gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n203), .A2(G141gat), .ZN(new_n206));
  NOR3_X1   g005(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  OAI22_X1  g008(.A1(new_n205), .A2(new_n206), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G141gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G148gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT76), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT2), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n204), .A2(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(new_n208), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n210), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G197gat), .B(G204gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT22), .ZN(new_n222));
  INV_X1    g021(.A(G211gat), .ZN(new_n223));
  INV_X1    g022(.A(G218gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G211gat), .B(G218gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n221), .A3(new_n225), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT29), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n220), .B1(new_n231), .B2(KEYINPUT3), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT81), .ZN(new_n233));
  XNOR2_X1  g032(.A(G141gat), .B(G148gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n208), .B(new_n218), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n237), .A3(new_n210), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n229), .A2(new_n230), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n240), .A2(new_n242), .B1(G228gat), .B2(G233gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT81), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n244), .B(new_n220), .C1(new_n231), .C2(KEYINPUT3), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n233), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G228gat), .A2(G233gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT73), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n241), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n229), .A2(KEYINPUT73), .A3(new_n230), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n240), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n248), .B1(new_n252), .B2(new_n232), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n247), .A2(G50gat), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G50gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n253), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(new_n246), .ZN(new_n257));
  NOR3_X1   g056(.A1(new_n254), .A2(new_n257), .A3(KEYINPUT31), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT31), .ZN(new_n259));
  OAI21_X1  g058(.A(G50gat), .B1(new_n247), .B2(new_n253), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n256), .A2(new_n255), .A3(new_n246), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G78gat), .B(G106gat), .Z(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(G22gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT80), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n258), .A2(new_n262), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT31), .B1(new_n254), .B2(new_n257), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n260), .A2(new_n259), .A3(new_n261), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n265), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n272), .B1(new_n273), .B2(KEYINPUT23), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT23), .ZN(new_n275));
  NOR3_X1   g074(.A1(new_n275), .A2(G169gat), .A3(G176gat), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT64), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT25), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AND3_X1   g080(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n277), .A2(new_n278), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n278), .B1(new_n277), .B2(new_n284), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT65), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT64), .ZN(new_n288));
  AND2_X1   g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  INV_X1    g088(.A(G169gat), .ZN(new_n290));
  INV_X1    g089(.A(G176gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n289), .B1(new_n292), .B2(new_n275), .ZN(new_n293));
  INV_X1    g092(.A(new_n276), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n288), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n282), .A2(new_n279), .A3(new_n280), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT25), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT65), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n277), .A2(new_n278), .A3(new_n284), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G183gat), .ZN(new_n301));
  INV_X1    g100(.A(G190gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT26), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n272), .B1(new_n273), .B2(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(KEYINPUT67), .A2(KEYINPUT26), .ZN(new_n306));
  NOR2_X1   g105(.A1(KEYINPUT67), .A2(KEYINPUT26), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n273), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n305), .B1(new_n308), .B2(KEYINPUT68), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT68), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n310), .B(new_n273), .C1(new_n306), .C2(new_n307), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n303), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT27), .B(G183gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n302), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT66), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT66), .ZN(new_n316));
  AND2_X1   g115(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n316), .B(new_n302), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(KEYINPUT28), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n316), .B1(new_n313), .B2(new_n302), .ZN(new_n322));
  INV_X1    g121(.A(new_n319), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n312), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n287), .A2(new_n300), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G134gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G127gat), .ZN(new_n328));
  INV_X1    g127(.A(G127gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G134gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT1), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G120gat), .ZN(new_n333));
  OR2_X1    g132(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G113gat), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT70), .B1(new_n337), .B2(G120gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT70), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(new_n333), .A3(G113gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n332), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n337), .A2(G120gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n333), .A2(G113gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n331), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT69), .B1(new_n329), .B2(G134gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT69), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(new_n327), .A3(G127gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n348), .A3(new_n330), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n342), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n326), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G227gat), .ZN(new_n353));
  INV_X1    g152(.A(G233gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n351), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n287), .A2(new_n300), .A3(new_n325), .A4(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n352), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT34), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT32), .ZN(new_n362));
  XNOR2_X1  g161(.A(G15gat), .B(G43gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(G71gat), .B(G99gat), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n363), .B(new_n364), .Z(new_n365));
  NAND2_X1  g164(.A1(new_n352), .A2(new_n358), .ZN(new_n366));
  AOI221_X4 g165(.A(new_n362), .B1(KEYINPUT33), .B2(new_n365), .C1(new_n366), .C2(new_n355), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n356), .B1(new_n352), .B2(new_n358), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n365), .B1(new_n368), .B2(KEYINPUT33), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n362), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n361), .B(KEYINPUT72), .C1(new_n367), .C2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT72), .B1(new_n371), .B2(new_n367), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n360), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n271), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n312), .A2(new_n320), .A3(new_n324), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n297), .A2(new_n299), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n239), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT74), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n326), .A2(new_n380), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n241), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT75), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n382), .A2(KEYINPUT75), .A3(new_n241), .A4(new_n383), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n250), .A2(new_n251), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n380), .B1(new_n326), .B2(new_n239), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n285), .A2(new_n286), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n381), .B1(new_n391), .B2(new_n325), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n389), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n386), .A2(new_n387), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G8gat), .B(G36gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(G64gat), .B(G92gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n397), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n386), .A2(new_n399), .A3(new_n387), .A4(new_n393), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(KEYINPUT30), .A3(new_n400), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n390), .A2(new_n392), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n402), .A2(new_n389), .B1(new_n384), .B2(new_n385), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT30), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n403), .A2(new_n404), .A3(new_n399), .A4(new_n387), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n238), .A2(new_n351), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT77), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n204), .A2(new_n212), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n214), .A2(new_n216), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n219), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n207), .A2(new_n209), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(new_n234), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n407), .B1(new_n413), .B2(new_n237), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n220), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n406), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G225gat), .A2(G233gat), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n413), .A2(new_n418), .A3(new_n350), .A4(new_n342), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT4), .B1(new_n351), .B2(new_n220), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n416), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n417), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n351), .A2(new_n220), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n350), .A2(new_n342), .B1(new_n236), .B2(new_n210), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT5), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT78), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT5), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n422), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n427), .B1(new_n422), .B2(new_n429), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(G57gat), .B(G85gat), .Z(new_n433));
  XNOR2_X1  g232(.A(G1gat), .B(G29gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n432), .A2(KEYINPUT6), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n437), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n439), .B1(new_n430), .B2(new_n431), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n429), .ZN(new_n441));
  INV_X1    g240(.A(new_n427), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n422), .A2(new_n427), .A3(new_n429), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n444), .A3(new_n437), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n440), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n401), .A2(new_n405), .B1(new_n438), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n202), .B1(new_n375), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n266), .B1(new_n258), .B2(new_n262), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n268), .A2(new_n265), .A3(new_n269), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n369), .B(new_n370), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n360), .ZN(new_n454));
  OR3_X1    g253(.A1(new_n371), .A2(new_n360), .A3(new_n367), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n452), .A2(new_n454), .A3(new_n455), .A4(new_n202), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n401), .A2(new_n405), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n447), .A2(new_n438), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT37), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n403), .B2(new_n387), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n386), .A2(new_n461), .A3(new_n387), .A4(new_n393), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n397), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT38), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n402), .A2(new_n389), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n241), .B1(new_n382), .B2(new_n383), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT37), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT38), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n468), .A2(new_n469), .A3(new_n397), .A4(new_n463), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n447), .A2(new_n438), .A3(new_n400), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n465), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT39), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT82), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n416), .A2(new_n421), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n474), .B1(new_n475), .B2(new_n423), .ZN(new_n476));
  AOI211_X1 g275(.A(KEYINPUT82), .B(new_n417), .C1(new_n416), .C2(new_n421), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n238), .A2(new_n351), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT77), .B1(new_n220), .B2(KEYINPUT3), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n481), .A2(new_n415), .B1(new_n420), .B2(new_n419), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT82), .B1(new_n482), .B2(new_n417), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n475), .A2(new_n474), .A3(new_n423), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n424), .A2(new_n425), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n473), .B1(new_n485), .B2(new_n417), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n478), .A2(new_n487), .A3(KEYINPUT40), .A4(new_n439), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT83), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n483), .A2(new_n484), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n437), .B1(new_n491), .B2(new_n473), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n492), .A2(KEYINPUT83), .A3(KEYINPUT40), .A4(new_n487), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n439), .A3(new_n487), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT40), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n495), .A2(new_n496), .B1(new_n432), .B2(new_n437), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n494), .A2(new_n405), .A3(new_n401), .A4(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n472), .A2(new_n498), .A3(new_n452), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n374), .A2(KEYINPUT36), .A3(new_n372), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n454), .A2(new_n455), .A3(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n500), .B(new_n502), .C1(new_n448), .C2(new_n452), .ZN(new_n503));
  OAI22_X1  g302(.A1(new_n449), .A2(new_n460), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G113gat), .B(G141gat), .ZN(new_n505));
  INV_X1    g304(.A(G197gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT11), .B(G169gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT12), .ZN(new_n510));
  NAND2_X1  g309(.A1(G229gat), .A2(G233gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT13), .ZN(new_n512));
  NOR2_X1   g311(.A1(G29gat), .A2(G36gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT14), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(G29gat), .A2(G36gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT84), .ZN(new_n517));
  XNOR2_X1  g316(.A(G43gat), .B(G50gat), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n515), .B(new_n517), .C1(KEYINPUT15), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(KEYINPUT15), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT85), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT85), .ZN(new_n523));
  INV_X1    g322(.A(new_n520), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n519), .A2(new_n524), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G15gat), .B(G22gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT16), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(G1gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT86), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n531), .B(new_n532), .C1(G1gat), .C2(new_n529), .ZN(new_n533));
  INV_X1    g332(.A(G8gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n535), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n522), .A2(new_n537), .A3(new_n527), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n512), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n535), .B(KEYINPUT87), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT17), .B1(new_n522), .B2(new_n527), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n521), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n540), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(new_n511), .A3(new_n538), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT18), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n539), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n544), .A2(KEYINPUT18), .A3(new_n511), .A4(new_n538), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n510), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(new_n548), .A3(new_n510), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n504), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(KEYINPUT88), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G57gat), .B(G64gat), .Z(new_n556));
  NAND2_X1  g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT90), .ZN(new_n560));
  NOR2_X1   g359(.A1(G71gat), .A2(G78gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n560), .B1(new_n561), .B2(KEYINPUT89), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT89), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n563), .B(KEYINPUT90), .C1(G71gat), .C2(G78gat), .ZN(new_n564));
  AOI22_X1  g363(.A1(new_n556), .A2(new_n559), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(new_n557), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n562), .A2(new_n564), .ZN(new_n567));
  INV_X1    g366(.A(G64gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(G57gat), .ZN(new_n569));
  INV_X1    g368(.A(G57gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(G64gat), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n559), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n567), .A2(new_n572), .A3(new_n557), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n559), .A3(new_n561), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n566), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT21), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n535), .ZN(new_n578));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G127gat), .B(G155gat), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n576), .A2(KEYINPUT21), .ZN(new_n585));
  XOR2_X1   g384(.A(G183gat), .B(G211gat), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT93), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n585), .B(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(KEYINPUT91), .B(KEYINPUT20), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n582), .A2(new_n583), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n582), .A2(new_n583), .ZN(new_n593));
  INV_X1    g392(.A(new_n590), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(G232gat), .A2(G233gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(KEYINPUT41), .ZN(new_n598));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT94), .B(KEYINPUT96), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G99gat), .A2(G106gat), .ZN(new_n604));
  INV_X1    g403(.A(G85gat), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(KEYINPUT8), .A2(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G85gat), .A2(G92gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT7), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G99gat), .B(G106gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT95), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n610), .A2(new_n611), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n613), .B1(new_n616), .B2(new_n607), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  AOI211_X1 g417(.A(KEYINPUT95), .B(new_n613), .C1(new_n616), .C2(new_n607), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n528), .A2(new_n542), .ZN(new_n622));
  INV_X1    g421(.A(new_n543), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n597), .A2(KEYINPUT41), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n528), .B2(new_n620), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n603), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n626), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n620), .B1(new_n541), .B2(new_n543), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n629), .A3(new_n602), .ZN(new_n630));
  XOR2_X1   g429(.A(G190gat), .B(G218gat), .Z(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n627), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n632), .B1(new_n627), .B2(new_n630), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n601), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n627), .A2(new_n630), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n631), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n627), .A2(new_n630), .A3(new_n632), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n637), .A2(new_n600), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n596), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G176gat), .B(G204gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OAI22_X1  g444(.A1(new_n618), .A2(new_n619), .B1(new_n566), .B2(new_n575), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n573), .A2(new_n574), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n565), .A2(new_n557), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT97), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n612), .A2(new_n649), .A3(new_n614), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n612), .A2(new_n614), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n616), .A2(new_n613), .A3(new_n607), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(KEYINPUT97), .A3(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n647), .A2(new_n648), .A3(new_n650), .A4(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT10), .B1(new_n646), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n576), .A2(KEYINPUT10), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(new_n620), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(G230gat), .A2(G233gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n659), .B(KEYINPUT98), .Z(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n659), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n646), .A2(new_n663), .A3(new_n654), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n645), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT99), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n658), .A2(new_n663), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n668), .A2(new_n645), .A3(new_n664), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n553), .B2(KEYINPUT88), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n555), .A2(new_n642), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n458), .B(KEYINPUT100), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G1gat), .ZN(G1324gat));
  INV_X1    g476(.A(new_n457), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT101), .B(KEYINPUT16), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(new_n534), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n674), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(KEYINPUT42), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT42), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n674), .A2(new_n678), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n684), .B2(G8gat), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n682), .B1(new_n685), .B2(new_n681), .ZN(G1325gat));
  NAND2_X1  g485(.A1(new_n500), .A2(new_n502), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n674), .A2(G15gat), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n454), .A2(new_n455), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(G15gat), .B1(new_n674), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n688), .A2(new_n691), .ZN(G1326gat));
  NOR2_X1   g491(.A1(new_n673), .A2(new_n452), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT43), .B(G22gat), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  NOR2_X1   g494(.A1(new_n596), .A2(new_n640), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n555), .A2(new_n672), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(G29gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n675), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT45), .Z(new_n701));
  INV_X1    g500(.A(new_n675), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n635), .A2(new_n639), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n504), .A2(KEYINPUT44), .A3(new_n703), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n591), .A2(new_n595), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n499), .B2(new_n503), .ZN(new_n708));
  INV_X1    g507(.A(new_n687), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n472), .A2(new_n498), .A3(new_n452), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n452), .B1(new_n457), .B2(new_n458), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n709), .A2(new_n710), .A3(new_n712), .A4(KEYINPUT102), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n449), .B2(new_n460), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n374), .A2(new_n372), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n452), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT35), .B1(new_n718), .B2(new_n459), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n689), .A2(new_n271), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(new_n202), .A3(new_n448), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n719), .A2(new_n721), .A3(KEYINPUT103), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n703), .B1(new_n714), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n706), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n547), .A2(new_n548), .A3(new_n510), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n549), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n671), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT104), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n503), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT102), .B1(new_n732), .B2(new_n710), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n499), .A2(new_n503), .A3(new_n707), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n716), .B(new_n722), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT44), .B1(new_n735), .B2(new_n703), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n737));
  INV_X1    g536(.A(new_n729), .ZN(new_n738));
  NOR4_X1   g537(.A1(new_n736), .A2(new_n737), .A3(new_n706), .A4(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n702), .B1(new_n731), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n701), .B1(new_n698), .B2(new_n741), .ZN(G1328gat));
  NOR2_X1   g541(.A1(new_n457), .A2(G36gat), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n555), .A2(new_n672), .A3(new_n696), .A4(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n745));
  OR3_X1    g544(.A1(new_n744), .A2(new_n745), .A3(KEYINPUT46), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n744), .B2(KEYINPUT46), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(KEYINPUT46), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n457), .B1(new_n731), .B2(new_n740), .ZN(new_n750));
  INV_X1    g549(.A(G36gat), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n746), .B(new_n749), .C1(new_n750), .C2(new_n751), .ZN(G1329gat));
  NOR3_X1   g551(.A1(new_n697), .A2(G43gat), .A3(new_n689), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n726), .A2(new_n729), .ZN(new_n755));
  OAI21_X1  g554(.A(G43gat), .B1(new_n755), .B2(new_n709), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(new_n756), .A3(KEYINPUT47), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n687), .B1(new_n730), .B2(new_n739), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n753), .B1(new_n758), .B2(G43gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n759), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g559(.A(KEYINPUT48), .B(G50gat), .C1(new_n755), .C2(new_n452), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n452), .A2(G50gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT106), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n697), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n761), .B(new_n764), .C1(new_n765), .C2(KEYINPUT48), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n697), .A2(new_n765), .A3(new_n763), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n271), .B1(new_n730), .B2(new_n739), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n768), .B2(G50gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n766), .B1(new_n769), .B2(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g569(.A1(new_n642), .A2(new_n735), .A3(new_n728), .A4(new_n671), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n675), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g572(.A(new_n457), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT108), .Z(new_n775));
  NAND2_X1  g574(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT109), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n771), .A2(new_n778), .A3(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n780), .B(new_n781), .ZN(G1333gat));
  NAND2_X1  g581(.A1(new_n771), .A2(new_n687), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n689), .A2(G71gat), .ZN(new_n784));
  AOI22_X1  g583(.A1(new_n783), .A2(G71gat), .B1(new_n771), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n271), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G78gat), .ZN(G1335gat));
  INV_X1    g587(.A(new_n671), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n552), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n726), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G85gat), .B1(new_n791), .B2(new_n702), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n596), .A2(new_n552), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n724), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n796));
  OR2_X1    g595(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(KEYINPUT110), .B(KEYINPUT51), .C1(new_n724), .C2(new_n794), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(new_n671), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n675), .A2(new_n605), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n792), .B1(new_n800), .B2(new_n801), .ZN(G1336gat));
  OAI21_X1  g601(.A(G92gat), .B1(new_n791), .B2(new_n457), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n457), .A2(G92gat), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT52), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n803), .B(new_n808), .C1(new_n800), .C2(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(G1337gat));
  OAI21_X1  g609(.A(G99gat), .B1(new_n791), .B2(new_n709), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n689), .A2(G99gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n800), .B2(new_n812), .ZN(G1338gat));
  OAI21_X1  g612(.A(G106gat), .B1(new_n791), .B2(new_n452), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n452), .A2(G106gat), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n798), .A2(new_n799), .A3(new_n671), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT53), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT111), .B1(new_n791), .B2(new_n452), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n726), .A2(new_n820), .A3(new_n271), .A4(new_n790), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n819), .A2(G106gat), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n816), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n818), .B1(new_n822), .B2(new_n824), .ZN(G1339gat));
  INV_X1    g624(.A(new_n655), .ZN(new_n826));
  INV_X1    g625(.A(new_n657), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n827), .A3(new_n661), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n828), .B(KEYINPUT54), .C1(new_n658), .C2(new_n663), .ZN(new_n829));
  XNOR2_X1  g628(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n660), .B(new_n830), .C1(new_n655), .C2(new_n657), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n831), .A2(KEYINPUT113), .A3(new_n645), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT113), .B1(new_n831), .B2(new_n645), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n829), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n829), .B(KEYINPUT55), .C1(new_n832), .C2(new_n833), .ZN(new_n837));
  AND4_X1   g636(.A1(KEYINPUT114), .A2(new_n836), .A3(new_n670), .A4(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n669), .B1(new_n834), .B2(new_n835), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT114), .B1(new_n839), .B2(new_n837), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n552), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n511), .B1(new_n544), .B2(new_n538), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n536), .A2(new_n538), .A3(new_n512), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n509), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n551), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n671), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n703), .B1(new_n841), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n639), .A3(new_n635), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n836), .A2(new_n670), .A3(new_n837), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n839), .A2(KEYINPUT114), .A3(new_n837), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n849), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n705), .B1(new_n848), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n642), .A2(new_n728), .A3(new_n789), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n702), .A2(new_n678), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n720), .ZN(new_n860));
  OAI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n728), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n375), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n334), .A2(new_n335), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n552), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n861), .B1(new_n862), .B2(new_n864), .ZN(G1340gat));
  OAI21_X1  g664(.A(G120gat), .B1(new_n860), .B2(new_n789), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n671), .A2(new_n333), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n862), .B2(new_n867), .ZN(G1341gat));
  OAI21_X1  g667(.A(G127gat), .B1(new_n860), .B2(new_n705), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n596), .A2(new_n329), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n862), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n871), .B(new_n872), .ZN(G1342gat));
  NAND4_X1  g672(.A1(new_n859), .A2(new_n327), .A3(new_n703), .A4(new_n375), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n860), .B2(new_n640), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G1343gat));
  NOR2_X1   g677(.A1(new_n687), .A2(new_n452), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n857), .A2(new_n858), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n552), .A2(new_n211), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(KEYINPUT58), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n271), .A2(KEYINPUT57), .ZN(new_n884));
  INV_X1    g683(.A(new_n850), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n552), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n703), .B1(new_n886), .B2(new_n847), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n705), .B1(new_n854), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n884), .B1(new_n888), .B2(new_n856), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n728), .B1(new_n852), .B2(new_n853), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n789), .A2(new_n845), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n640), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n640), .A2(new_n845), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n893), .B1(new_n840), .B2(new_n838), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n596), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n641), .A2(new_n552), .A3(new_n671), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n271), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n889), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n858), .A2(new_n709), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n899), .A2(new_n728), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G141gat), .B1(new_n901), .B2(KEYINPUT117), .ZN(new_n902));
  INV_X1    g701(.A(new_n900), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT57), .B1(new_n857), .B2(new_n271), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n552), .B(new_n903), .C1(new_n904), .C2(new_n889), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT117), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n883), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n882), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n909), .B1(new_n901), .B2(new_n211), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT116), .B1(new_n910), .B2(KEYINPUT58), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n882), .B1(new_n905), .B2(G141gat), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT116), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT58), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n908), .B1(new_n911), .B2(new_n915), .ZN(G1344gat));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n897), .A2(KEYINPUT57), .ZN(new_n918));
  INV_X1    g717(.A(new_n887), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n893), .A2(new_n885), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n596), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n898), .B(new_n271), .C1(new_n921), .C2(new_n896), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n900), .B(KEYINPUT118), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n918), .A2(new_n671), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G148gat), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n671), .B(new_n903), .C1(new_n904), .C2(new_n889), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n203), .A2(KEYINPUT59), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n925), .A2(KEYINPUT59), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n880), .A2(G148gat), .A3(new_n789), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n917), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n929), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n926), .A2(new_n927), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT59), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n933), .B1(new_n924), .B2(G148gat), .ZN(new_n934));
  OAI211_X1 g733(.A(KEYINPUT119), .B(new_n931), .C1(new_n932), .C2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n930), .A2(new_n935), .ZN(G1345gat));
  INV_X1    g735(.A(new_n880), .ZN(new_n937));
  AOI21_X1  g736(.A(G155gat), .B1(new_n937), .B2(new_n596), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n899), .A2(new_n900), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n596), .A2(G155gat), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT120), .Z(new_n941));
  AOI21_X1  g740(.A(new_n938), .B1(new_n939), .B2(new_n941), .ZN(G1346gat));
  INV_X1    g741(.A(G162gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n937), .A2(new_n943), .A3(new_n703), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n899), .A2(new_n640), .A3(new_n900), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(new_n943), .ZN(G1347gat));
  AOI21_X1  g745(.A(new_n675), .B1(new_n855), .B2(new_n856), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n718), .A2(new_n457), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT121), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n290), .A3(new_n552), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n689), .A2(new_n457), .A3(new_n271), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n947), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(G169gat), .B1(new_n953), .B2(new_n728), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n951), .A2(new_n954), .ZN(G1348gat));
  AOI21_X1  g754(.A(G176gat), .B1(new_n950), .B2(new_n671), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n947), .A2(G176gat), .A3(new_n671), .A4(new_n952), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(KEYINPUT122), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(KEYINPUT122), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(G1349gat));
  NAND3_X1  g759(.A1(new_n950), .A2(new_n596), .A3(new_n313), .ZN(new_n961));
  OAI21_X1  g760(.A(G183gat), .B1(new_n953), .B2(new_n705), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n964), .A2(KEYINPUT60), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(KEYINPUT60), .ZN(new_n966));
  XOR2_X1   g765(.A(new_n966), .B(KEYINPUT124), .Z(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  OR3_X1    g767(.A1(new_n963), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n963), .B2(new_n965), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1350gat));
  OAI21_X1  g770(.A(G190gat), .B1(new_n953), .B2(new_n640), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT61), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n950), .A2(new_n302), .A3(new_n703), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(G1351gat));
  NOR3_X1   g774(.A1(new_n687), .A2(new_n457), .A3(new_n675), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n918), .A2(new_n922), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(G197gat), .B1(new_n977), .B2(new_n728), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n687), .A2(new_n452), .A3(new_n457), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n947), .A2(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n981), .A2(new_n506), .A3(new_n552), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n978), .A2(new_n982), .ZN(G1352gat));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n789), .A2(G204gat), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n981), .A2(KEYINPUT125), .A3(new_n985), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT125), .ZN(new_n987));
  INV_X1    g786(.A(new_n985), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n987), .B1(new_n980), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n984), .B1(new_n990), .B2(KEYINPUT62), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT62), .ZN(new_n993));
  NAND4_X1  g792(.A1(new_n986), .A2(KEYINPUT126), .A3(new_n993), .A4(new_n989), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n918), .A2(new_n671), .A3(new_n922), .ZN(new_n995));
  INV_X1    g794(.A(new_n976), .ZN(new_n996));
  OAI21_X1  g795(.A(G204gat), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND4_X1  g796(.A1(new_n991), .A2(new_n992), .A3(new_n994), .A4(new_n997), .ZN(G1353gat));
  NAND4_X1  g797(.A1(new_n918), .A2(new_n596), .A3(new_n922), .A4(new_n976), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(G211gat), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT63), .ZN(new_n1001));
  OAI21_X1  g800(.A(KEYINPUT127), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n1004));
  NAND4_X1  g803(.A1(new_n999), .A2(new_n1004), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n981), .A2(new_n223), .A3(new_n596), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1006), .A2(new_n1007), .ZN(G1354gat));
  NOR3_X1   g807(.A1(new_n977), .A2(new_n224), .A3(new_n640), .ZN(new_n1009));
  AOI21_X1  g808(.A(G218gat), .B1(new_n981), .B2(new_n703), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n1009), .A2(new_n1010), .ZN(G1355gat));
endmodule


