//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1224, new_n1225,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NAND2_X1  g0005(.A1(G107), .A2(G264), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  INV_X1    g0007(.A(G226), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G58), .ZN(new_n210));
  INV_X1    g0010(.A(G232), .ZN(new_n211));
  INV_X1    g0011(.A(G77), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n209), .B(new_n214), .C1(G116), .C2(G270), .ZN(new_n215));
  AND2_X1   g0015(.A1(KEYINPUT66), .A2(G68), .ZN(new_n216));
  NOR2_X1   g0016(.A1(KEYINPUT66), .A2(G68), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(KEYINPUT67), .B(G238), .Z(new_n219));
  OAI21_X1  g0019(.A(new_n215), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT68), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n205), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT64), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n207), .B1(new_n202), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n226), .B1(new_n225), .B2(new_n202), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT65), .Z(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n205), .A2(G13), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT0), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n224), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G97), .B(G107), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  XNOR2_X1  g0052(.A(KEYINPUT73), .B(G200), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G222), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n261), .A2(new_n262), .B1(new_n212), .B2(new_n259), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n260), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT70), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n263), .B1(new_n268), .B2(G223), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G1), .A3(G13), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(new_n271), .A3(G274), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n271), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(new_n275), .ZN(new_n279));
  XOR2_X1   g0079(.A(KEYINPUT69), .B(G226), .Z(new_n280));
  AOI21_X1  g0080(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n254), .B1(new_n272), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT71), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(new_n205), .B2(new_n256), .ZN(new_n285));
  NAND4_X1  g0085(.A1(KEYINPUT71), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G1), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G13), .A3(G20), .ZN(new_n288));
  AND4_X1   g0088(.A1(new_n229), .A2(new_n285), .A3(new_n286), .A4(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n230), .A2(G1), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(G50), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n285), .A2(new_n229), .A3(new_n286), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT8), .B(G58), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n230), .A2(G33), .ZN(new_n295));
  INV_X1    g0095(.A(G150), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n294), .A2(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n230), .B1(new_n201), .B2(new_n207), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n293), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n292), .B(new_n301), .C1(G50), .C2(new_n288), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT9), .ZN(new_n303));
  OAI211_X1 g0103(.A(G190), .B(new_n281), .C1(new_n269), .C2(new_n271), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n283), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n283), .A2(new_n303), .A3(new_n307), .A4(new_n304), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G179), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n277), .B1(G244), .B2(new_n279), .ZN(new_n311));
  INV_X1    g0111(.A(G107), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n261), .A2(new_n211), .B1(new_n312), .B2(new_n259), .ZN(new_n313));
  INV_X1    g0113(.A(new_n219), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n268), .B2(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n310), .B(new_n311), .C1(new_n315), .C2(new_n271), .ZN(new_n316));
  INV_X1    g0116(.A(new_n294), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n317), .A2(new_n297), .B1(G20), .B2(G77), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT72), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT15), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(G87), .ZN(new_n321));
  INV_X1    g0121(.A(G87), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(KEYINPUT15), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n319), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(KEYINPUT15), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n320), .A2(G87), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT72), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n318), .B1(new_n328), .B2(new_n295), .ZN(new_n329));
  INV_X1    g0129(.A(new_n288), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n329), .A2(new_n293), .B1(new_n212), .B2(new_n330), .ZN(new_n331));
  NOR4_X1   g0131(.A1(new_n293), .A2(new_n212), .A3(new_n330), .A4(new_n290), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n315), .A2(new_n271), .ZN(new_n335));
  INV_X1    g0135(.A(new_n311), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n316), .B(new_n334), .C1(new_n337), .C2(G169), .ZN(new_n338));
  INV_X1    g0138(.A(new_n334), .ZN(new_n339));
  OAI211_X1 g0139(.A(G190), .B(new_n311), .C1(new_n315), .C2(new_n271), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n339), .B(new_n340), .C1(new_n337), .C2(new_n253), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n272), .A2(new_n282), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n310), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n344), .B(new_n302), .C1(G169), .C2(new_n343), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n309), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n218), .A2(G20), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n347), .B1(new_n207), .B2(new_n298), .C1(new_n212), .C2(new_n295), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n293), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT11), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G13), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(G1), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n218), .A2(KEYINPUT12), .A3(G20), .A4(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT12), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n288), .B2(G68), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n351), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n289), .A2(G68), .A3(new_n291), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n349), .B2(new_n350), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  XOR2_X1   g0160(.A(new_n276), .B(KEYINPUT74), .Z(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G97), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n211), .A2(G1698), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(G226), .B2(G1698), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n362), .B1(new_n364), .B2(new_n266), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n365), .A2(new_n278), .B1(new_n279), .B2(G238), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT13), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT13), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n361), .A2(new_n369), .A3(new_n366), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G190), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n360), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n371), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT75), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT75), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n371), .A2(new_n377), .A3(G200), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n373), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G169), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n368), .B2(new_n370), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT14), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n381), .A2(new_n382), .B1(new_n371), .B2(new_n310), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n381), .A2(KEYINPUT76), .A3(new_n382), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT76), .B1(new_n381), .B2(new_n382), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n384), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n360), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n379), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n294), .A2(new_n290), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n289), .A2(new_n391), .B1(new_n330), .B2(new_n294), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT77), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT7), .B1(new_n266), .B2(new_n230), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n230), .A4(new_n258), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n395), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n257), .A2(new_n230), .A3(new_n258), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n395), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n218), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g0204(.A(KEYINPUT66), .B(G68), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n201), .B1(new_n405), .B2(G58), .ZN(new_n406));
  INV_X1    g0206(.A(G159), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n406), .A2(new_n230), .B1(new_n407), .B2(new_n298), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n394), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n293), .ZN(new_n410));
  INV_X1    g0210(.A(G68), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n400), .A2(new_n401), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(new_n397), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n410), .B1(new_n414), .B2(KEYINPUT16), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n393), .B1(new_n409), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n287), .B1(G41), .B2(G45), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n271), .A2(G232), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT78), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n276), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n419), .B1(new_n276), .B2(new_n418), .ZN(new_n421));
  OR2_X1    g0221(.A1(G223), .A2(G1698), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n208), .A2(G1698), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n422), .B(new_n423), .C1(new_n264), .C2(new_n265), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G33), .A2(G87), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n271), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n420), .A2(new_n421), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G179), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n276), .A2(new_n418), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT78), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n424), .A2(new_n425), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n278), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n276), .A2(new_n418), .A3(new_n419), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G169), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT18), .B1(new_n416), .B2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n430), .A2(new_n432), .A3(new_n372), .A4(new_n433), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n427), .B2(G200), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n416), .A2(KEYINPUT17), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT77), .B1(new_n412), .B2(new_n397), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n405), .B1(new_n442), .B2(new_n402), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n202), .B1(new_n218), .B2(new_n210), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n444), .A2(G20), .B1(G159), .B2(new_n297), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT16), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(G68), .B1(new_n396), .B2(new_n398), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n447), .A3(KEYINPUT16), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n293), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n440), .B(new_n392), .C1(new_n446), .C2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n392), .B1(new_n446), .B2(new_n449), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT18), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(new_n436), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n438), .A2(new_n441), .A3(new_n452), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n346), .A2(new_n390), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT79), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n346), .A2(new_n390), .A3(KEYINPUT79), .A4(new_n457), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n327), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT72), .B1(new_n325), .B2(new_n326), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT84), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n287), .A2(G33), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n465), .A2(new_n289), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n286), .A2(new_n229), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n469), .A2(new_n285), .A3(new_n288), .A4(new_n467), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT84), .B1(new_n470), .B2(new_n328), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n230), .B(G68), .C1(new_n264), .C2(new_n265), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n230), .A2(G33), .A3(G97), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT19), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT82), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT82), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT19), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n230), .B1(new_n481), .B2(new_n362), .ZN(new_n482));
  OR2_X1    g0282(.A1(KEYINPUT83), .A2(G87), .ZN(new_n483));
  NOR2_X1   g0283(.A1(G97), .A2(G107), .ZN(new_n484));
  NAND2_X1  g0284(.A1(KEYINPUT83), .A2(G87), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n480), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n487), .A2(new_n410), .B1(new_n288), .B2(new_n465), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT85), .B1(new_n472), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n482), .A2(new_n486), .ZN(new_n490));
  INV_X1    g0290(.A(new_n480), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n492), .A2(new_n293), .B1(new_n330), .B2(new_n328), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT85), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n468), .A2(new_n471), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n259), .A2(G244), .A3(G1698), .ZN(new_n497));
  OAI211_X1 g0297(.A(G238), .B(new_n260), .C1(new_n264), .C2(new_n265), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G116), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n278), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n271), .B(G250), .C1(G1), .C2(new_n274), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n274), .A2(G1), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n271), .A2(G274), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n501), .A2(G179), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n505), .B1(new_n500), .B2(new_n278), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n380), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n489), .A2(new_n496), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n470), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n488), .B1(G87), .B2(new_n511), .ZN(new_n512));
  AOI211_X1 g0312(.A(new_n372), .B(new_n505), .C1(new_n278), .C2(new_n500), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n253), .B1(new_n501), .B2(new_n506), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n510), .A2(KEYINPUT86), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT86), .B1(new_n510), .B2(new_n516), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n259), .A2(G250), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n260), .B1(new_n520), .B2(KEYINPUT4), .ZN(new_n521));
  AND2_X1   g0321(.A1(KEYINPUT4), .A2(G244), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n260), .B(new_n522), .C1(new_n264), .C2(new_n265), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G283), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n213), .B1(new_n257), .B2(new_n258), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n523), .B(new_n524), .C1(new_n525), .C2(KEYINPUT4), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n278), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g0327(.A(KEYINPUT5), .B(G41), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n528), .A2(G274), .A3(new_n271), .A4(new_n503), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n278), .B1(new_n503), .B2(new_n528), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n530), .B1(G257), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT80), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT80), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n527), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(G190), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT81), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT81), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n534), .A2(new_n539), .A3(G190), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n533), .A2(G200), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n312), .B1(new_n399), .B2(new_n403), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT6), .ZN(new_n543));
  INV_X1    g0343(.A(G97), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n543), .A2(new_n544), .A3(G107), .ZN(new_n545));
  XNOR2_X1  g0345(.A(G97), .B(G107), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(new_n543), .ZN(new_n547));
  OAI22_X1  g0347(.A1(new_n547), .A2(new_n230), .B1(new_n212), .B2(new_n298), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n293), .B1(new_n542), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n288), .A2(G97), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n511), .B2(G97), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n541), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n538), .A2(new_n540), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n534), .A2(new_n536), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n380), .ZN(new_n555));
  INV_X1    g0355(.A(new_n533), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n549), .A2(new_n551), .B1(new_n556), .B2(new_n310), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n259), .A2(G264), .A3(G1698), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n259), .A2(G257), .A3(new_n260), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n266), .A2(G303), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n278), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n271), .A2(G274), .A3(new_n503), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n531), .A2(G270), .B1(new_n565), .B2(new_n528), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(new_n375), .ZN(new_n569));
  AOI21_X1  g0369(.A(G20), .B1(G33), .B2(G283), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n256), .A2(G97), .ZN(new_n571));
  INV_X1    g0371(.A(G116), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n570), .A2(new_n571), .B1(G20), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n293), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT20), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n293), .A2(KEYINPUT20), .A3(new_n573), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n289), .A2(KEYINPUT87), .A3(G116), .A4(new_n467), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT87), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n470), .B2(new_n572), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n353), .A2(G20), .A3(new_n572), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n578), .A2(new_n579), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n567), .A2(new_n372), .ZN(new_n584));
  OR3_X1    g0384(.A1(new_n569), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n259), .A2(G257), .A3(G1698), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n259), .A2(G250), .A3(new_n260), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G294), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n278), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n531), .A2(G264), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(new_n529), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G200), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n230), .B(G87), .C1(new_n264), .C2(new_n265), .ZN(new_n594));
  NAND2_X1  g0394(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n259), .A2(new_n230), .A3(G87), .A4(new_n595), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT24), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n499), .A2(G20), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT23), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n230), .B2(G107), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n312), .A2(KEYINPUT23), .A3(G20), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n599), .A2(new_n600), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n600), .B1(new_n599), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n293), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n330), .A2(new_n312), .ZN(new_n609));
  XNOR2_X1  g0409(.A(new_n609), .B(KEYINPUT25), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n511), .B2(G107), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n590), .A2(G190), .A3(new_n529), .A4(new_n591), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n593), .A2(new_n608), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n585), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n583), .A2(G169), .A3(new_n567), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT21), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI211_X1 g0417(.A(new_n616), .B(new_n380), .C1(new_n564), .C2(new_n566), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n567), .A2(new_n310), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n583), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n608), .A2(new_n611), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n592), .A2(new_n380), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(G179), .B2(new_n592), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n617), .B(new_n620), .C1(new_n621), .C2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n614), .A2(new_n624), .ZN(new_n625));
  AND4_X1   g0425(.A1(new_n462), .A2(new_n519), .A3(new_n559), .A4(new_n625), .ZN(G372));
  INV_X1    g0426(.A(new_n345), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n338), .A2(KEYINPUT89), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n338), .A2(KEYINPUT89), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n376), .A2(new_n378), .ZN(new_n631));
  INV_X1    g0431(.A(new_n373), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n630), .A2(new_n633), .B1(new_n389), .B2(new_n388), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n441), .A2(new_n452), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n438), .B(new_n455), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n627), .B1(new_n636), .B2(new_n309), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n555), .A2(new_n557), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n519), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n493), .A2(new_n495), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n512), .A2(new_n515), .B1(new_n509), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n642), .A2(new_n555), .A3(new_n643), .A4(new_n557), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n509), .A2(new_n641), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n516), .A2(new_n613), .A3(new_n645), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n553), .A2(new_n647), .A3(new_n624), .A4(new_n558), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n640), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n462), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n637), .A2(new_n651), .ZN(G369));
  NAND2_X1  g0452(.A1(new_n617), .A2(new_n620), .ZN(new_n653));
  INV_X1    g0453(.A(new_n353), .ZN(new_n654));
  OR3_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .A3(G20), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT27), .B1(new_n654), .B2(G20), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n583), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g0460(.A(new_n653), .B(new_n660), .Z(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n585), .ZN(new_n662));
  INV_X1    g0462(.A(G330), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n621), .A2(new_n623), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(new_n659), .ZN(new_n666));
  INV_X1    g0466(.A(new_n659), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n613), .B1(new_n621), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n666), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n659), .B1(new_n617), .B2(new_n620), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT90), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n666), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(G399));
  INV_X1    g0474(.A(new_n233), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n486), .A2(G116), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G1), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n227), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n647), .A2(new_n624), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT92), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n559), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n638), .A2(new_n642), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n686), .A2(KEYINPUT26), .B1(new_n641), .B2(new_n509), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n648), .A2(KEYINPUT92), .ZN(new_n688));
  INV_X1    g0488(.A(new_n518), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n510), .A2(KEYINPUT86), .A3(new_n516), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n689), .A2(new_n643), .A3(new_n690), .A4(new_n638), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n685), .A2(new_n687), .A3(new_n688), .A4(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n682), .B1(new_n692), .B2(new_n667), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n650), .A2(new_n667), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(KEYINPUT29), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n590), .A2(new_n591), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n501), .A2(new_n506), .ZN(new_n697));
  NOR4_X1   g0497(.A1(new_n567), .A2(new_n696), .A3(new_n697), .A4(new_n310), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(new_n534), .A3(new_n536), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT30), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n568), .A2(G179), .A3(new_n508), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(new_n533), .A3(new_n592), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT91), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n667), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n519), .A2(new_n625), .A3(new_n559), .A4(new_n667), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n704), .B1(KEYINPUT31), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n700), .A2(new_n702), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n708), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  AOI211_X1 g0511(.A(new_n693), .B(new_n695), .C1(G330), .C2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n681), .B1(new_n712), .B2(G1), .ZN(G364));
  XNOR2_X1  g0513(.A(new_n664), .B(KEYINPUT93), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n352), .A2(G20), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n287), .B1(new_n715), .B2(G45), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n676), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n662), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n719), .B1(new_n720), .B2(G330), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n714), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g0522(.A(new_n722), .B(KEYINPUT94), .Z(new_n723));
  AOI21_X1  g0523(.A(new_n229), .B1(G20), .B2(new_n380), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n230), .A2(new_n310), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G200), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G190), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  XOR2_X1   g0529(.A(KEYINPUT33), .B(G317), .Z(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n726), .A2(G190), .A3(new_n375), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n230), .A2(G179), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G190), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n733), .A2(G322), .B1(new_n737), .B2(G329), .ZN(new_n738));
  INV_X1    g0538(.A(G311), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n726), .A2(new_n735), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n738), .B(new_n266), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n734), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n253), .A2(new_n742), .A3(G190), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n731), .B(new_n741), .C1(G283), .C2(new_n743), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n372), .A2(G179), .A3(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n230), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n727), .A2(new_n372), .ZN(new_n748));
  AOI22_X1  g0548(.A1(G294), .A2(new_n747), .B1(new_n748), .B2(G326), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n749), .B(KEYINPUT96), .Z(new_n750));
  INV_X1    g0550(.A(G303), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n253), .A2(new_n742), .A3(new_n372), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT95), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(KEYINPUT95), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n744), .B(new_n750), .C1(new_n751), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n746), .A2(new_n544), .ZN(new_n757));
  INV_X1    g0557(.A(new_n748), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n207), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n757), .B(new_n759), .C1(G68), .C2(new_n728), .ZN(new_n760));
  INV_X1    g0560(.A(new_n755), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n483), .A2(new_n485), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n743), .A2(G107), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n259), .B1(new_n740), .B2(new_n212), .C1(new_n210), .C2(new_n732), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT32), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(new_n736), .B2(new_n407), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n737), .A2(KEYINPUT32), .A3(G159), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n760), .A2(new_n763), .A3(new_n764), .A4(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n725), .B1(new_n756), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G13), .A2(G33), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n724), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n228), .A2(new_n274), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n675), .A2(new_n259), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n776), .B(new_n777), .C1(new_n274), .C2(new_n248), .ZN(new_n778));
  INV_X1    g0578(.A(G355), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n259), .A2(new_n233), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n778), .B1(G116), .B2(new_n233), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n719), .B(new_n771), .C1(new_n775), .C2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n774), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n720), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n723), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT97), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(G396));
  NAND2_X1  g0587(.A1(new_n711), .A2(G330), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n339), .A2(new_n667), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n628), .A2(new_n629), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n342), .B1(new_n339), .B2(new_n667), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n694), .A2(new_n793), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n342), .A2(new_n667), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n643), .B1(new_n519), .B2(new_n638), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n646), .A2(new_n648), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n719), .B1(new_n788), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n801), .A2(KEYINPUT98), .B1(new_n788), .B2(new_n799), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(KEYINPUT98), .B2(new_n801), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n724), .A2(new_n772), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n718), .B1(G77), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n729), .A2(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n757), .B(new_n808), .C1(G303), .C2(new_n748), .ZN(new_n809));
  INV_X1    g0609(.A(new_n743), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n322), .ZN(new_n811));
  INV_X1    g0611(.A(G294), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n266), .B1(new_n732), .B2(new_n812), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n740), .A2(new_n572), .B1(new_n736), .B2(new_n739), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n809), .B(new_n815), .C1(new_n312), .C2(new_n755), .ZN(new_n816));
  INV_X1    g0616(.A(new_n740), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n733), .A2(G143), .B1(new_n817), .B2(G159), .ZN(new_n818));
  INV_X1    g0618(.A(G137), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n818), .B1(new_n729), .B2(new_n296), .C1(new_n819), .C2(new_n758), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT34), .Z(new_n821));
  NOR2_X1   g0621(.A1(new_n746), .A2(new_n210), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n266), .B(new_n822), .C1(G132), .C2(new_n737), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n823), .B1(new_n411), .B2(new_n810), .C1(new_n755), .C2(new_n207), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n816), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n806), .B1(new_n825), .B2(new_n724), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n792), .B2(new_n773), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n803), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G384));
  INV_X1    g0629(.A(new_n547), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n830), .A2(KEYINPUT35), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(KEYINPUT35), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n831), .A2(G116), .A3(new_n231), .A4(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(KEYINPUT99), .B(KEYINPUT36), .Z(new_n834));
  XNOR2_X1  g0634(.A(new_n833), .B(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n227), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n836), .B(G77), .C1(new_n210), .C2(new_n218), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n207), .A2(G68), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n287), .B(G13), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n450), .B(new_n841), .C1(new_n416), .C2(new_n657), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT100), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n453), .A2(new_n844), .A3(new_n436), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT100), .B1(new_n416), .B2(new_n437), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n843), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n414), .A2(KEYINPUT16), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n392), .B1(new_n848), .B2(new_n449), .ZN(new_n849));
  INV_X1    g0649(.A(new_n657), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n849), .B1(new_n436), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n450), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n847), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n456), .A2(new_n850), .A3(new_n849), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(KEYINPUT38), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n841), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n450), .B1(new_n416), .B2(new_n657), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n416), .A2(new_n437), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n846), .A2(new_n845), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n860), .B1(new_n842), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT102), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n456), .A2(new_n453), .A3(new_n850), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n860), .B(KEYINPUT102), .C1(new_n842), .C2(new_n861), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT103), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n868), .B1(new_n867), .B2(new_n869), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n856), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n704), .A2(KEYINPUT31), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n706), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n389), .A2(new_n659), .ZN(new_n876));
  INV_X1    g0676(.A(new_n387), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n383), .B1(new_n877), .B2(new_n385), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n633), .B(new_n876), .C1(new_n878), .C2(new_n360), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n389), .B(new_n659), .C1(new_n388), .C2(new_n379), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n881), .A2(new_n792), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n873), .A2(KEYINPUT40), .A3(new_n875), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n854), .A2(new_n855), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n869), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n856), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n875), .A2(new_n886), .A3(new_n882), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n462), .A2(new_n875), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n663), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n891), .B2(new_n890), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n850), .B1(new_n438), .B2(new_n455), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n338), .A2(new_n659), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n798), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n881), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n894), .B1(new_n900), .B2(new_n886), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n856), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n866), .A2(new_n865), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT102), .B1(new_n847), .B2(new_n860), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n869), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT103), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n903), .B1(new_n907), .B2(new_n870), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n902), .B1(new_n885), .B2(new_n856), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n878), .A2(new_n360), .A3(new_n659), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n901), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n462), .B1(new_n695), .B2(new_n693), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n637), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n913), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n893), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n287), .B2(new_n715), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n893), .A2(new_n916), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n840), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT104), .ZN(G367));
  NOR2_X1   g0721(.A1(new_n512), .A2(new_n667), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n642), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n645), .B2(new_n923), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT105), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n549), .A2(new_n551), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n559), .B1(new_n928), .B2(new_n667), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n638), .A2(new_n659), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(new_n669), .A3(new_n672), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT42), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n558), .B1(new_n929), .B2(new_n665), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n667), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n932), .A2(KEYINPUT42), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n927), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n938), .B(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n670), .B1(new_n929), .B2(new_n930), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n940), .B(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n676), .B(new_n943), .Z(new_n944));
  XOR2_X1   g0744(.A(new_n669), .B(new_n672), .Z(new_n945));
  NOR2_X1   g0745(.A1(new_n714), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n664), .B2(new_n945), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n712), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n673), .A2(new_n931), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT45), .Z(new_n951));
  NOR2_X1   g0751(.A1(new_n673), .A2(new_n931), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT44), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n951), .A2(new_n670), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n953), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(new_n664), .A3(new_n669), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n949), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n944), .B1(new_n957), .B2(new_n712), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n942), .B1(new_n958), .B2(new_n717), .ZN(new_n959));
  INV_X1    g0759(.A(new_n777), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n775), .B1(new_n233), .B2(new_n328), .C1(new_n244), .C2(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n961), .A2(new_n718), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n817), .A2(G283), .B1(new_n737), .B2(G317), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n963), .B(new_n266), .C1(new_n751), .C2(new_n732), .ZN(new_n964));
  AOI22_X1  g0764(.A1(G294), .A2(new_n728), .B1(new_n748), .B2(G311), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n312), .B2(new_n746), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n964), .B(new_n966), .C1(G97), .C2(new_n743), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n761), .A2(KEYINPUT46), .A3(G116), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT46), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n755), .B2(new_n572), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n746), .A2(new_n411), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n729), .A2(new_n407), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(G143), .C2(new_n748), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n733), .A2(G150), .B1(new_n737), .B2(G137), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n743), .A2(G77), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n266), .B1(new_n817), .B2(G50), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n974), .B(new_n978), .C1(new_n210), .C2(new_n755), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n971), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT47), .Z(new_n981));
  OAI221_X1 g0781(.A(new_n962), .B1(new_n925), .B2(new_n783), .C1(new_n981), .C2(new_n725), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n959), .A2(new_n982), .ZN(G387));
  OR2_X1    g0783(.A1(new_n669), .A2(new_n783), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n777), .B1(new_n241), .B2(new_n274), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n678), .B2(new_n780), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n294), .A2(G50), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT107), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n988), .A2(KEYINPUT50), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(KEYINPUT50), .ZN(new_n990));
  AOI21_X1  g0790(.A(G45), .B1(G68), .B2(G77), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n989), .A2(new_n678), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n986), .A2(new_n992), .B1(new_n312), .B2(new_n675), .ZN(new_n993));
  INV_X1    g0793(.A(new_n775), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n718), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n465), .A2(new_n747), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n207), .B2(new_n732), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT108), .Z(new_n998));
  NAND2_X1  g0798(.A1(new_n761), .A2(G77), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n259), .B1(new_n736), .B2(new_n296), .C1(new_n411), .C2(new_n740), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n407), .A2(new_n758), .B1(new_n729), .B2(new_n294), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(G97), .C2(new_n743), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n998), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n259), .B1(new_n737), .B2(G326), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n733), .A2(G317), .B1(new_n817), .B2(G303), .ZN(new_n1005));
  INV_X1    g0805(.A(G322), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1005), .B1(new_n729), .B2(new_n739), .C1(new_n1006), .C2(new_n758), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT48), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n807), .B2(new_n746), .C1(new_n812), .C2(new_n755), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT49), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1004), .B1(new_n572), .B2(new_n810), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1003), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n995), .B1(new_n1013), .B2(new_n724), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n947), .A2(new_n717), .B1(new_n984), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n676), .B(KEYINPUT109), .Z(new_n1016));
  NAND2_X1  g0816(.A1(new_n948), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n947), .A2(new_n712), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT110), .ZN(G393));
  NAND2_X1  g0820(.A1(new_n956), .A2(KEYINPUT111), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(new_n954), .Z(new_n1022));
  OAI211_X1 g0822(.A(new_n957), .B(new_n1016), .C1(new_n1022), .C2(new_n949), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n929), .A2(new_n774), .A3(new_n930), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n266), .B(new_n811), .C1(G143), .C2(new_n737), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n218), .B2(new_n755), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT113), .Z(new_n1027));
  AOI22_X1  g0827(.A1(G150), .A2(new_n748), .B1(new_n733), .B2(G159), .ZN(new_n1028));
  XOR2_X1   g0828(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n746), .A2(new_n212), .B1(new_n740), .B2(new_n294), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(G50), .C2(new_n728), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1027), .A2(new_n1031), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n266), .B1(new_n736), .B2(new_n1006), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n729), .A2(new_n751), .B1(new_n572), .B2(new_n746), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(G294), .C2(new_n817), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G317), .A2(new_n748), .B1(new_n733), .B2(G311), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT52), .Z(new_n1040));
  NAND2_X1  g0840(.A1(new_n761), .A2(G283), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1038), .A2(new_n764), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n725), .B1(new_n1035), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n251), .A2(new_n777), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n994), .B1(G97), .B2(new_n675), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n719), .B(new_n1043), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT114), .Z(new_n1047));
  AOI22_X1  g0847(.A1(new_n1022), .A2(new_n717), .B1(new_n1024), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1023), .A2(new_n1048), .ZN(G390));
  NAND2_X1  g0849(.A1(new_n910), .A2(new_n772), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n737), .A2(G125), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n259), .B1(new_n810), .B2(new_n207), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT117), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n1053), .B2(new_n1052), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT118), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G159), .A2(new_n747), .B1(new_n728), .B2(G137), .ZN(new_n1057));
  XOR2_X1   g0857(.A(KEYINPUT54), .B(G143), .Z(new_n1058));
  AOI22_X1  g0858(.A1(new_n733), .A2(G132), .B1(new_n817), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(G128), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1057), .B(new_n1059), .C1(new_n1060), .C2(new_n758), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n761), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT53), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n755), .B2(new_n296), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1061), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1056), .A2(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n758), .A2(new_n807), .B1(new_n212), .B2(new_n746), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G107), .B2(new_n728), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n266), .B1(new_n736), .B2(new_n812), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n732), .A2(new_n572), .B1(new_n740), .B2(new_n544), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(G68), .C2(new_n743), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1068), .B(new_n1071), .C1(new_n322), .C2(new_n755), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n725), .B1(new_n1066), .B2(new_n1072), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n719), .B(new_n1073), .C1(new_n294), .C2(new_n804), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1050), .A2(new_n1074), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1075), .A2(KEYINPUT119), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1075), .A2(KEYINPUT119), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n882), .B(G330), .C1(new_n706), .C2(new_n874), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n856), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n907), .B2(new_n870), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n692), .A2(new_n667), .A3(new_n792), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n899), .B1(new_n1083), .B2(new_n896), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n1082), .A2(new_n1084), .A3(new_n911), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n911), .B1(new_n897), .B2(new_n881), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n908), .A2(new_n909), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1080), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(KEYINPUT115), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1083), .A2(new_n896), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n881), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n873), .A2(new_n912), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n903), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n871), .B2(new_n872), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1086), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n909), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n711), .A2(G330), .A3(new_n792), .A4(new_n881), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1092), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT115), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1100), .B(new_n1080), .C1(new_n1085), .C2(new_n1087), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1089), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1078), .B1(new_n1102), .B2(new_n716), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT120), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1078), .B(KEYINPUT120), .C1(new_n1102), .C2(new_n716), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1016), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n462), .A2(new_n875), .A3(G330), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n914), .A2(new_n1108), .A3(new_n637), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1090), .ZN(new_n1111));
  OAI211_X1 g0911(.A(G330), .B(new_n792), .C1(new_n706), .C2(new_n874), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n899), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1098), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(G330), .B(new_n792), .C1(new_n706), .C2(new_n709), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n899), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n898), .B1(new_n1079), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1110), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1107), .B1(new_n1102), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1079), .A2(new_n1117), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n897), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1109), .B1(new_n1122), .B2(new_n1114), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1089), .A2(new_n1099), .A3(new_n1101), .A4(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(KEYINPUT116), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1101), .A2(new_n1099), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1092), .A2(new_n1097), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1100), .B1(new_n1127), .B2(new_n1080), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1119), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  AND4_X1   g0929(.A1(KEYINPUT116), .A2(new_n1129), .A3(new_n1016), .A4(new_n1124), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1105), .B(new_n1106), .C1(new_n1125), .C2(new_n1130), .ZN(G378));
  NAND3_X1  g0931(.A1(new_n883), .A2(G330), .A3(new_n889), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n309), .A2(new_n345), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n302), .A2(new_n850), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1133), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1138), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1133), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1140), .A2(new_n1136), .A3(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1132), .A2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1143), .B(KEYINPUT121), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1145), .A2(new_n883), .A3(G330), .A4(new_n889), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1144), .A2(new_n1146), .A3(new_n913), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n913), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n717), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n758), .A2(new_n572), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n972), .B(new_n1151), .C1(G97), .C2(new_n728), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n465), .A2(new_n817), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n259), .A2(G41), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1154), .B1(new_n807), .B2(new_n736), .C1(new_n312), .C2(new_n732), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G58), .B2(new_n743), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1152), .A2(new_n999), .A3(new_n1153), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT58), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1154), .ZN(new_n1159));
  AOI21_X1  g0959(.A(G50), .B1(new_n256), .B2(new_n273), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1157), .A2(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n1158), .B2(new_n1157), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n761), .A2(new_n1058), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n732), .A2(new_n1060), .B1(new_n740), .B2(new_n819), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G132), .B2(new_n728), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G150), .A2(new_n747), .B1(new_n748), .B2(G125), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1163), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1167), .A2(KEYINPUT59), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(KEYINPUT59), .ZN(new_n1169));
  AOI211_X1 g0969(.A(G33), .B(G41), .C1(new_n737), .C2(G124), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n407), .B2(new_n810), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n724), .B1(new_n1162), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n719), .B1(new_n207), .B2(new_n804), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(new_n1145), .C2(new_n773), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1150), .A2(new_n1175), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n1126), .A2(new_n1128), .A3(new_n1119), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1109), .B(KEYINPUT122), .Z(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(KEYINPUT123), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT123), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1124), .A2(new_n1181), .A3(new_n1178), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT57), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1147), .A2(new_n1148), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1107), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1124), .A2(new_n1181), .A3(new_n1178), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1181), .B1(new_n1124), .B2(new_n1178), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1149), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1184), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1176), .B1(new_n1186), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(G375));
  NOR3_X1   g0992(.A1(new_n1110), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1193), .A2(new_n944), .A3(new_n1123), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT124), .Z(new_n1195));
  OAI21_X1  g0995(.A(new_n718), .B1(G68), .B2(new_n805), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n728), .A2(new_n1058), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n207), .B2(new_n746), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G132), .B2(new_n748), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n259), .B1(new_n740), .B2(new_n296), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n732), .A2(new_n819), .B1(new_n736), .B2(new_n1060), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(G58), .C2(new_n743), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1199), .B(new_n1202), .C1(new_n407), .C2(new_n755), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n572), .A2(new_n729), .B1(new_n758), .B2(new_n812), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n266), .B1(new_n740), .B2(new_n312), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n732), .A2(new_n807), .B1(new_n736), .B2(new_n751), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1207), .A2(new_n976), .A3(new_n996), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n755), .A2(new_n544), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1203), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1196), .B1(new_n1210), .B2(new_n724), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n881), .B2(new_n773), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1212), .B1(new_n1213), .B2(new_n716), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1195), .A2(new_n1214), .ZN(G381));
  INV_X1    g1015(.A(G390), .ZN(new_n1216));
  INV_X1    g1016(.A(G387), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n828), .A3(new_n1217), .ZN(new_n1218));
  NOR4_X1   g1018(.A1(new_n1218), .A2(G381), .A3(G396), .A4(G393), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1105), .A2(new_n1220), .A3(new_n1106), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1219), .A2(new_n1191), .A3(new_n1222), .ZN(G407));
  NAND2_X1  g1023(.A1(new_n658), .A2(G213), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1191), .A2(new_n1222), .A3(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(G407), .A2(G213), .A3(new_n1226), .ZN(G409));
  INV_X1    g1027(.A(G2897), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1224), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT125), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1213), .A2(new_n1109), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT60), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1231), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1193), .A2(KEYINPUT125), .A3(KEYINPUT60), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1107), .B(new_n1123), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1214), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(G384), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(G384), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1230), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1238), .A2(G384), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1214), .B(new_n828), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1242), .A2(new_n1243), .A3(new_n1229), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1150), .A2(new_n1175), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n944), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1247), .B(new_n1149), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1221), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1191), .B2(G378), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1245), .B1(new_n1250), .B2(new_n1225), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT57), .B1(new_n1183), .B2(new_n1149), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1185), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1016), .ZN(new_n1254));
  OAI211_X1 g1054(.A(G378), .B(new_n1246), .C1(new_n1252), .C2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1222), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT62), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1224), .A4(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT61), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1251), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1225), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1259), .B1(new_n1264), .B2(new_n1260), .ZN(new_n1265));
  OAI21_X1  g1065(.A(KEYINPUT127), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1265), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1258), .A2(new_n1224), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT61), .B1(new_n1268), .B2(new_n1245), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT127), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1267), .A2(new_n1269), .A3(new_n1270), .A4(new_n1261), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1216), .A2(G387), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1217), .A2(G390), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(G393), .B(new_n786), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1275), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1266), .A2(new_n1271), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1264), .A2(new_n1260), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT63), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1276), .A2(new_n1262), .A3(new_n1278), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT126), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1283), .B1(new_n1284), .B2(new_n1251), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1268), .A2(KEYINPUT126), .A3(new_n1245), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1282), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1280), .A2(new_n1287), .ZN(G405));
  OAI21_X1  g1088(.A(new_n1255), .B1(new_n1191), .B2(new_n1221), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1289), .A2(new_n1260), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1260), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  XOR2_X1   g1092(.A(new_n1292), .B(new_n1279), .Z(G402));
endmodule


