//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n536, new_n538,
    new_n539, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n551, new_n552, new_n553, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n581,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1145, new_n1146, new_n1148;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n462), .A2(new_n464), .A3(G137), .A4(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n468), .B1(G2105), .B2(new_n471), .ZN(G160));
  AND3_X1   g047(.A1(new_n462), .A2(new_n464), .A3(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n465), .A2(G112), .ZN(new_n475));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n465), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n477), .B1(G136), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT67), .ZN(G162));
  NAND4_X1  g057(.A1(new_n462), .A2(new_n464), .A3(G138), .A4(new_n465), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n483), .B(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT69), .B1(new_n465), .B2(G114), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(new_n488), .A3(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g068(.A1(G126), .A2(G2105), .ZN(new_n494));
  AOI21_X1  g069(.A(KEYINPUT68), .B1(new_n478), .B2(new_n494), .ZN(new_n495));
  AND4_X1   g070(.A1(KEYINPUT68), .A2(new_n462), .A3(new_n464), .A4(new_n494), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n485), .A2(new_n497), .ZN(G164));
  NAND2_X1  g073(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  XNOR2_X1  g075(.A(new_n499), .B(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(G543), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n504), .A2(new_n510), .ZN(G303));
  INV_X1    g086(.A(G303), .ZN(G166));
  INV_X1    g087(.A(new_n506), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n513), .A2(G89), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  INV_X1    g092(.A(G51), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n515), .B(new_n517), .C1(new_n518), .C2(new_n509), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n514), .A2(new_n519), .ZN(G286));
  INV_X1    g095(.A(G286), .ZN(G168));
  AOI22_X1  g096(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n522), .A2(new_n503), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT72), .B(G90), .ZN(new_n524));
  INV_X1    g099(.A(G52), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n506), .A2(new_n524), .B1(new_n525), .B2(new_n509), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(G171));
  AOI22_X1  g102(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n503), .ZN(new_n529));
  INV_X1    g104(.A(G81), .ZN(new_n530));
  INV_X1    g105(.A(G43), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n506), .A2(new_n530), .B1(new_n531), .B2(new_n509), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G860), .ZN(new_n534));
  XOR2_X1   g109(.A(new_n534), .B(KEYINPUT73), .Z(G153));
  AND3_X1   g110(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G36), .ZN(G176));
  NAND2_X1  g112(.A1(G1), .A2(G3), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT8), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n539), .ZN(G188));
  NAND3_X1  g115(.A1(new_n505), .A2(G53), .A3(G543), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT9), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(KEYINPUT74), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n541), .A2(new_n543), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n544), .A2(new_n545), .B1(new_n513), .B2(G91), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n501), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n503), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(G299));
  INV_X1    g124(.A(G171), .ZN(G301));
  INV_X1    g125(.A(new_n509), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n513), .A2(G87), .B1(G49), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g127(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(G288));
  NAND2_X1  g129(.A1(new_n551), .A2(G48), .ZN(new_n555));
  INV_X1    g130(.A(G86), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n556), .B2(new_n506), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n501), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(new_n503), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(G305));
  NAND2_X1  g136(.A1(G72), .A2(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n499), .B(G543), .ZN(new_n563));
  INV_X1    g138(.A(G60), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n503), .B1(new_n565), .B2(KEYINPUT75), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n566), .B1(KEYINPUT75), .B2(new_n565), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT76), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n513), .A2(G85), .B1(G47), .B2(new_n551), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(G290));
  NAND2_X1  g145(.A1(G301), .A2(G868), .ZN(new_n571));
  AND3_X1   g146(.A1(new_n501), .A2(G92), .A3(new_n505), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT10), .ZN(new_n573));
  NAND2_X1  g148(.A1(G79), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G66), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n563), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(new_n551), .B2(G54), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n571), .B1(new_n578), .B2(G868), .ZN(G284));
  OAI21_X1  g154(.A(new_n571), .B1(new_n578), .B2(G868), .ZN(G321));
  XOR2_X1   g155(.A(G299), .B(KEYINPUT77), .Z(new_n581));
  MUX2_X1   g156(.A(new_n581), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g157(.A(new_n581), .B(G286), .S(G868), .Z(G280));
  INV_X1    g158(.A(G559), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n578), .B1(new_n584), .B2(G860), .ZN(G148));
  NAND2_X1  g160(.A1(new_n578), .A2(new_n584), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G868), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(KEYINPUT78), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(KEYINPUT78), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n588), .B(new_n589), .C1(G868), .C2(new_n533), .ZN(G323));
  XOR2_X1   g165(.A(KEYINPUT79), .B(KEYINPUT11), .Z(new_n591));
  XNOR2_X1  g166(.A(G323), .B(new_n591), .ZN(G282));
  NAND2_X1  g167(.A1(new_n480), .A2(G2104), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT12), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT13), .ZN(new_n595));
  INV_X1    g170(.A(G2100), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n473), .A2(G123), .ZN(new_n599));
  INV_X1    g174(.A(G135), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n465), .A2(G111), .ZN(new_n601));
  OAI21_X1  g176(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n602));
  OAI221_X1 g177(.A(new_n599), .B1(new_n600), .B2(new_n479), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(G2096), .Z(new_n604));
  NAND3_X1  g179(.A1(new_n597), .A2(new_n598), .A3(new_n604), .ZN(G156));
  XNOR2_X1  g180(.A(G2427), .B(G2438), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(G2430), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT15), .B(G2435), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n609), .A2(KEYINPUT14), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(G1341), .B(G1348), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n611), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(G2451), .B(G2454), .ZN(new_n616));
  XNOR2_X1  g191(.A(G2443), .B(G2446), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n616), .B(new_n617), .Z(new_n618));
  OR2_X1    g193(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n615), .A2(new_n618), .ZN(new_n620));
  AND3_X1   g195(.A1(new_n619), .A2(G14), .A3(new_n620), .ZN(G401));
  XOR2_X1   g196(.A(G2072), .B(G2078), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT81), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT17), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2067), .B(G2678), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2084), .B(G2090), .ZN(new_n626));
  NOR3_X1   g201(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n623), .B2(new_n625), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n624), .B2(new_n625), .ZN(new_n629));
  INV_X1    g204(.A(new_n625), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n630), .A2(new_n626), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT18), .ZN(new_n633));
  NOR3_X1   g208(.A1(new_n627), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2096), .B(G2100), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(G227));
  XOR2_X1   g211(.A(G1971), .B(G1976), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT19), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1956), .B(G2474), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1961), .B(G1966), .ZN(new_n640));
  AND2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  NOR3_X1   g218(.A1(new_n638), .A2(new_n643), .A3(new_n641), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n638), .A2(new_n643), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n646));
  AOI211_X1 g221(.A(new_n642), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n645), .B2(new_n646), .ZN(new_n648));
  XOR2_X1   g223(.A(G1991), .B(G1996), .Z(new_n649));
  XOR2_X1   g224(.A(new_n648), .B(new_n649), .Z(new_n650));
  XNOR2_X1  g225(.A(G1981), .B(G1986), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT83), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n650), .B(new_n654), .ZN(G229));
  INV_X1    g230(.A(G16), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(G20), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT23), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(G299), .B2(G16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT95), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G1956), .ZN(new_n661));
  NOR2_X1   g236(.A1(G168), .A2(new_n656), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n656), .B2(G21), .ZN(new_n663));
  INV_X1    g238(.A(G1966), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT31), .B(G11), .ZN(new_n666));
  INV_X1    g241(.A(G29), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT30), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n667), .B1(new_n668), .B2(G28), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n669), .A2(KEYINPUT91), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(G28), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n669), .B2(KEYINPUT91), .ZN(new_n672));
  OAI221_X1 g247(.A(new_n666), .B1(new_n670), .B2(new_n672), .C1(new_n603), .C2(new_n667), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n656), .A2(G5), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(G171), .B2(new_n656), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n673), .B1(new_n675), .B2(G1961), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n663), .A2(new_n664), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n665), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT92), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n667), .A2(G26), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT88), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  OR2_X1    g257(.A1(G104), .A2(G2105), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n683), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n684));
  INV_X1    g259(.A(G140), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n479), .B2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT87), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n478), .A2(G2105), .ZN(new_n688));
  INV_X1    g263(.A(G128), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n473), .A2(KEYINPUT87), .A3(G128), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n686), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n682), .B1(new_n693), .B2(G29), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G2067), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n667), .A2(G33), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT25), .Z(new_n698));
  INV_X1    g273(.A(G139), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(new_n479), .ZN(new_n700));
  AOI22_X1  g275(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n701), .A2(new_n465), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT89), .Z(new_n704));
  OAI21_X1  g279(.A(new_n696), .B1(new_n704), .B2(new_n667), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n695), .B1(new_n705), .B2(G2072), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n667), .A2(G35), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G162), .B2(new_n667), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G2090), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI211_X1 g287(.A(new_n706), .B(new_n712), .C1(G2072), .C2(new_n705), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT26), .Z(new_n715));
  INV_X1    g290(.A(G129), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n688), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n718));
  INV_X1    g293(.A(G141), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n479), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(new_n667), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n667), .B2(G32), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT27), .B(G1996), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(G160), .A2(G29), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT90), .B(KEYINPUT24), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G34), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n726), .B1(G29), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n725), .B1(G2084), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n656), .A2(G19), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n533), .B2(new_n656), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(G1341), .Z(new_n734));
  INV_X1    g309(.A(G2084), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n723), .A2(new_n724), .B1(new_n735), .B2(new_n729), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n731), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G27), .A2(G29), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G164), .B2(G29), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT93), .B(G2078), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G1961), .B2(new_n675), .ZN(new_n742));
  NOR2_X1   g317(.A1(G4), .A2(G16), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n578), .B2(G16), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1348), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n737), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n679), .A2(new_n713), .A3(new_n746), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n661), .B(new_n747), .C1(new_n711), .C2(new_n710), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n473), .A2(G119), .ZN(new_n749));
  INV_X1    g324(.A(G131), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n465), .A2(G107), .ZN(new_n751));
  OAI21_X1  g326(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n749), .B1(new_n750), .B2(new_n479), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  MUX2_X1   g328(.A(G25), .B(new_n753), .S(G29), .Z(new_n754));
  XOR2_X1   g329(.A(KEYINPUT35), .B(G1991), .Z(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n754), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n656), .A2(G24), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT84), .Z(new_n759));
  INV_X1    g334(.A(G290), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(new_n656), .ZN(new_n761));
  INV_X1    g336(.A(G1986), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n656), .A2(G22), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G166), .B2(new_n656), .ZN(new_n765));
  INV_X1    g340(.A(G1971), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n656), .A2(G23), .ZN(new_n768));
  INV_X1    g343(.A(G288), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(new_n656), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT33), .B(G1976), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT85), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n770), .B(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G6), .A2(G16), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n560), .B2(G16), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT32), .B(G1981), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n767), .A2(new_n773), .A3(new_n777), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n778), .A2(KEYINPUT34), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n763), .A2(new_n779), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n757), .B(new_n780), .C1(KEYINPUT34), .C2(new_n778), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT86), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n781), .A2(new_n782), .A3(KEYINPUT36), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT86), .B(KEYINPUT36), .Z(new_n784));
  OR2_X1    g359(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n748), .A2(new_n783), .A3(new_n785), .ZN(G150));
  INV_X1    g361(.A(G150), .ZN(G311));
  NAND2_X1  g362(.A1(new_n578), .A2(G559), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT38), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(new_n503), .ZN(new_n791));
  INV_X1    g366(.A(G93), .ZN(new_n792));
  INV_X1    g367(.A(G55), .ZN(new_n793));
  OAI22_X1  g368(.A1(new_n506), .A2(new_n792), .B1(new_n793), .B2(new_n509), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n533), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n533), .A2(new_n795), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n789), .B(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(KEYINPUT39), .ZN(new_n801));
  INV_X1    g376(.A(G860), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(KEYINPUT39), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n795), .A2(new_n802), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT37), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n806), .ZN(G145));
  XNOR2_X1  g382(.A(new_n594), .B(new_n753), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n693), .A2(G164), .ZN(new_n810));
  INV_X1    g385(.A(new_n484), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n483), .B(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n462), .A2(new_n464), .A3(new_n494), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT68), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n478), .A2(KEYINPUT68), .A3(new_n494), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n815), .A2(new_n816), .B1(new_n490), .B2(new_n492), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n692), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n810), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n721), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n810), .A2(new_n721), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(new_n704), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT96), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n822), .A2(new_n826), .A3(new_n823), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n826), .B1(new_n822), .B2(new_n823), .ZN(new_n829));
  OAI22_X1  g404(.A1(new_n828), .A2(new_n829), .B1(new_n702), .B2(new_n700), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n825), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n824), .A2(KEYINPUT96), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n703), .B1(new_n833), .B2(new_n827), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n834), .A2(KEYINPUT97), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n480), .A2(G142), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT98), .ZN(new_n837));
  OR2_X1    g412(.A1(G106), .A2(G2105), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n838), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n839));
  INV_X1    g414(.A(G130), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n688), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n832), .A2(new_n835), .A3(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n842), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n834), .A2(KEYINPUT97), .B1(new_n704), .B2(new_n824), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n830), .A2(new_n831), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n809), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n468), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n471), .A2(G2105), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n603), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(G162), .B(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n842), .B1(new_n832), .B2(new_n835), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n845), .A2(new_n846), .A3(new_n844), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n854), .A2(new_n808), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n848), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n848), .A2(KEYINPUT99), .A3(new_n853), .A4(new_n856), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n853), .B1(new_n848), .B2(new_n856), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n862), .A2(G37), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n861), .A2(KEYINPUT40), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT40), .B1(new_n861), .B2(new_n863), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(G395));
  NOR2_X1   g441(.A1(new_n578), .A2(G299), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT101), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n578), .A2(G299), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT100), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT102), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n798), .B(new_n586), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n868), .A2(KEYINPUT41), .A3(new_n870), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT41), .B1(new_n868), .B2(new_n870), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n874), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(G290), .B(new_n560), .ZN(new_n879));
  XNOR2_X1  g454(.A(G303), .B(G288), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT42), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n878), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(G868), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(G868), .B2(new_n795), .ZN(G295));
  OAI21_X1  g460(.A(new_n884), .B1(G868), .B2(new_n795), .ZN(G331));
  INV_X1    g461(.A(new_n881), .ZN(new_n887));
  NAND2_X1  g462(.A1(G301), .A2(KEYINPUT103), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n889));
  NAND2_X1  g464(.A1(G171), .A2(new_n889), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n888), .A2(G168), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(G168), .B1(new_n888), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n799), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n798), .B1(new_n891), .B2(new_n892), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n875), .B2(new_n876), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n898), .A3(new_n895), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n893), .A2(KEYINPUT104), .A3(new_n799), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n871), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n887), .A2(new_n897), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n897), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n881), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT43), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n901), .B1(new_n910), .B2(new_n875), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n877), .A2(KEYINPUT105), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n872), .A2(new_n895), .A3(new_n894), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n887), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n915), .A2(new_n905), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT44), .B1(new_n909), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n916), .B1(new_n906), .B2(new_n908), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n915), .A2(new_n905), .A3(KEYINPUT43), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n918), .B1(new_n921), .B2(KEYINPUT44), .ZN(G397));
  NAND3_X1  g497(.A1(new_n849), .A2(new_n850), .A3(G40), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT106), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n925));
  NAND3_X1  g500(.A1(G160), .A2(new_n925), .A3(G40), .ZN(new_n926));
  AOI21_X1  g501(.A(G1384), .B1(new_n812), .B2(new_n817), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT50), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n924), .B(new_n926), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G1384), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n485), .B2(new_n497), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n931), .A2(KEYINPUT50), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(KEYINPUT108), .A3(new_n711), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n924), .A2(new_n926), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n927), .A2(new_n928), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n931), .A2(KEYINPUT50), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n935), .A2(new_n711), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n924), .B(new_n926), .C1(new_n927), .C2(KEYINPUT45), .ZN(new_n941));
  OAI211_X1 g516(.A(KEYINPUT45), .B(new_n930), .C1(new_n485), .C2(new_n497), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n934), .B(new_n940), .C1(G1971), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(G303), .A2(G8), .ZN(new_n946));
  XNOR2_X1  g521(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n946), .B(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(G8), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT49), .ZN(new_n950));
  INV_X1    g525(.A(new_n559), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n513), .A2(G86), .ZN(new_n952));
  XOR2_X1   g527(.A(KEYINPUT110), .B(G1981), .Z(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n951), .A2(new_n952), .A3(new_n555), .A4(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G1981), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n560), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n950), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n924), .A2(new_n927), .A3(new_n926), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G8), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n955), .B(KEYINPUT49), .C1(new_n560), .C2(new_n957), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n959), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n769), .A2(G1976), .ZN(new_n966));
  INV_X1    g541(.A(G1976), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT52), .B1(G288), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n963), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(G8), .A3(new_n960), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT52), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n965), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n949), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n942), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n818), .A2(KEYINPUT112), .A3(KEYINPUT45), .A4(new_n930), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n664), .B1(new_n977), .B2(new_n941), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n935), .A2(new_n735), .A3(new_n936), .A4(new_n937), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n962), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(G168), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT63), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n944), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n984), .A2(new_n766), .B1(new_n938), .B2(new_n939), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n962), .B1(new_n985), .B2(new_n934), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n948), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(new_n986), .B2(new_n987), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n973), .B(new_n983), .C1(new_n988), .C2(new_n990), .ZN(new_n991));
  AOI22_X1  g566(.A1(new_n984), .A2(new_n766), .B1(new_n933), .B2(new_n711), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n989), .B1(new_n992), .B2(new_n962), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n949), .A2(new_n993), .A3(new_n972), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n982), .B1(new_n994), .B2(new_n981), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n965), .A2(new_n967), .A3(new_n769), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n963), .B1(new_n996), .B2(new_n956), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n986), .A2(new_n972), .A3(new_n948), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT111), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n991), .A2(new_n995), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G286), .A2(G8), .ZN(new_n1004));
  XOR2_X1   g579(.A(new_n1004), .B(KEYINPUT118), .Z(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(new_n980), .B2(KEYINPUT119), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n1007));
  AOI211_X1 g582(.A(new_n1007), .B(new_n962), .C1(new_n978), .C2(new_n979), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT51), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT120), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT120), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1011), .B(KEYINPUT51), .C1(new_n1006), .C2(new_n1008), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1010), .A2(new_n978), .A3(new_n979), .A4(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n980), .A2(KEYINPUT51), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1005), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G2078), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n931), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n935), .A2(new_n1018), .A3(new_n1020), .A4(new_n942), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1022));
  NAND3_X1  g597(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n1023));
  INV_X1    g598(.A(G1961), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n1021), .A2(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT123), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n927), .A2(KEYINPUT45), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1026), .B1(new_n1027), .B2(new_n923), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1020), .A2(KEYINPUT123), .A3(G40), .A4(G160), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1031));
  AND2_X1   g606(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n942), .B(KEYINPUT53), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT125), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT125), .ZN(new_n1036));
  AOI211_X1 g611(.A(new_n1036), .B(new_n1033), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1025), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT126), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g615(.A(KEYINPUT126), .B(new_n1025), .C1(new_n1035), .C2(new_n1037), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(G171), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1025), .ZN(new_n1044));
  INV_X1    g619(.A(new_n941), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1045), .A2(new_n1018), .A3(new_n976), .A4(new_n975), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT121), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1044), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1043), .B1(new_n1051), .B2(G301), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n994), .B1(new_n1042), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT114), .B1(new_n544), .B2(new_n545), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(KEYINPUT57), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G299), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n546), .B(new_n548), .C1(new_n1054), .C2(KEYINPUT57), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1956), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(new_n929), .B2(new_n932), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n1061));
  XNOR2_X1  g636(.A(new_n1061), .B(G2072), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n935), .A2(new_n1020), .A3(new_n942), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1058), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1060), .A2(new_n1063), .A3(new_n1058), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n578), .ZN(new_n1067));
  INV_X1    g642(.A(G1348), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1023), .A2(new_n1068), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n960), .A2(G2067), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1064), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT61), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n1065), .B2(new_n1064), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1996), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n935), .A2(new_n1077), .A3(new_n1020), .A4(new_n942), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT58), .B(G1341), .Z(new_n1079));
  NAND2_X1  g654(.A1(new_n960), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n533), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT116), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(new_n1084), .A3(new_n533), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(KEYINPUT59), .A3(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(KEYINPUT117), .B(new_n1073), .C1(new_n1065), .C2(new_n1064), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1084), .B1(new_n1081), .B2(new_n533), .ZN(new_n1089));
  INV_X1    g664(.A(new_n533), .ZN(new_n1090));
  AOI211_X1 g665(.A(KEYINPUT116), .B(new_n1090), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1088), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1076), .A2(new_n1086), .A3(new_n1087), .A4(new_n1092), .ZN(new_n1093));
  OR3_X1    g668(.A1(new_n1065), .A2(new_n1064), .A3(new_n1073), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1069), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT60), .B1(new_n1095), .B2(new_n1071), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1069), .A2(new_n1097), .A3(new_n578), .A4(new_n1070), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1072), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g675(.A(G301), .B(new_n1025), .C1(new_n1035), .C2(new_n1037), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1051), .B2(G301), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1043), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1053), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1003), .B1(new_n1017), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT127), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1017), .A2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(KEYINPUT62), .B(new_n1013), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n994), .A2(G301), .A3(new_n1051), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1003), .B(KEYINPUT127), .C1(new_n1017), .C2(new_n1104), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1107), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n924), .A2(new_n926), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(new_n1020), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n721), .B(G1996), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n692), .B(G2067), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n753), .B(new_n755), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1117), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n760), .A2(new_n762), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1124), .A2(KEYINPUT107), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n760), .A2(new_n762), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1117), .B1(new_n1124), .B2(KEYINPUT107), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1123), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1114), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1117), .B1(new_n721), .B2(new_n1119), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1116), .A2(KEYINPUT46), .A3(new_n1077), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT46), .B1(new_n1116), .B2(new_n1077), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT47), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1123), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1126), .A2(new_n1117), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1136), .B1(new_n1137), .B2(KEYINPUT48), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1138), .B1(KEYINPUT48), .B2(new_n1137), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n753), .A2(new_n756), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1120), .A2(new_n1140), .B1(G2067), .B2(new_n693), .ZN(new_n1141));
  AOI211_X1 g716(.A(new_n1135), .B(new_n1139), .C1(new_n1116), .C2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1130), .A2(new_n1142), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g718(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1145));
  OAI21_X1  g719(.A(new_n1145), .B1(new_n919), .B2(new_n920), .ZN(new_n1146));
  AOI21_X1  g720(.A(new_n1146), .B1(new_n861), .B2(new_n863), .ZN(G308));
  NAND2_X1  g721(.A1(new_n861), .A2(new_n863), .ZN(new_n1148));
  OAI211_X1 g722(.A(new_n1148), .B(new_n1145), .C1(new_n919), .C2(new_n920), .ZN(G225));
endmodule


