

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  XNOR2_X1 U324 ( .A(n354), .B(n353), .ZN(n356) );
  AND2_X1 U325 ( .A1(n399), .A2(n398), .ZN(n401) );
  INV_X1 U326 ( .A(KEYINPUT115), .ZN(n400) );
  NOR2_X1 U327 ( .A1(n452), .A2(n543), .ZN(n453) );
  XNOR2_X1 U328 ( .A(n396), .B(n292), .ZN(n366) );
  XNOR2_X1 U329 ( .A(n352), .B(KEYINPUT8), .ZN(n353) );
  NOR2_X1 U330 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U331 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U332 ( .A(n401), .B(n400), .ZN(n411) );
  XNOR2_X1 U333 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U334 ( .A(n394), .B(n393), .ZN(n395) );
  AND2_X1 U335 ( .A1(n570), .A2(n550), .ZN(n457) );
  XNOR2_X1 U336 ( .A(n436), .B(n421), .ZN(n292) );
  XOR2_X1 U337 ( .A(G113GAT), .B(G197GAT), .Z(n293) );
  XOR2_X1 U338 ( .A(KEYINPUT54), .B(n413), .Z(n294) );
  XNOR2_X1 U339 ( .A(n402), .B(KEYINPUT113), .ZN(n403) );
  XNOR2_X1 U340 ( .A(n404), .B(n403), .ZN(n407) );
  XNOR2_X1 U341 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n408) );
  XOR2_X1 U342 ( .A(G1GAT), .B(G15GAT), .Z(n388) );
  XNOR2_X1 U343 ( .A(n359), .B(KEYINPUT10), .ZN(n360) );
  INV_X1 U344 ( .A(G29GAT), .ZN(n352) );
  XNOR2_X1 U345 ( .A(n368), .B(n360), .ZN(n364) );
  NOR2_X1 U346 ( .A1(n528), .A2(n294), .ZN(n414) );
  XNOR2_X1 U347 ( .A(n427), .B(n293), .ZN(n393) );
  XOR2_X1 U348 ( .A(KEYINPUT36), .B(n550), .Z(n588) );
  XNOR2_X1 U349 ( .A(n366), .B(n365), .ZN(n405) );
  XNOR2_X1 U350 ( .A(n383), .B(n382), .ZN(n580) );
  XNOR2_X1 U351 ( .A(n453), .B(KEYINPUT122), .ZN(n570) );
  XNOR2_X1 U352 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U353 ( .A(n460), .B(n459), .ZN(G1349GAT) );
  XOR2_X1 U354 ( .A(G85GAT), .B(G162GAT), .Z(n296) );
  XNOR2_X1 U355 ( .A(G29GAT), .B(G134GAT), .ZN(n295) );
  XNOR2_X1 U356 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U357 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n298) );
  XNOR2_X1 U358 ( .A(KEYINPUT90), .B(G57GAT), .ZN(n297) );
  XNOR2_X1 U359 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U360 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U361 ( .A(KEYINPUT5), .B(G148GAT), .Z(n302) );
  NAND2_X1 U362 ( .A1(G225GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U363 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U364 ( .A(KEYINPUT4), .B(n303), .ZN(n304) );
  XNOR2_X1 U365 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U366 ( .A(KEYINPUT91), .B(G120GAT), .Z(n307) );
  XNOR2_X1 U367 ( .A(G141GAT), .B(G1GAT), .ZN(n306) );
  XNOR2_X1 U368 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U369 ( .A(n309), .B(n308), .Z(n314) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n310), .B(G127GAT), .ZN(n439) );
  XOR2_X1 U372 ( .A(G155GAT), .B(KEYINPUT3), .Z(n312) );
  XNOR2_X1 U373 ( .A(KEYINPUT2), .B(KEYINPUT88), .ZN(n311) );
  XNOR2_X1 U374 ( .A(n312), .B(n311), .ZN(n426) );
  XNOR2_X1 U375 ( .A(n439), .B(n426), .ZN(n313) );
  XNOR2_X1 U376 ( .A(n314), .B(n313), .ZN(n528) );
  INV_X1 U377 ( .A(G204GAT), .ZN(n315) );
  NAND2_X1 U378 ( .A1(G64GAT), .A2(n315), .ZN(n318) );
  INV_X1 U379 ( .A(G64GAT), .ZN(n316) );
  NAND2_X1 U380 ( .A1(n316), .A2(G204GAT), .ZN(n317) );
  NAND2_X1 U381 ( .A1(n318), .A2(n317), .ZN(n320) );
  XNOR2_X1 U382 ( .A(G176GAT), .B(KEYINPUT74), .ZN(n319) );
  XNOR2_X1 U383 ( .A(n320), .B(n319), .ZN(n369) );
  XOR2_X1 U384 ( .A(KEYINPUT92), .B(G92GAT), .Z(n322) );
  NAND2_X1 U385 ( .A1(G226GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U386 ( .A(n322), .B(n321), .ZN(n325) );
  XOR2_X1 U387 ( .A(G211GAT), .B(KEYINPUT21), .Z(n324) );
  XNOR2_X1 U388 ( .A(G197GAT), .B(KEYINPUT87), .ZN(n323) );
  XNOR2_X1 U389 ( .A(n324), .B(n323), .ZN(n424) );
  XOR2_X1 U390 ( .A(n325), .B(n424), .Z(n329) );
  XOR2_X1 U391 ( .A(G183GAT), .B(KEYINPUT19), .Z(n327) );
  XNOR2_X1 U392 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n326) );
  XNOR2_X1 U393 ( .A(n327), .B(n326), .ZN(n435) );
  XNOR2_X1 U394 ( .A(G190GAT), .B(n435), .ZN(n328) );
  XNOR2_X1 U395 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U396 ( .A(n330), .B(G218GAT), .Z(n332) );
  XOR2_X1 U397 ( .A(G169GAT), .B(G8GAT), .Z(n386) );
  XNOR2_X1 U398 ( .A(G36GAT), .B(n386), .ZN(n331) );
  XNOR2_X1 U399 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U400 ( .A(n369), .B(n333), .Z(n490) );
  XOR2_X1 U401 ( .A(G211GAT), .B(G155GAT), .Z(n335) );
  XNOR2_X1 U402 ( .A(G127GAT), .B(G183GAT), .ZN(n334) );
  XNOR2_X1 U403 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U404 ( .A(n336), .B(G64GAT), .Z(n338) );
  XNOR2_X1 U405 ( .A(G8GAT), .B(n388), .ZN(n337) );
  XNOR2_X1 U406 ( .A(n338), .B(n337), .ZN(n343) );
  XNOR2_X1 U407 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n339) );
  XNOR2_X1 U408 ( .A(n339), .B(KEYINPUT71), .ZN(n377) );
  XOR2_X1 U409 ( .A(n377), .B(KEYINPUT12), .Z(n341) );
  NAND2_X1 U410 ( .A1(G231GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U411 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U412 ( .A(n343), .B(n342), .Z(n351) );
  XOR2_X1 U413 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n345) );
  XNOR2_X1 U414 ( .A(KEYINPUT81), .B(KEYINPUT79), .ZN(n344) );
  XNOR2_X1 U415 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U416 ( .A(G78GAT), .B(KEYINPUT80), .Z(n347) );
  XNOR2_X1 U417 ( .A(G22GAT), .B(G71GAT), .ZN(n346) );
  XNOR2_X1 U418 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U419 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U420 ( .A(n351), .B(n350), .ZN(n461) );
  XNOR2_X1 U421 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n354) );
  XNOR2_X1 U422 ( .A(G43GAT), .B(G50GAT), .ZN(n355) );
  XNOR2_X1 U423 ( .A(n356), .B(n355), .ZN(n396) );
  XOR2_X1 U424 ( .A(G190GAT), .B(G134GAT), .Z(n436) );
  XOR2_X1 U425 ( .A(G162GAT), .B(G218GAT), .Z(n421) );
  XOR2_X1 U426 ( .A(G106GAT), .B(G92GAT), .Z(n358) );
  XNOR2_X1 U427 ( .A(G99GAT), .B(G85GAT), .ZN(n357) );
  XNOR2_X1 U428 ( .A(n358), .B(n357), .ZN(n368) );
  AND2_X1 U429 ( .A1(G232GAT), .A2(G233GAT), .ZN(n359) );
  XOR2_X1 U430 ( .A(KEYINPUT11), .B(KEYINPUT77), .Z(n362) );
  XNOR2_X1 U431 ( .A(KEYINPUT9), .B(KEYINPUT65), .ZN(n361) );
  XNOR2_X1 U432 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U433 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U434 ( .A(n405), .B(KEYINPUT78), .ZN(n550) );
  NOR2_X1 U435 ( .A1(n461), .A2(n588), .ZN(n367) );
  XNOR2_X1 U436 ( .A(n367), .B(KEYINPUT45), .ZN(n399) );
  XNOR2_X1 U437 ( .A(n369), .B(n368), .ZN(n375) );
  XOR2_X1 U438 ( .A(KEYINPUT73), .B(KEYINPUT75), .Z(n371) );
  NAND2_X1 U439 ( .A1(G230GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U440 ( .A(n371), .B(n370), .ZN(n373) );
  INV_X1 U441 ( .A(KEYINPUT33), .ZN(n372) );
  XNOR2_X1 U442 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U443 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U444 ( .A(G148GAT), .B(G78GAT), .Z(n420) );
  XNOR2_X1 U445 ( .A(n376), .B(n420), .ZN(n383) );
  XOR2_X1 U446 ( .A(G120GAT), .B(G71GAT), .Z(n437) );
  XOR2_X1 U447 ( .A(n437), .B(n377), .Z(n381) );
  XOR2_X1 U448 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n379) );
  XNOR2_X1 U449 ( .A(KEYINPUT76), .B(KEYINPUT32), .ZN(n378) );
  XNOR2_X1 U450 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U451 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n385) );
  XNOR2_X1 U452 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n385), .B(n384), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n387), .B(n386), .ZN(n392) );
  XOR2_X1 U455 ( .A(n388), .B(KEYINPUT30), .Z(n390) );
  NAND2_X1 U456 ( .A1(G229GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U457 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n392), .B(n391), .ZN(n394) );
  XOR2_X1 U459 ( .A(G141GAT), .B(G22GAT), .Z(n427) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n577) );
  XNOR2_X1 U461 ( .A(n577), .B(KEYINPUT70), .ZN(n567) );
  INV_X1 U462 ( .A(n567), .ZN(n397) );
  AND2_X1 U463 ( .A1(n580), .A2(n397), .ZN(n398) );
  XNOR2_X1 U464 ( .A(KEYINPUT41), .B(n580), .ZN(n558) );
  NAND2_X1 U465 ( .A1(n577), .A2(n558), .ZN(n404) );
  INV_X1 U466 ( .A(KEYINPUT46), .ZN(n402) );
  INV_X1 U467 ( .A(n461), .ZN(n585) );
  NOR2_X1 U468 ( .A1(n405), .A2(n585), .ZN(n406) );
  NAND2_X1 U469 ( .A1(n407), .A2(n406), .ZN(n409) );
  XNOR2_X1 U470 ( .A(KEYINPUT48), .B(n412), .ZN(n538) );
  NOR2_X1 U471 ( .A1(n490), .A2(n538), .ZN(n413) );
  XOR2_X1 U472 ( .A(KEYINPUT64), .B(n414), .Z(n576) );
  XOR2_X1 U473 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n416) );
  XNOR2_X1 U474 ( .A(G204GAT), .B(KEYINPUT89), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n433) );
  XOR2_X1 U476 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n418) );
  NAND2_X1 U477 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U479 ( .A(KEYINPUT86), .B(n419), .ZN(n431) );
  XOR2_X1 U480 ( .A(n420), .B(G106GAT), .Z(n423) );
  XNOR2_X1 U481 ( .A(G50GAT), .B(n421), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U483 ( .A(n425), .B(n424), .Z(n429) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n473) );
  NOR2_X1 U488 ( .A1(n576), .A2(n473), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n434), .B(KEYINPUT55), .ZN(n452) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n443) );
  XOR2_X1 U492 ( .A(n439), .B(KEYINPUT82), .Z(n441) );
  NAND2_X1 U493 ( .A1(G227GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U495 ( .A(n443), .B(n442), .Z(n451) );
  XOR2_X1 U496 ( .A(G176GAT), .B(G99GAT), .Z(n445) );
  XNOR2_X1 U497 ( .A(G169GAT), .B(G43GAT), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U499 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n447) );
  XNOR2_X1 U500 ( .A(G15GAT), .B(KEYINPUT83), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U503 ( .A(n451), .B(n450), .ZN(n543) );
  XNOR2_X1 U504 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n455) );
  INV_X1 U505 ( .A(G190GAT), .ZN(n454) );
  XNOR2_X1 U506 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  NAND2_X1 U507 ( .A1(n558), .A2(n570), .ZN(n460) );
  XOR2_X1 U508 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n458) );
  XNOR2_X1 U509 ( .A(n458), .B(G176GAT), .ZN(n459) );
  XOR2_X1 U510 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n488) );
  NAND2_X1 U511 ( .A1(n567), .A2(n580), .ZN(n504) );
  NOR2_X1 U512 ( .A1(n461), .A2(n550), .ZN(n462) );
  XNOR2_X1 U513 ( .A(n462), .B(KEYINPUT16), .ZN(n485) );
  XNOR2_X1 U514 ( .A(n490), .B(KEYINPUT93), .ZN(n463) );
  XNOR2_X1 U515 ( .A(n463), .B(KEYINPUT27), .ZN(n478) );
  NAND2_X1 U516 ( .A1(n528), .A2(n478), .ZN(n539) );
  XOR2_X1 U517 ( .A(KEYINPUT28), .B(KEYINPUT66), .Z(n464) );
  XOR2_X1 U518 ( .A(n473), .B(n464), .Z(n541) );
  NOR2_X1 U519 ( .A1(n539), .A2(n541), .ZN(n465) );
  XNOR2_X1 U520 ( .A(KEYINPUT94), .B(n465), .ZN(n466) );
  NAND2_X1 U521 ( .A1(n466), .A2(n543), .ZN(n467) );
  XOR2_X1 U522 ( .A(KEYINPUT95), .B(n467), .Z(n484) );
  INV_X1 U523 ( .A(n528), .ZN(n482) );
  XOR2_X1 U524 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n468) );
  XNOR2_X1 U525 ( .A(KEYINPUT25), .B(n468), .ZN(n472) );
  NOR2_X1 U526 ( .A1(n543), .A2(n490), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n469), .B(KEYINPUT98), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n473), .A2(n470), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n472), .B(n471), .ZN(n480) );
  XOR2_X1 U530 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n475) );
  NAND2_X1 U531 ( .A1(n543), .A2(n473), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U533 ( .A(KEYINPUT96), .B(n476), .ZN(n575) );
  INV_X1 U534 ( .A(n575), .ZN(n477) );
  NAND2_X1 U535 ( .A1(n478), .A2(n477), .ZN(n479) );
  NAND2_X1 U536 ( .A1(n480), .A2(n479), .ZN(n481) );
  NAND2_X1 U537 ( .A1(n482), .A2(n481), .ZN(n483) );
  NAND2_X1 U538 ( .A1(n484), .A2(n483), .ZN(n500) );
  NAND2_X1 U539 ( .A1(n485), .A2(n500), .ZN(n486) );
  XOR2_X1 U540 ( .A(KEYINPUT101), .B(n486), .Z(n515) );
  NOR2_X1 U541 ( .A1(n504), .A2(n515), .ZN(n497) );
  NAND2_X1 U542 ( .A1(n497), .A2(n528), .ZN(n487) );
  XNOR2_X1 U543 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U544 ( .A(G1GAT), .B(n489), .Z(G1324GAT) );
  XOR2_X1 U545 ( .A(G8GAT), .B(KEYINPUT103), .Z(n492) );
  INV_X1 U546 ( .A(n490), .ZN(n530) );
  NAND2_X1 U547 ( .A1(n497), .A2(n530), .ZN(n491) );
  XNOR2_X1 U548 ( .A(n492), .B(n491), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT105), .B(KEYINPUT35), .Z(n494) );
  INV_X1 U550 ( .A(n543), .ZN(n532) );
  NAND2_X1 U551 ( .A1(n497), .A2(n532), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n494), .B(n493), .ZN(n496) );
  XOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT104), .Z(n495) );
  XNOR2_X1 U554 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  NAND2_X1 U555 ( .A1(n541), .A2(n497), .ZN(n498) );
  XNOR2_X1 U556 ( .A(n498), .B(KEYINPUT106), .ZN(n499) );
  XNOR2_X1 U557 ( .A(G22GAT), .B(n499), .ZN(G1327GAT) );
  XNOR2_X1 U558 ( .A(KEYINPUT37), .B(KEYINPUT107), .ZN(n503) );
  NOR2_X1 U559 ( .A1(n585), .A2(n588), .ZN(n501) );
  NAND2_X1 U560 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U561 ( .A(n503), .B(n502), .ZN(n527) );
  NOR2_X1 U562 ( .A1(n527), .A2(n504), .ZN(n506) );
  XNOR2_X1 U563 ( .A(KEYINPUT108), .B(KEYINPUT38), .ZN(n505) );
  XNOR2_X1 U564 ( .A(n506), .B(n505), .ZN(n512) );
  NAND2_X1 U565 ( .A1(n528), .A2(n512), .ZN(n508) );
  XOR2_X1 U566 ( .A(G29GAT), .B(KEYINPUT39), .Z(n507) );
  XNOR2_X1 U567 ( .A(n508), .B(n507), .ZN(G1328GAT) );
  NAND2_X1 U568 ( .A1(n512), .A2(n530), .ZN(n509) );
  XNOR2_X1 U569 ( .A(G36GAT), .B(n509), .ZN(G1329GAT) );
  NAND2_X1 U570 ( .A1(n532), .A2(n512), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n510), .B(KEYINPUT40), .ZN(n511) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n511), .ZN(G1330GAT) );
  NAND2_X1 U573 ( .A1(n541), .A2(n512), .ZN(n513) );
  XNOR2_X1 U574 ( .A(n513), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n517) );
  INV_X1 U576 ( .A(n577), .ZN(n514) );
  NAND2_X1 U577 ( .A1(n514), .A2(n558), .ZN(n526) );
  NOR2_X1 U578 ( .A1(n515), .A2(n526), .ZN(n523) );
  NAND2_X1 U579 ( .A1(n523), .A2(n528), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(n518), .ZN(G1332GAT) );
  NAND2_X1 U582 ( .A1(n530), .A2(n523), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n519), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n521) );
  NAND2_X1 U585 ( .A1(n523), .A2(n532), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U587 ( .A(G71GAT), .B(n522), .ZN(G1334GAT) );
  XOR2_X1 U588 ( .A(G78GAT), .B(KEYINPUT43), .Z(n525) );
  NAND2_X1 U589 ( .A1(n523), .A2(n541), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n535) );
  NAND2_X1 U592 ( .A1(n528), .A2(n535), .ZN(n529) );
  XNOR2_X1 U593 ( .A(G85GAT), .B(n529), .ZN(G1336GAT) );
  NAND2_X1 U594 ( .A1(n530), .A2(n535), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n531), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U596 ( .A1(n532), .A2(n535), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n533), .B(KEYINPUT112), .ZN(n534) );
  XNOR2_X1 U598 ( .A(G99GAT), .B(n534), .ZN(G1338GAT) );
  NAND2_X1 U599 ( .A1(n541), .A2(n535), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n536), .B(KEYINPUT44), .ZN(n537) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n537), .ZN(G1339GAT) );
  NOR2_X1 U602 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U603 ( .A(n540), .B(KEYINPUT116), .Z(n555) );
  OR2_X1 U604 ( .A1(n541), .A2(n555), .ZN(n542) );
  NOR2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n551), .A2(n567), .ZN(n544) );
  XNOR2_X1 U607 ( .A(n544), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U609 ( .A1(n551), .A2(n558), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n548) );
  NAND2_X1 U612 ( .A1(n551), .A2(n585), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U618 ( .A(G134GAT), .B(n554), .ZN(G1343GAT) );
  XOR2_X1 U619 ( .A(G141GAT), .B(KEYINPUT119), .Z(n557) );
  NOR2_X1 U620 ( .A1(n555), .A2(n575), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n563), .A2(n577), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n560) );
  NAND2_X1 U624 ( .A1(n563), .A2(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(n561), .ZN(G1345GAT) );
  NAND2_X1 U627 ( .A1(n585), .A2(n563), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n565) );
  NAND2_X1 U630 ( .A1(n563), .A2(n405), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G162GAT), .B(n566), .ZN(G1347GAT) );
  XOR2_X1 U633 ( .A(G169GAT), .B(KEYINPUT123), .Z(n569) );
  NAND2_X1 U634 ( .A1(n567), .A2(n570), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1348GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n585), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n573) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(n574), .Z(n579) );
  NOR2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n584) );
  NAND2_X1 U643 ( .A1(n584), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n582) );
  INV_X1 U646 ( .A(n584), .ZN(n587) );
  OR2_X1 U647 ( .A1(n587), .A2(n580), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U649 ( .A(G204GAT), .B(n583), .Z(G1353GAT) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(n589), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

