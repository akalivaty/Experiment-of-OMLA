//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G227), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT79), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  OR2_X1    g013(.A1(KEYINPUT0), .A2(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT0), .A3(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G107), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n208), .A2(KEYINPUT3), .A3(G104), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT3), .B1(new_n208), .B2(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT80), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n208), .A2(G104), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n206), .B2(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n208), .A2(KEYINPUT3), .A3(G104), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT80), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n213), .A2(G101), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n205), .B1(new_n220), .B2(KEYINPUT4), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT82), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n224));
  INV_X1    g038(.A(G101), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n225), .B(new_n207), .C1(new_n209), .C2(new_n210), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT81), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n224), .B1(new_n220), .B2(new_n228), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n213), .A2(new_n227), .A3(new_n219), .A4(G101), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n223), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(G101), .B1(new_n218), .B2(KEYINPUT80), .ZN(new_n232));
  AOI211_X1 g046(.A(new_n212), .B(new_n214), .C1(new_n216), .C2(new_n217), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n228), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n234), .A2(new_n230), .A3(new_n223), .A4(KEYINPUT4), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n222), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT87), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT83), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n207), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n206), .A2(KEYINPUT83), .A3(G107), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n240), .B(new_n241), .C1(new_n206), .C2(G107), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G101), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n243), .A2(new_n226), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT85), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n195), .A2(new_n245), .A3(KEYINPUT1), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G128), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n245), .B1(new_n195), .B2(KEYINPUT1), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n198), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT84), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n202), .A2(G128), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n252), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n254), .A2(KEYINPUT84), .A3(G128), .A4(new_n202), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n249), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n244), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT10), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n252), .B2(new_n195), .ZN(new_n261));
  OAI22_X1  g075(.A1(new_n261), .A2(new_n202), .B1(new_n251), .B2(new_n252), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n244), .A2(new_n262), .A3(KEYINPUT10), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n237), .A2(new_n238), .A3(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n234), .A2(new_n230), .A3(KEYINPUT4), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT82), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n221), .B1(new_n267), .B2(new_n235), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n259), .A2(new_n263), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT87), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G134), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G137), .ZN(new_n272));
  INV_X1    g086(.A(G137), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT64), .B1(new_n273), .B2(G134), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT11), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n272), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT64), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(new_n271), .B2(G137), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(KEYINPUT11), .ZN(new_n279));
  OAI21_X1  g093(.A(G131), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n273), .A2(G134), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n282), .B1(new_n278), .B2(KEYINPUT11), .ZN(new_n283));
  INV_X1    g097(.A(G131), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n274), .A2(new_n275), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n280), .A2(new_n281), .A3(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(KEYINPUT65), .B(G131), .C1(new_n276), .C2(new_n279), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n265), .A2(new_n270), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n237), .A2(new_n289), .A3(new_n264), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n193), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n262), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n243), .A2(new_n226), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n289), .B1(new_n257), .B2(new_n296), .ZN(new_n297));
  OR2_X1    g111(.A1(KEYINPUT86), .A2(KEYINPUT12), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT86), .B(KEYINPUT12), .Z(new_n300));
  OAI21_X1  g114(.A(new_n299), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n292), .A2(new_n193), .A3(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n187), .B(new_n188), .C1(new_n293), .C2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n187), .A2(new_n188), .ZN(new_n304));
  INV_X1    g118(.A(new_n193), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n268), .A2(new_n269), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n306), .B2(new_n289), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n292), .A2(new_n301), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n291), .A2(new_n307), .B1(new_n308), .B2(new_n305), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n304), .B1(new_n309), .B2(G469), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n303), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT9), .B(G234), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT78), .ZN(new_n313));
  OAI21_X1  g127(.A(G221), .B1(new_n313), .B2(G902), .ZN(new_n314));
  XNOR2_X1  g128(.A(G113), .B(G122), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(new_n206), .ZN(new_n316));
  XNOR2_X1  g130(.A(G125), .B(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n194), .ZN(new_n318));
  INV_X1    g132(.A(G125), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT75), .B1(new_n319), .B2(KEYINPUT74), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G125), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n321), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(KEYINPUT94), .B(new_n318), .C1(new_n327), .C2(new_n194), .ZN(new_n328));
  INV_X1    g142(.A(G237), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT68), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT68), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G237), .ZN(new_n332));
  AOI21_X1  g146(.A(G953), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT93), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G143), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n196), .A2(KEYINPUT93), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n333), .A2(G214), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n335), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n339), .B1(new_n333), .B2(G214), .ZN(new_n340));
  OAI211_X1 g154(.A(KEYINPUT18), .B(G131), .C1(new_n338), .C2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT94), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n342), .B(G146), .C1(new_n323), .C2(new_n326), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n330), .A2(new_n332), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(G214), .A3(new_n189), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n335), .ZN(new_n346));
  NAND2_X1  g160(.A1(KEYINPUT18), .A2(G131), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n333), .A2(G214), .A3(new_n337), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n328), .A2(new_n341), .A3(new_n343), .A4(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(G131), .B1(new_n338), .B2(new_n340), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT17), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n346), .A2(new_n284), .A3(new_n348), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT16), .B1(new_n323), .B2(new_n326), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT16), .B1(new_n321), .B2(G125), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n194), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT16), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n320), .A2(new_n325), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G140), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n359), .B1(new_n361), .B2(new_n322), .ZN(new_n362));
  OAI21_X1  g176(.A(G146), .B1(new_n362), .B2(new_n356), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n354), .A2(new_n358), .A3(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(KEYINPUT17), .B(G131), .C1(new_n338), .C2(new_n340), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT95), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n284), .B1(new_n346), .B2(new_n348), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(KEYINPUT95), .A3(KEYINPUT17), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n316), .B(new_n350), .C1(new_n364), .C2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT19), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n317), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n194), .B(new_n373), .C1(new_n327), .C2(new_n372), .ZN(new_n374));
  INV_X1    g188(.A(new_n353), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n363), .B(new_n374), .C1(new_n375), .C2(new_n368), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n350), .ZN(new_n377));
  INV_X1    g191(.A(new_n316), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n371), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT20), .ZN(new_n381));
  NOR2_X1   g195(.A1(G475), .A2(G902), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT96), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT96), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n380), .A2(new_n385), .A3(new_n381), .A4(new_n382), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n380), .A2(new_n382), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT20), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n384), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n196), .A2(G128), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n260), .A2(G143), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n392), .B(new_n271), .ZN(new_n393));
  XNOR2_X1  g207(.A(G116), .B(G122), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n208), .ZN(new_n395));
  INV_X1    g209(.A(G116), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT14), .A3(G122), .ZN(new_n397));
  INV_X1    g211(.A(new_n394), .ZN(new_n398));
  OAI211_X1 g212(.A(G107), .B(new_n397), .C1(new_n398), .C2(KEYINPUT14), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n393), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n394), .B(new_n208), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n392), .A2(new_n271), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT13), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n390), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n196), .A2(KEYINPUT13), .A3(G128), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n404), .A2(new_n405), .A3(new_n391), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n401), .B(new_n402), .C1(new_n271), .C2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G217), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n313), .A2(new_n408), .A3(G953), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n400), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n409), .B1(new_n400), .B2(new_n407), .ZN(new_n411));
  OAI211_X1 g225(.A(KEYINPUT97), .B(new_n188), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G478), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(KEYINPUT15), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n400), .A2(new_n407), .ZN(new_n416));
  INV_X1    g230(.A(new_n409), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n400), .A2(new_n409), .A3(new_n407), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n414), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n420), .A2(KEYINPUT97), .A3(new_n188), .A4(new_n421), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n415), .A2(new_n422), .A3(KEYINPUT98), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT98), .B1(new_n415), .B2(new_n422), .ZN(new_n424));
  NAND2_X1  g238(.A1(G234), .A2(G237), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n425), .A2(G952), .A3(new_n189), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(G898), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT99), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n425), .A2(G902), .A3(G953), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n426), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n423), .A2(new_n424), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n371), .ZN(new_n433));
  INV_X1    g247(.A(new_n358), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n194), .B1(new_n355), .B2(new_n357), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n436), .A2(new_n354), .A3(new_n367), .A4(new_n369), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n316), .B1(new_n437), .B2(new_n350), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n188), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G475), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n389), .A2(new_n432), .A3(new_n440), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n311), .A2(new_n314), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G214), .B1(G237), .B2(G902), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n445));
  INV_X1    g259(.A(G119), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G116), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n396), .A2(G119), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT2), .B(G113), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n449), .B(new_n450), .Z(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n220), .B2(KEYINPUT4), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n231), .B2(new_n236), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT5), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G113), .B1(new_n447), .B2(KEYINPUT5), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n449), .A2(new_n450), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n244), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n455), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G110), .B(G122), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n445), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n462), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n267), .A2(new_n235), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n467), .B1(new_n468), .B2(new_n454), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT88), .B1(new_n469), .B2(new_n464), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n453), .B1(new_n267), .B2(new_n235), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n472));
  NOR4_X1   g286(.A1(new_n471), .A2(new_n472), .A3(new_n467), .A4(new_n465), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n466), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n463), .A2(new_n445), .A3(new_n465), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n204), .A2(G125), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n262), .B2(G125), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n189), .A2(G224), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n477), .B(new_n478), .Z(new_n479));
  NAND3_X1  g293(.A1(new_n474), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n455), .A2(new_n462), .A3(new_n464), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n472), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n469), .A2(KEYINPUT88), .A3(new_n464), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n478), .A2(KEYINPUT7), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n477), .B(new_n485), .ZN(new_n486));
  XOR2_X1   g300(.A(new_n464), .B(KEYINPUT8), .Z(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n295), .B2(new_n461), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT89), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n458), .B1(new_n456), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n457), .A2(KEYINPUT89), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n460), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n488), .B1(new_n295), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT90), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n494), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n486), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(G902), .B1(new_n484), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n480), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G210), .B1(G237), .B2(G902), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n500), .B(KEYINPUT91), .Z(new_n501));
  XOR2_X1   g315(.A(new_n501), .B(KEYINPUT92), .Z(new_n502));
  NAND2_X1  g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n501), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n480), .A2(new_n498), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n444), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n408), .B1(G234), .B2(new_n188), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT22), .B(G137), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  XOR2_X1   g326(.A(G119), .B(G128), .Z(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT24), .B(G110), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(KEYINPUT73), .B1(new_n446), .B2(G128), .ZN(new_n516));
  OR2_X1    g330(.A1(new_n516), .A2(KEYINPUT23), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n516), .A2(KEYINPUT23), .B1(new_n446), .B2(G128), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n515), .B1(new_n519), .B2(G110), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(new_n358), .B2(new_n363), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n513), .A2(new_n514), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n519), .B2(G110), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n318), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(new_n435), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n512), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n520), .B1(new_n434), .B2(new_n435), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n363), .A2(new_n524), .A3(new_n318), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n511), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n188), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT76), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT25), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n527), .A2(new_n530), .A3(new_n188), .A4(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n508), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n527), .A2(new_n530), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n508), .A2(new_n188), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(KEYINPUT77), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n333), .A2(G210), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT26), .B(G101), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n287), .A2(new_n205), .A3(new_n288), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n271), .A2(G137), .ZN(new_n551));
  OAI21_X1  g365(.A(G131), .B1(new_n551), .B2(new_n282), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n262), .A2(new_n286), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n451), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT71), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n550), .A2(new_n451), .A3(new_n553), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT71), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n555), .B(new_n556), .C1(new_n559), .C2(new_n554), .ZN(new_n560));
  INV_X1    g374(.A(new_n557), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n561), .A2(KEYINPUT28), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n549), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT31), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n550), .A2(KEYINPUT30), .A3(new_n553), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n452), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n550), .A2(new_n553), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT30), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT67), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n567), .A2(KEYINPUT67), .A3(new_n568), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n566), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n561), .A2(new_n548), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n564), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n565), .A2(new_n452), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT67), .B1(new_n567), .B2(new_n568), .ZN(new_n578));
  AOI211_X1 g392(.A(new_n570), .B(KEYINPUT30), .C1(new_n550), .C2(new_n553), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(KEYINPUT31), .A3(new_n574), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n563), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(G472), .A2(G902), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT32), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n560), .A2(new_n562), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n548), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n580), .A2(KEYINPUT31), .A3(new_n574), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT31), .B1(new_n580), .B2(new_n574), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT32), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n583), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n586), .A2(new_n548), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n549), .B1(new_n580), .B2(new_n557), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n594), .A2(KEYINPUT29), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n554), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT72), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(new_n598), .A3(new_n557), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n567), .A2(KEYINPUT72), .A3(new_n452), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(KEYINPUT28), .A3(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n601), .A2(KEYINPUT29), .A3(new_n562), .A4(new_n549), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n188), .ZN(new_n603));
  OAI21_X1  g417(.A(G472), .B1(new_n596), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n543), .B1(new_n593), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n442), .A2(new_n506), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  INV_X1    g421(.A(G472), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n590), .B2(new_n188), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n582), .A2(new_n584), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n609), .A2(new_n610), .A3(new_n543), .ZN(new_n611));
  INV_X1    g425(.A(new_n314), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n303), .B2(new_n310), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n420), .A2(KEYINPUT33), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n418), .A2(new_n616), .A3(new_n419), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(G478), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n420), .A2(new_n413), .A3(new_n188), .ZN(new_n620));
  NAND2_X1  g434(.A1(G478), .A2(G902), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AOI211_X1 g436(.A(new_n431), .B(new_n622), .C1(new_n389), .C2(new_n440), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n480), .A2(new_n498), .A3(new_n504), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n504), .B1(new_n480), .B2(new_n498), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n623), .B(new_n443), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n499), .A2(new_n501), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n444), .B1(new_n629), .B2(new_n505), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT100), .B1(new_n630), .B2(new_n623), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n614), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT102), .B(G104), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT101), .B(KEYINPUT34), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  INV_X1    g450(.A(new_n383), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n381), .B1(new_n380), .B2(new_n382), .ZN(new_n638));
  OAI221_X1 g452(.A(new_n440), .B1(new_n423), .B2(new_n424), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n431), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n614), .A2(new_n630), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n528), .A2(new_n529), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n512), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT103), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n645), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n541), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n538), .A2(new_n644), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n649), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT104), .B1(new_n537), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n653), .A2(new_n610), .A3(new_n609), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n442), .A2(new_n506), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  AOI21_X1  g471(.A(new_n653), .B1(new_n593), .B2(new_n604), .ZN(new_n658));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n430), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n426), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n639), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n630), .A2(new_n658), .A3(new_n613), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  XNOR2_X1  g480(.A(new_n662), .B(KEYINPUT39), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n613), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT40), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n599), .A2(new_n548), .A3(new_n600), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n670), .A2(KEYINPUT105), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(KEYINPUT105), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n580), .A2(new_n574), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n675), .B2(G902), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT106), .B1(new_n593), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n593), .A2(KEYINPUT106), .A3(new_n676), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n502), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n480), .B2(new_n498), .ZN(new_n682));
  OAI21_X1  g496(.A(KEYINPUT38), .B1(new_n624), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT38), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n503), .A2(new_n684), .A3(new_n505), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n389), .A2(new_n440), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n423), .A2(new_n424), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n444), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n538), .A2(new_n649), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n669), .A2(new_n680), .A3(new_n686), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G143), .ZN(G45));
  INV_X1    g508(.A(new_n622), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n687), .A2(new_n695), .A3(new_n662), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n630), .A2(new_n658), .A3(new_n613), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  NAND2_X1  g513(.A1(new_n291), .A2(new_n292), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n302), .B1(new_n700), .B2(new_n305), .ZN(new_n701));
  OAI21_X1  g515(.A(G469), .B1(new_n701), .B2(G902), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n702), .A2(new_n314), .A3(new_n303), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n605), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n626), .A2(new_n627), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n630), .A2(KEYINPUT100), .A3(new_n623), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT41), .B(G113), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND4_X1  g523(.A1(new_n630), .A2(new_n605), .A3(new_n703), .A4(new_n640), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  NAND4_X1  g525(.A1(new_n630), .A2(new_n658), .A3(new_n703), .A4(new_n441), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  AOI21_X1  g527(.A(new_n690), .B1(new_n629), .B2(new_n505), .ZN(new_n714));
  OAI21_X1  g528(.A(G472), .B1(new_n582), .B2(G902), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n537), .B1(new_n541), .B2(new_n539), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n588), .A2(new_n589), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n549), .B1(new_n601), .B2(new_n562), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n583), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n715), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n431), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n714), .A2(new_n721), .A3(new_n703), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n714), .A2(new_n721), .A3(new_n703), .A4(KEYINPUT107), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  NAND3_X1  g541(.A1(new_n715), .A2(new_n719), .A3(new_n691), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n696), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n630), .A2(new_n729), .A3(new_n703), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  NOR3_X1   g545(.A1(new_n624), .A2(new_n682), .A3(new_n444), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n304), .B(KEYINPUT108), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n309), .B2(G469), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n612), .B1(new_n303), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n732), .A2(new_n605), .A3(new_n697), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n497), .B1(new_n470), .B2(new_n473), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n188), .ZN(new_n741));
  INV_X1    g555(.A(new_n475), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n742), .B1(new_n484), .B2(new_n466), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n741), .B1(new_n743), .B2(new_n479), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n443), .B(new_n505), .C1(new_n744), .C2(new_n681), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n303), .A2(new_n735), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n314), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n738), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n605), .A3(new_n697), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n739), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  NAND4_X1  g566(.A1(new_n732), .A2(new_n605), .A3(new_n664), .A4(new_n736), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G134), .ZN(G36));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n687), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n389), .A2(KEYINPUT111), .A3(new_n440), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(KEYINPUT43), .A3(new_n695), .A4(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n687), .B2(new_n622), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n691), .B1(new_n609), .B2(new_n610), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n762), .A2(KEYINPUT112), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(KEYINPUT112), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n309), .A2(KEYINPUT45), .ZN(new_n768));
  OAI21_X1  g582(.A(G469), .B1(new_n309), .B2(KEYINPUT45), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n733), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT46), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(KEYINPUT46), .B(new_n733), .C1(new_n768), .C2(new_n769), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n303), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n314), .ZN(new_n775));
  INV_X1    g589(.A(new_n667), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT110), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n774), .A2(new_n778), .A3(new_n314), .A4(new_n667), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n745), .B1(new_n765), .B2(new_n766), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n767), .A2(new_n777), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  NAND2_X1  g596(.A1(new_n775), .A2(KEYINPUT47), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT47), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n774), .A2(new_n784), .A3(new_n314), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n697), .A2(new_n593), .A3(new_n604), .A4(new_n543), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n745), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n783), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  NAND3_X1  g603(.A1(new_n702), .A2(new_n314), .A3(new_n303), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n745), .A2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n791), .A2(new_n426), .A3(new_n761), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n605), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT48), .ZN(new_n794));
  INV_X1    g608(.A(G952), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n661), .B(new_n720), .C1(new_n758), .C2(new_n760), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n630), .A2(new_n703), .ZN(new_n797));
  AOI211_X1 g611(.A(new_n795), .B(G953), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n679), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n677), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n687), .A2(new_n695), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n543), .A2(new_n661), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n800), .A2(new_n802), .A3(new_n791), .A4(new_n803), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n798), .A2(KEYINPUT119), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT119), .B1(new_n798), .B2(new_n804), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n794), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n703), .A2(new_n444), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n808), .B1(new_n686), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n790), .A2(new_n443), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(KEYINPUT116), .A3(new_n683), .A4(new_n685), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n796), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n810), .A2(KEYINPUT50), .A3(new_n796), .A4(new_n812), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n728), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n792), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n687), .A2(new_n695), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n800), .A2(new_n791), .A3(new_n803), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n817), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n702), .A2(KEYINPUT115), .A3(new_n303), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT115), .B1(new_n702), .B2(new_n303), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n314), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n783), .A2(new_n785), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n796), .A2(new_n732), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT51), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT118), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n828), .A2(new_n829), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n822), .B1(new_n815), .B2(new_n816), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(KEYINPUT51), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n807), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n824), .A2(KEYINPUT117), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n832), .B1(new_n833), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n837), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n836), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n665), .A2(new_n730), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n691), .A2(new_n663), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n714), .A2(new_n736), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n680), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n843), .A2(new_n846), .A3(new_n847), .A4(new_n698), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n665), .A2(new_n698), .A3(new_n730), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n714), .A2(new_n736), .A3(new_n844), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n800), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT52), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n415), .A2(new_n422), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n389), .A2(new_n440), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n431), .B1(new_n801), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n506), .A2(new_n613), .A3(new_n856), .A4(new_n611), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n857), .A2(new_n606), .A3(new_n655), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n732), .A2(new_n729), .A3(new_n736), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n854), .A2(new_n663), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n440), .B(new_n860), .C1(new_n637), .C2(new_n638), .ZN(new_n861));
  AOI211_X1 g675(.A(new_n612), .B(new_n861), .C1(new_n303), .C2(new_n310), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n732), .A2(new_n658), .A3(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n753), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n751), .A2(new_n858), .A3(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n710), .A2(new_n712), .ZN(new_n866));
  INV_X1    g680(.A(new_n704), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n628), .B2(new_n631), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n726), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT53), .B1(new_n853), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n753), .A2(new_n863), .A3(new_n859), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n750), .B2(new_n739), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n710), .A2(new_n712), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n707), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n873), .A2(new_n726), .A3(new_n875), .A4(new_n858), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n848), .A2(new_n852), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n665), .A2(new_n730), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT53), .B1(new_n878), .B2(KEYINPUT52), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT54), .B1(new_n871), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n878), .A2(KEYINPUT52), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT53), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n865), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n869), .A2(KEYINPUT114), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT114), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n875), .A2(new_n886), .A3(new_n726), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n853), .A2(new_n884), .A3(new_n885), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n876), .B2(new_n877), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT54), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n881), .A2(new_n892), .ZN(new_n893));
  OAI22_X1  g707(.A1(new_n842), .A2(new_n893), .B1(G952), .B2(G953), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n702), .A2(new_n303), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT49), .ZN(new_n896));
  NOR4_X1   g710(.A1(new_n543), .A2(new_n444), .A3(new_n622), .A4(new_n612), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n896), .A2(new_n756), .A3(new_n757), .A4(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n895), .A2(KEYINPUT49), .ZN(new_n899));
  NOR4_X1   g713(.A1(new_n680), .A2(new_n898), .A3(new_n686), .A4(new_n899), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT113), .Z(new_n901));
  NAND2_X1  g715(.A1(new_n894), .A2(new_n901), .ZN(G75));
  NOR2_X1   g716(.A1(new_n189), .A2(G952), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT120), .Z(new_n904));
  AOI21_X1  g718(.A(new_n188), .B1(new_n888), .B2(new_n890), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n905), .A2(new_n502), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n743), .B(new_n479), .Z(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n904), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n905), .A2(new_n501), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n908), .B1(new_n912), .B2(new_n909), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n911), .A2(new_n913), .ZN(G51));
  XOR2_X1   g728(.A(new_n733), .B(KEYINPUT57), .Z(new_n915));
  AND3_X1   g729(.A1(new_n888), .A2(new_n891), .A3(new_n890), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n891), .B1(new_n888), .B2(new_n890), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n701), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n768), .A2(new_n769), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n905), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n903), .B1(new_n920), .B2(new_n922), .ZN(G54));
  NAND2_X1  g737(.A1(KEYINPUT58), .A2(G475), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n905), .A2(new_n380), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n380), .B1(new_n905), .B2(new_n925), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n903), .ZN(G60));
  INV_X1    g742(.A(new_n618), .ZN(new_n929));
  XNOR2_X1  g743(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n621), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n929), .B(new_n931), .C1(new_n916), .C2(new_n917), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n904), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n929), .B1(new_n893), .B2(new_n931), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n933), .A2(new_n934), .ZN(G63));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n936));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT60), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n888), .B2(new_n890), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n648), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n904), .B1(new_n939), .B2(new_n539), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n539), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n888), .A2(new_n890), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n944), .B1(new_n945), .B2(new_n938), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n946), .A2(KEYINPUT61), .A3(new_n904), .A4(new_n940), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n943), .A2(new_n947), .ZN(G66));
  AOI21_X1  g762(.A(new_n189), .B1(new_n428), .B2(G224), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT122), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n875), .A2(new_n726), .A3(new_n858), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n950), .B1(new_n951), .B2(G953), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT123), .ZN(new_n953));
  INV_X1    g767(.A(G898), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n743), .B1(new_n954), .B2(G953), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n953), .B(new_n955), .ZN(G69));
  OAI21_X1  g770(.A(new_n565), .B1(new_n578), .B2(new_n579), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n373), .B1(new_n327), .B2(new_n372), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n957), .B(new_n958), .Z(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(G900), .B2(G953), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n777), .A2(new_n605), .A3(new_n714), .A4(new_n779), .ZN(new_n961));
  AND4_X1   g775(.A1(new_n751), .A2(new_n961), .A3(new_n753), .A4(new_n788), .ZN(new_n962));
  INV_X1    g776(.A(new_n849), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n781), .A2(KEYINPUT125), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT125), .B1(new_n781), .B2(new_n963), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n960), .B1(new_n966), .B2(G953), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n693), .A2(KEYINPUT62), .A3(new_n963), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT62), .B1(new_n693), .B2(new_n963), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n801), .A2(new_n855), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n668), .A2(new_n605), .A3(new_n732), .A4(new_n972), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT124), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n974), .A2(new_n788), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n781), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n189), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n959), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT126), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n967), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n980), .B1(new_n967), .B2(new_n978), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n981), .A2(new_n982), .ZN(G72));
  OAI21_X1  g797(.A(new_n549), .B1(new_n573), .B2(new_n561), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n975), .A2(new_n781), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n985), .B(new_n951), .C1(new_n970), .C2(new_n969), .ZN(new_n986));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  AOI21_X1  g802(.A(new_n984), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n580), .A2(new_n557), .A3(new_n548), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n962), .B(new_n951), .C1(new_n964), .C2(new_n965), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n990), .B1(new_n991), .B2(new_n988), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n871), .A2(new_n880), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n988), .B1(new_n674), .B2(new_n595), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR4_X1   g809(.A1(new_n989), .A2(new_n992), .A3(new_n995), .A4(new_n903), .ZN(G57));
endmodule


