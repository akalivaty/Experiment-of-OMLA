//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(G134gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G127gat), .ZN(new_n204));
  INV_X1    g003(.A(G127gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G134gat), .ZN(new_n206));
  NOR3_X1   g005(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT1), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT73), .ZN(new_n209));
  INV_X1    g008(.A(G113gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(G120gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(G120gat), .ZN(new_n212));
  INV_X1    g011(.A(G120gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT73), .A3(G113gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n211), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT74), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n211), .A2(new_n214), .A3(KEYINPUT74), .A4(new_n212), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n208), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(G113gat), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT1), .B1(new_n220), .B2(new_n212), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  OR2_X1    g021(.A1(KEYINPUT70), .A2(KEYINPUT71), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT70), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(new_n203), .A3(G127gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(KEYINPUT70), .A2(KEYINPUT71), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n205), .A2(G134gat), .ZN(new_n227));
  AND4_X1   g026(.A1(new_n223), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n225), .A2(new_n227), .B1(new_n223), .B2(new_n226), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n222), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT72), .ZN(new_n231));
  NOR3_X1   g030(.A1(new_n205), .A2(KEYINPUT70), .A3(G134gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(KEYINPUT70), .A2(KEYINPUT71), .ZN(new_n233));
  INV_X1    g032(.A(new_n226), .ZN(new_n234));
  OAI22_X1  g033(.A1(new_n232), .A2(new_n204), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n225), .A2(new_n223), .A3(new_n226), .A4(new_n227), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT72), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n238), .A3(new_n222), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n219), .B1(new_n231), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G169gat), .ZN(new_n248));
  INV_X1    g047(.A(G176gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n250), .A2(KEYINPUT26), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n243), .A2(new_n247), .A3(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT27), .B(G183gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT28), .ZN(new_n254));
  INV_X1    g053(.A(G190gat), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n253), .A2(KEYINPUT68), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G183gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT27), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT27), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G183gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n260), .A3(new_n255), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n254), .A2(KEYINPUT68), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n261), .A2(new_n262), .B1(G183gat), .B2(G190gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n252), .A2(new_n256), .A3(new_n263), .ZN(new_n264));
  AND3_X1   g063(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266));
  OAI22_X1  g065(.A1(new_n265), .A2(new_n244), .B1(KEYINPUT23), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NOR3_X1   g068(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT24), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT24), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(G183gat), .A3(G190gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n267), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT23), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT65), .B1(new_n250), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n266), .A2(new_n280), .A3(KEYINPUT23), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT25), .B1(new_n277), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n250), .A2(new_n278), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT25), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n285), .B1(new_n266), .B2(KEYINPUT23), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n247), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n276), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT67), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n276), .A2(KEYINPUT67), .A3(new_n289), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n287), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n264), .B1(new_n283), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n240), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n270), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n276), .A2(new_n297), .A3(new_n268), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n245), .A2(new_n246), .B1(new_n278), .B2(new_n250), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n282), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(new_n285), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT67), .B1(new_n276), .B2(new_n289), .ZN(new_n302));
  AOI211_X1 g101(.A(new_n291), .B(new_n288), .C1(new_n273), .C2(new_n275), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n299), .B(new_n286), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n263), .A2(new_n256), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n301), .A2(new_n304), .B1(new_n305), .B2(new_n252), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n217), .A2(new_n218), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n207), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n238), .B1(new_n237), .B2(new_n222), .ZN(new_n309));
  AOI211_X1 g108(.A(KEYINPUT72), .B(new_n221), .C1(new_n235), .C2(new_n236), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n296), .A2(new_n312), .A3(G227gat), .A4(G233gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT32), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT33), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(G15gat), .B(G43gat), .Z(new_n317));
  XNOR2_X1  g116(.A(G71gat), .B(G99gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n314), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n319), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n313), .B(KEYINPUT32), .C1(new_n315), .C2(new_n321), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n320), .A2(KEYINPUT77), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT77), .B1(new_n320), .B2(new_n322), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n296), .A2(new_n312), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G227gat), .A2(G233gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n296), .A2(new_n312), .A3(KEYINPUT75), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT34), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT34), .B1(G227gat), .B2(G233gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n325), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n325), .A2(KEYINPUT76), .A3(new_n332), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n323), .A2(new_n324), .A3(new_n338), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n330), .A2(KEYINPUT34), .B1(new_n335), .B2(new_n336), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n320), .A2(new_n322), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n202), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n324), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT77), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n340), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n323), .B1(new_n324), .B2(new_n338), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT36), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT84), .ZN(new_n352));
  XNOR2_X1  g151(.A(G78gat), .B(G106gat), .ZN(new_n353));
  INV_X1    g152(.A(G50gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n352), .B(new_n355), .Z(new_n356));
  INV_X1    g155(.A(G228gat), .ZN(new_n357));
  INV_X1    g156(.A(G233gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  OR2_X1    g159(.A1(KEYINPUT80), .A2(G141gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(KEYINPUT80), .A2(G141gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(G148gat), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G148gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G141gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT2), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G141gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G148gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n368), .ZN(new_n375));
  INV_X1    g174(.A(new_n367), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n376), .A2(new_n370), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n366), .A2(new_n371), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT79), .B(KEYINPUT29), .ZN(new_n379));
  AND2_X1   g178(.A1(G211gat), .A2(G218gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(G211gat), .A2(G218gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G204gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT78), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(G197gat), .ZN(new_n386));
  INV_X1    g185(.A(G197gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n387), .A2(KEYINPUT78), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n384), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(KEYINPUT78), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n385), .A2(G197gat), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n391), .A3(G204gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n380), .A2(KEYINPUT22), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n383), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  AOI211_X1 g195(.A(new_n382), .B(new_n394), .C1(new_n389), .C2(new_n392), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n379), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n378), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n379), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n378), .B2(new_n399), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n390), .A2(new_n391), .A3(G204gat), .ZN(new_n403));
  AOI21_X1  g202(.A(G204gat), .B1(new_n390), .B2(new_n391), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n395), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n382), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n393), .A2(new_n383), .A3(new_n395), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n360), .B1(new_n400), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n396), .B2(new_n397), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n378), .B1(new_n412), .B2(new_n399), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n359), .B1(new_n402), .B2(new_n408), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT85), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n378), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT29), .B1(new_n406), .B2(new_n407), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(KEYINPUT3), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n396), .A2(new_n397), .ZN(new_n420));
  XNOR2_X1  g219(.A(G141gat), .B(G148gat), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n370), .B(new_n376), .C1(new_n421), .C2(KEYINPUT2), .ZN(new_n422));
  INV_X1    g221(.A(new_n365), .ZN(new_n423));
  INV_X1    g222(.A(new_n362), .ZN(new_n424));
  NOR2_X1   g223(.A1(KEYINPUT80), .A2(G141gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n423), .B1(new_n426), .B2(G148gat), .ZN(new_n427));
  INV_X1    g226(.A(new_n371), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n422), .B(new_n399), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n379), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n360), .B1(new_n420), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT85), .B1(new_n419), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n410), .B1(new_n416), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(G22gat), .ZN(new_n434));
  INV_X1    g233(.A(G22gat), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n435), .B(new_n410), .C1(new_n416), .C2(new_n432), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n356), .B1(new_n437), .B2(KEYINPUT86), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT87), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n439), .B1(new_n437), .B2(KEYINPUT86), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT86), .ZN(new_n441));
  AOI211_X1 g240(.A(new_n441), .B(KEYINPUT87), .C1(new_n434), .C2(new_n436), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n438), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n356), .ZN(new_n444));
  INV_X1    g243(.A(new_n436), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n415), .B1(new_n413), .B2(new_n414), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n419), .A2(new_n431), .A3(KEYINPUT85), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n435), .B1(new_n448), .B2(new_n410), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n444), .B1(new_n450), .B2(new_n441), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT86), .B1(new_n445), .B2(new_n449), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT87), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n437), .A2(KEYINPUT86), .A3(new_n439), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n443), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(G225gat), .A2(G233gat), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n376), .A2(new_n370), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n460), .B1(new_n374), .B2(new_n368), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n363), .A2(new_n365), .B1(new_n370), .B2(new_n369), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT3), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n463), .A2(new_n429), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n459), .B1(new_n311), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT4), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n466), .B1(new_n240), .B2(new_n378), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n308), .B(new_n378), .C1(new_n309), .C2(new_n310), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n468), .A2(KEYINPUT4), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n465), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT81), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT5), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n311), .A2(new_n417), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(new_n468), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n473), .B1(new_n475), .B2(new_n459), .ZN(new_n476));
  OAI211_X1 g275(.A(KEYINPUT81), .B(new_n465), .C1(new_n467), .C2(new_n469), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n472), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n240), .A2(KEYINPUT82), .A3(new_n466), .A4(new_n378), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n311), .A2(new_n464), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n468), .A2(KEYINPUT4), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n231), .A2(new_n239), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n483), .A2(new_n466), .A3(new_n308), .A4(new_n378), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT82), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n481), .A2(new_n473), .A3(new_n486), .A4(new_n458), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n478), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G1gat), .B(G29gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT0), .ZN(new_n490));
  XNOR2_X1  g289(.A(G57gat), .B(G85gat), .ZN(new_n491));
  XOR2_X1   g290(.A(new_n490), .B(new_n491), .Z(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n492), .A3(new_n487), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n492), .B1(new_n478), .B2(new_n487), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G8gat), .B(G36gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(G64gat), .B(G92gat), .ZN(new_n502));
  XOR2_X1   g301(.A(new_n501), .B(new_n502), .Z(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G226gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(new_n358), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(new_n306), .B2(KEYINPUT29), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n295), .A2(new_n506), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n508), .A2(new_n408), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n507), .B1(new_n306), .B2(new_n401), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n408), .B1(new_n511), .B2(new_n509), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n504), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n506), .B1(new_n295), .B2(new_n379), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n306), .A2(new_n507), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n420), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n508), .A2(new_n408), .A3(new_n509), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n503), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n513), .A2(KEYINPUT30), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT30), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n516), .A2(new_n517), .A3(new_n520), .A4(new_n503), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n500), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n350), .B1(new_n457), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n458), .B1(new_n481), .B2(new_n486), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT39), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n493), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n482), .A2(new_n484), .A3(new_n485), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n479), .A2(new_n480), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n459), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT88), .B1(new_n475), .B2(new_n459), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT88), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n474), .A2(new_n533), .A3(new_n468), .A4(new_n458), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n534), .A2(KEYINPUT39), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT40), .B1(new_n528), .B2(new_n536), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n537), .A2(new_n522), .A3(new_n498), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n528), .A2(KEYINPUT40), .A3(new_n536), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n455), .A2(new_n443), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT89), .B(KEYINPUT38), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT90), .B(KEYINPUT37), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n516), .A2(new_n517), .A3(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n543), .A2(new_n504), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT37), .B1(new_n510), .B2(new_n512), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n408), .B1(new_n514), .B2(new_n515), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n508), .A2(new_n420), .A3(new_n509), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT37), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n549), .A2(new_n543), .A3(new_n504), .A4(new_n541), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n518), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT91), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n498), .A2(new_n553), .A3(KEYINPUT6), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n498), .B2(KEYINPUT6), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n497), .B(new_n552), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n525), .B1(new_n540), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n537), .ZN(new_n558));
  INV_X1    g357(.A(new_n522), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n558), .A2(new_n494), .A3(new_n559), .A4(new_n539), .ZN(new_n560));
  AND4_X1   g359(.A1(new_n525), .A2(new_n556), .A3(new_n456), .A4(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n524), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n347), .A2(new_n348), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n456), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT35), .B1(new_n564), .B2(new_n523), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n497), .B1(new_n554), .B2(new_n555), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n559), .A2(KEYINPUT35), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n456), .A2(new_n566), .A3(new_n563), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G229gat), .A2(G233gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n571), .B(KEYINPUT13), .Z(new_n572));
  XNOR2_X1  g371(.A(G43gat), .B(G50gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT15), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G29gat), .A2(G36gat), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NOR3_X1   g377(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n573), .A2(KEYINPUT15), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n576), .A3(new_n574), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n579), .A2(KEYINPUT94), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(KEYINPUT94), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n578), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n581), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G8gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(G15gat), .B(G22gat), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n589), .A2(G1gat), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT16), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n589), .B1(new_n591), .B2(G1gat), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n588), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n590), .A2(new_n588), .A3(new_n592), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT96), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n595), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT96), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n597), .A2(new_n598), .A3(new_n593), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n587), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n596), .A2(new_n599), .A3(new_n587), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n572), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n587), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT17), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n597), .A2(new_n593), .ZN(new_n606));
  XOR2_X1   g405(.A(KEYINPUT95), .B(KEYINPUT17), .Z(new_n607));
  OAI211_X1 g406(.A(new_n605), .B(new_n606), .C1(new_n604), .C2(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n608), .A2(KEYINPUT18), .A3(new_n600), .A4(new_n571), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n600), .A3(new_n571), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G113gat), .B(G141gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(G197gat), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT11), .B(G169gat), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT93), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n610), .B(new_n613), .C1(KEYINPUT98), .C2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n603), .A2(new_n609), .A3(KEYINPUT98), .ZN(new_n622));
  INV_X1    g421(.A(new_n613), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n603), .A2(new_n609), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n622), .B(new_n619), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n621), .A2(new_n625), .A3(KEYINPUT99), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G99gat), .A2(G106gat), .ZN(new_n631));
  INV_X1    g430(.A(G85gat), .ZN(new_n632));
  INV_X1    g431(.A(G92gat), .ZN(new_n633));
  AOI22_X1  g432(.A1(KEYINPUT8), .A2(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT7), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(new_n632), .B2(new_n633), .ZN(new_n636));
  NAND3_X1  g435(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G99gat), .B(G106gat), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n605), .B(new_n643), .C1(new_n604), .C2(new_n607), .ZN(new_n644));
  AND3_X1   g443(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n645));
  INV_X1    g444(.A(new_n643), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n645), .B1(new_n646), .B2(new_n587), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(G190gat), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n644), .A2(new_n647), .A3(new_n255), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(G218gat), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT101), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n649), .A2(G218gat), .A3(new_n650), .ZN(new_n654));
  XNOR2_X1  g453(.A(G134gat), .B(G162gat), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n657), .B1(new_n653), .B2(new_n654), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(G71gat), .A2(G78gat), .ZN(new_n662));
  OR2_X1    g461(.A1(G71gat), .A2(G78gat), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT9), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(G57gat), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT100), .B1(new_n666), .B2(G64gat), .ZN(new_n667));
  INV_X1    g466(.A(G64gat), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n667), .B1(G57gat), .B2(new_n668), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n666), .A2(KEYINPUT100), .A3(G64gat), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n666), .A2(G64gat), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n668), .A2(G57gat), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT9), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n662), .A3(new_n663), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT21), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(G231gat), .A2(G233gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(new_n205), .ZN(new_n681));
  INV_X1    g480(.A(new_n676), .ZN(new_n682));
  AOI211_X1 g481(.A(new_n599), .B(new_n596), .C1(KEYINPUT21), .C2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n685));
  INV_X1    g484(.A(G155gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(G183gat), .B(G211gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n684), .B(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n661), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(G120gat), .B(G148gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT103), .ZN(new_n694));
  XNOR2_X1  g493(.A(G176gat), .B(G204gat), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n694), .B(new_n695), .Z(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n641), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n643), .A2(new_n699), .A3(new_n682), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n641), .B(new_n642), .C1(new_n676), .C2(new_n698), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(G230gat), .A2(G233gat), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n697), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT10), .B1(new_n700), .B2(new_n701), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n646), .A2(KEYINPUT10), .A3(new_n682), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  OAI211_X1 g510(.A(KEYINPUT104), .B(new_n703), .C1(new_n706), .C2(new_n707), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n711), .A2(new_n712), .B1(new_n704), .B2(new_n702), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n709), .B1(new_n713), .B2(new_n696), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(KEYINPUT105), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n716), .B(new_n709), .C1(new_n713), .C2(new_n696), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n692), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n570), .A2(new_n630), .A3(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n500), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n559), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT16), .B(G8gat), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT106), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT42), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n729));
  OAI211_X1 g528(.A(KEYINPUT106), .B(new_n729), .C1(new_n725), .C2(new_n726), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n725), .A2(G8gat), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n728), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT107), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n728), .A2(new_n734), .A3(new_n730), .A4(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(G1325gat));
  INV_X1    g535(.A(new_n350), .ZN(new_n737));
  OAI21_X1  g536(.A(G15gat), .B1(new_n720), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(G15gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n563), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n720), .B2(new_n740), .ZN(G1326gat));
  INV_X1    g540(.A(new_n570), .ZN(new_n742));
  INV_X1    g541(.A(new_n630), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n457), .A3(new_n719), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT108), .ZN(new_n746));
  XNOR2_X1  g545(.A(KEYINPUT43), .B(G22gat), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1327gat));
  NOR2_X1   g547(.A1(new_n691), .A2(new_n718), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n626), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n660), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n658), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n562), .A2(KEYINPUT109), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n524), .B(new_n759), .C1(new_n557), .C2(new_n561), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n757), .B1(new_n761), .B2(new_n569), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n756), .B1(new_n570), .B2(new_n755), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n753), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G29gat), .B1(new_n767), .B2(new_n500), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n750), .A2(new_n661), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n744), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(G29gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n722), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n769), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  OR3_X1    g573(.A1(new_n771), .A2(new_n769), .A3(new_n773), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n768), .A2(new_n774), .A3(new_n775), .ZN(G1328gat));
  OAI21_X1  g575(.A(G36gat), .B1(new_n767), .B2(new_n522), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n522), .A2(G36gat), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT46), .B1(new_n771), .B2(new_n778), .ZN(new_n779));
  OR3_X1    g578(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n778), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(G1329gat));
  OAI211_X1 g580(.A(new_n350), .B(new_n752), .C1(new_n762), .C2(new_n764), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G43gat), .ZN(new_n783));
  INV_X1    g582(.A(new_n771), .ZN(new_n784));
  INV_X1    g583(.A(G43gat), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(new_n785), .A3(new_n563), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(G1330gat));
  NAND2_X1  g588(.A1(new_n766), .A2(new_n457), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G50gat), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n771), .A2(G50gat), .A3(new_n456), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(KEYINPUT48), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT48), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n354), .B1(new_n766), .B2(new_n457), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(new_n792), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n797), .ZN(G1331gat));
  NAND2_X1  g597(.A1(new_n761), .A2(new_n569), .ZN(new_n799));
  INV_X1    g598(.A(new_n718), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n692), .A2(new_n626), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(new_n500), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(new_n666), .ZN(G1332gat));
  NOR2_X1   g603(.A1(new_n802), .A2(new_n522), .ZN(new_n805));
  NOR2_X1   g604(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n806));
  AND2_X1   g605(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n805), .B2(new_n806), .ZN(G1333gat));
  OAI21_X1  g608(.A(G71gat), .B1(new_n802), .B2(new_n737), .ZN(new_n810));
  INV_X1    g609(.A(G71gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n563), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n802), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g612(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n814));
  XNOR2_X1  g613(.A(new_n813), .B(new_n814), .ZN(G1334gat));
  NOR2_X1   g614(.A1(new_n802), .A2(new_n456), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g616(.A1(new_n690), .A2(new_n751), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n800), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n819), .B1(new_n762), .B2(new_n764), .ZN(new_n820));
  OAI21_X1  g619(.A(G85gat), .B1(new_n820), .B2(new_n500), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n758), .A2(new_n760), .B1(new_n565), .B2(new_n568), .ZN(new_n822));
  INV_X1    g621(.A(new_n818), .ZN(new_n823));
  OR2_X1    g622(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n755), .A3(new_n824), .ZN(new_n825));
  OAI211_X1 g624(.A(KEYINPUT112), .B(KEYINPUT51), .C1(new_n822), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n827));
  INV_X1    g626(.A(new_n825), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n799), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n718), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n722), .A2(new_n632), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n821), .B1(new_n831), .B2(new_n832), .ZN(G1336gat));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n522), .A2(G92gat), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n826), .A2(new_n829), .A3(new_n718), .A4(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n834), .B1(new_n836), .B2(KEYINPUT113), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n559), .B(new_n819), .C1(new_n762), .C2(new_n764), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G92gat), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n836), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n837), .B(new_n840), .ZN(G1337gat));
  INV_X1    g640(.A(G99gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n563), .A2(new_n842), .A3(new_n718), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT114), .Z(new_n844));
  NAND2_X1  g643(.A1(new_n830), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(G99gat), .B1(new_n820), .B2(new_n737), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1338gat));
  OAI211_X1 g646(.A(new_n457), .B(new_n819), .C1(new_n762), .C2(new_n764), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G106gat), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n456), .A2(G106gat), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n826), .A2(new_n829), .A3(new_n718), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n849), .B(new_n853), .C1(new_n850), .C2(KEYINPUT53), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(G1339gat));
  NOR3_X1   g657(.A1(new_n601), .A2(new_n602), .A3(new_n572), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n571), .B1(new_n608), .B2(new_n600), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n617), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n610), .A2(new_n620), .A3(new_n613), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n865), .B1(new_n715), .B2(new_n717), .ZN(new_n866));
  XNOR2_X1  g665(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n711), .A2(new_n712), .A3(new_n867), .ZN(new_n868));
  OR3_X1    g667(.A1(new_n706), .A2(new_n707), .A3(new_n703), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n708), .A3(KEYINPUT54), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n868), .A2(new_n697), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n868), .A2(KEYINPUT55), .A3(new_n870), .A4(new_n697), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n709), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n751), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n661), .B1(new_n866), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n865), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n873), .A2(new_n709), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n755), .A2(new_n878), .A3(new_n874), .A4(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n691), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n692), .A2(new_n626), .A3(new_n718), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT118), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n882), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n879), .A2(new_n626), .A3(new_n874), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n878), .A2(new_n718), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n755), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n661), .A2(new_n865), .A3(new_n875), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n690), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n884), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n883), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n457), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n500), .A2(new_n559), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n563), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G113gat), .B1(new_n895), .B2(new_n743), .ZN(new_n896));
  NOR4_X1   g695(.A1(new_n892), .A2(new_n500), .A3(new_n559), .A4(new_n564), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n210), .A3(new_n626), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT119), .Z(G1340gat));
  NOR3_X1   g699(.A1(new_n895), .A2(new_n213), .A3(new_n800), .ZN(new_n901));
  AOI21_X1  g700(.A(G120gat), .B1(new_n897), .B2(new_n718), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(G1341gat));
  OAI21_X1  g702(.A(G127gat), .B1(new_n895), .B2(new_n690), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n897), .A2(new_n205), .A3(new_n691), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1342gat));
  NAND3_X1  g705(.A1(new_n897), .A2(new_n203), .A3(new_n755), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n907), .A2(KEYINPUT56), .ZN(new_n908));
  OAI21_X1  g707(.A(G134gat), .B1(new_n895), .B2(new_n661), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(KEYINPUT56), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(G1343gat));
  NAND2_X1  g710(.A1(new_n737), .A2(new_n457), .ZN(new_n912));
  NOR4_X1   g711(.A1(new_n892), .A2(new_n500), .A3(new_n559), .A4(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n743), .A2(G141gat), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT58), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n873), .A2(KEYINPUT121), .A3(new_n709), .A4(new_n874), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n875), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n630), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n755), .B1(new_n919), .B2(new_n886), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n690), .B1(new_n920), .B2(new_n888), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT122), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n923), .B(new_n690), .C1(new_n920), .C2(new_n888), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n922), .A2(new_n884), .A3(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT57), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n456), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n883), .A2(new_n891), .A3(new_n457), .ZN(new_n928));
  XNOR2_X1  g727(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n929));
  AOI22_X1  g728(.A1(new_n925), .A2(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n737), .A2(new_n894), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n930), .A2(new_n743), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n915), .B1(new_n932), .B2(new_n426), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n934), .B1(new_n930), .B2(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n928), .A2(new_n929), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n924), .A2(new_n884), .ZN(new_n937));
  AOI22_X1  g736(.A1(new_n628), .A2(new_n629), .B1(new_n875), .B2(new_n917), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n866), .B1(new_n938), .B2(new_n916), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n880), .B1(new_n939), .B2(new_n755), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n923), .B1(new_n940), .B2(new_n690), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n927), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n936), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n943), .A2(KEYINPUT123), .A3(new_n737), .A4(new_n894), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n935), .A2(new_n944), .A3(new_n626), .ZN(new_n945));
  INV_X1    g744(.A(new_n426), .ZN(new_n946));
  AOI22_X1  g745(.A1(new_n945), .A2(new_n946), .B1(new_n913), .B2(new_n914), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT58), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n933), .B1(new_n947), .B2(new_n948), .ZN(G1344gat));
  NAND3_X1  g748(.A1(new_n935), .A2(new_n944), .A3(new_n718), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n364), .A2(KEYINPUT59), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n928), .A2(new_n929), .ZN(new_n953));
  AOI22_X1  g752(.A1(new_n940), .A2(new_n690), .B1(new_n743), .B2(new_n719), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n926), .B1(new_n954), .B2(new_n456), .ZN(new_n955));
  AOI211_X1 g754(.A(new_n800), .B(new_n931), .C1(new_n953), .C2(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(KEYINPUT59), .B1(new_n956), .B2(new_n364), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n952), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n913), .A2(new_n364), .A3(new_n718), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1345gat));
  AOI21_X1  g759(.A(G155gat), .B1(new_n913), .B2(new_n691), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n935), .A2(new_n944), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n690), .A2(new_n686), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT124), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n961), .B1(new_n962), .B2(new_n964), .ZN(G1346gat));
  NAND2_X1  g764(.A1(new_n962), .A2(new_n755), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G162gat), .ZN(new_n967));
  INV_X1    g766(.A(G162gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n913), .A2(new_n968), .A3(new_n755), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1347gat));
  NOR2_X1   g769(.A1(new_n722), .A2(new_n522), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n893), .A2(new_n563), .A3(new_n971), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n972), .A2(new_n248), .A3(new_n743), .ZN(new_n973));
  NOR4_X1   g772(.A1(new_n892), .A2(new_n722), .A3(new_n522), .A4(new_n564), .ZN(new_n974));
  AOI21_X1  g773(.A(G169gat), .B1(new_n974), .B2(new_n626), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n973), .A2(new_n975), .ZN(G1348gat));
  OAI21_X1  g775(.A(G176gat), .B1(new_n972), .B2(new_n800), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n974), .A2(new_n249), .A3(new_n718), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(G1349gat));
  OAI21_X1  g778(.A(G183gat), .B1(new_n972), .B2(new_n690), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n691), .A2(new_n253), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT125), .ZN(new_n982));
  AOI22_X1  g781(.A1(new_n974), .A2(new_n981), .B1(new_n982), .B2(KEYINPUT60), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n982), .A2(KEYINPUT60), .ZN(new_n985));
  XOR2_X1   g784(.A(new_n984), .B(new_n985), .Z(G1350gat));
  NAND3_X1  g785(.A1(new_n974), .A2(new_n255), .A3(new_n755), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n972), .A2(new_n661), .ZN(new_n988));
  NOR2_X1   g787(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n255), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n989), .B1(new_n988), .B2(new_n990), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n987), .B1(new_n992), .B2(new_n993), .ZN(G1351gat));
  NOR2_X1   g793(.A1(new_n892), .A2(new_n722), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n912), .A2(new_n522), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g797(.A(G197gat), .B1(new_n998), .B2(new_n626), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n737), .A2(new_n971), .ZN(new_n1000));
  XNOR2_X1  g799(.A(new_n1000), .B(KEYINPUT127), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n1001), .B1(new_n953), .B2(new_n955), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n743), .A2(new_n387), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n999), .B1(new_n1002), .B2(new_n1003), .ZN(G1352gat));
  NAND2_X1  g803(.A1(new_n718), .A2(new_n384), .ZN(new_n1005));
  OAI21_X1  g804(.A(KEYINPUT62), .B1(new_n997), .B2(new_n1005), .ZN(new_n1006));
  OR3_X1    g805(.A1(new_n997), .A2(KEYINPUT62), .A3(new_n1005), .ZN(new_n1007));
  AND2_X1   g806(.A1(new_n1002), .A2(new_n718), .ZN(new_n1008));
  OAI211_X1 g807(.A(new_n1006), .B(new_n1007), .C1(new_n1008), .C2(new_n384), .ZN(G1353gat));
  INV_X1    g808(.A(G211gat), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n953), .A2(new_n955), .ZN(new_n1011));
  NOR2_X1   g810(.A1(new_n1000), .A2(new_n690), .ZN(new_n1012));
  AOI21_X1  g811(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g812(.A(new_n1013), .B(KEYINPUT63), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n998), .A2(new_n1010), .A3(new_n691), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1014), .A2(new_n1015), .ZN(G1354gat));
  AOI21_X1  g815(.A(G218gat), .B1(new_n998), .B2(new_n755), .ZN(new_n1017));
  NOR2_X1   g816(.A1(new_n661), .A2(new_n652), .ZN(new_n1018));
  AOI21_X1  g817(.A(new_n1017), .B1(new_n1002), .B2(new_n1018), .ZN(G1355gat));
endmodule


