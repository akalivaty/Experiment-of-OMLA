//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT64), .B1(new_n188), .B2(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(KEYINPUT64), .A3(G143), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n191), .A2(new_n192), .A3(G128), .A4(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  OAI21_X1  g010(.A(G128), .B1(new_n196), .B2(new_n192), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n190), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G137), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT11), .A3(G134), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(G137), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n204), .A2(new_n206), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n203), .A2(G137), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n205), .A2(G134), .ZN(new_n211));
  OAI21_X1  g025(.A(G131), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n201), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n204), .A2(new_n206), .A3(new_n208), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G131), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT65), .A3(new_n209), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n218), .A3(G131), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT0), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n221), .B1(new_n199), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(new_n195), .B2(G146), .ZN(new_n225));
  OAI211_X1 g039(.A(G128), .B(new_n193), .C1(new_n225), .C2(new_n196), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n199), .A2(G128), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n223), .A2(new_n226), .B1(new_n227), .B2(new_n221), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n214), .B1(new_n220), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT30), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT2), .ZN(new_n232));
  INV_X1    g046(.A(G113), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n233), .A3(KEYINPUT66), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(KEYINPUT2), .B2(G113), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(KEYINPUT2), .A2(G113), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(KEYINPUT67), .A2(G116), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT67), .A2(G116), .ZN(new_n241));
  OAI21_X1  g055(.A(G119), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G116), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(G119), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n239), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n237), .A2(new_n242), .A3(new_n238), .A4(new_n245), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n223), .A2(new_n226), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n227), .A2(new_n221), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(new_n219), .A3(new_n217), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT30), .A3(new_n214), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n231), .A2(new_n249), .A3(new_n254), .ZN(new_n255));
  AND4_X1   g069(.A1(new_n237), .A2(new_n242), .A3(new_n238), .A4(new_n245), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n237), .A2(new_n238), .B1(new_n242), .B2(new_n245), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n258), .B(new_n214), .C1(new_n220), .C2(new_n228), .ZN(new_n259));
  NOR2_X1   g073(.A1(G237), .A2(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G210), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n255), .A2(new_n259), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT31), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT31), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n255), .A2(new_n267), .A3(new_n259), .A4(new_n264), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT28), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n259), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n253), .A2(KEYINPUT28), .A3(new_n258), .A4(new_n214), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n229), .A2(new_n249), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT68), .ZN(new_n274));
  INV_X1    g088(.A(new_n264), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n274), .B1(new_n273), .B2(new_n275), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n266), .B(new_n268), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n273), .A2(new_n275), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT68), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n266), .A4(new_n268), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(G472), .A2(G902), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT70), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n289));
  INV_X1    g103(.A(new_n287), .ZN(new_n290));
  AOI211_X1 g104(.A(new_n289), .B(new_n290), .C1(new_n279), .C2(new_n285), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n187), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n290), .B1(new_n279), .B2(new_n285), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT32), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n272), .A2(new_n296), .A3(new_n259), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n229), .A2(KEYINPUT71), .A3(new_n249), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(KEYINPUT28), .A3(new_n298), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n299), .A2(KEYINPUT29), .A3(new_n264), .A4(new_n270), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n255), .A2(new_n259), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n275), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n273), .A2(new_n275), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n295), .B(new_n300), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G472), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n292), .A2(new_n294), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G101), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n310));
  INV_X1    g124(.A(G107), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n311), .A3(G104), .ZN(new_n312));
  INV_X1    g126(.A(G104), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT3), .B1(new_n313), .B2(G107), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(G107), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n309), .B(new_n312), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n311), .A2(G104), .ZN(new_n317));
  OAI21_X1  g131(.A(G101), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n242), .A2(KEYINPUT5), .A3(new_n245), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT5), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n233), .B1(new_n244), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(new_n324), .A3(new_n248), .ZN(new_n325));
  XNOR2_X1  g139(.A(G110), .B(G122), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G101), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(KEYINPUT4), .A3(new_n316), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n330), .A3(G101), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n325), .B(new_n326), .C1(new_n332), .C2(new_n258), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT6), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n249), .A2(new_n331), .A3(new_n329), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n326), .B1(new_n335), .B2(new_n325), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT82), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n325), .ZN(new_n338));
  INV_X1    g152(.A(new_n326), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT82), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT6), .A4(new_n333), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT83), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n340), .B2(KEYINPUT6), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT6), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n336), .A2(KEYINPUT83), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n201), .A2(G125), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(G125), .B2(new_n228), .ZN(new_n350));
  INV_X1    g164(.A(G224), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(G953), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n350), .B(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n343), .A2(new_n348), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n350), .A2(KEYINPUT7), .A3(new_n353), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n324), .A2(new_n248), .A3(new_n319), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n326), .B(KEYINPUT8), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n323), .B(KEYINPUT84), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n256), .B1(new_n359), .B2(new_n321), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n357), .B(new_n358), .C1(new_n360), .C2(new_n319), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n356), .A2(new_n333), .A3(new_n361), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n349), .A2(KEYINPUT85), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n349), .A2(KEYINPUT85), .ZN(new_n364));
  INV_X1    g178(.A(G125), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n363), .B(new_n364), .C1(new_n365), .C2(new_n252), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT7), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n366), .B1(new_n367), .B2(new_n352), .ZN(new_n368));
  AOI21_X1  g182(.A(G902), .B1(new_n362), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n355), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G210), .B1(G237), .B2(G902), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n355), .A2(new_n369), .A3(new_n371), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G214), .B1(G237), .B2(G902), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT81), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n243), .A2(G122), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT67), .B(G116), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(G122), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT90), .B(G107), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G122), .ZN(new_n385));
  INV_X1    g199(.A(new_n241), .ZN(new_n386));
  NAND2_X1  g200(.A1(KEYINPUT67), .A2(G116), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n382), .B1(new_n388), .B2(new_n379), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT92), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n195), .A2(G128), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n222), .A2(G143), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT91), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT91), .B1(new_n392), .B2(new_n393), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n203), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT13), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n393), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n392), .A2(new_n398), .ZN(new_n401));
  OAI21_X1  g215(.A(G134), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n390), .A2(new_n391), .A3(new_n397), .A4(new_n402), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n397), .A2(new_n384), .A3(new_n402), .A4(new_n389), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT92), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n407));
  OAI21_X1  g221(.A(G107), .B1(new_n379), .B2(new_n407), .ZN(new_n408));
  XOR2_X1   g222(.A(new_n381), .B(new_n408), .Z(new_n409));
  OR3_X1    g223(.A1(new_n395), .A2(new_n203), .A3(new_n396), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n397), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  XOR2_X1   g226(.A(KEYINPUT9), .B(G234), .Z(new_n413));
  INV_X1    g227(.A(G953), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(G217), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n406), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n416), .B1(new_n406), .B2(new_n412), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n295), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT15), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n420), .A3(G478), .ZN(new_n421));
  INV_X1    g235(.A(G478), .ZN(new_n422));
  OAI221_X1 g236(.A(new_n295), .B1(KEYINPUT15), .B2(new_n422), .C1(new_n417), .C2(new_n418), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(G234), .A2(G237), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(G952), .A3(new_n414), .ZN(new_n426));
  XOR2_X1   g240(.A(KEYINPUT21), .B(G898), .Z(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(G902), .A3(G953), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G237), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n414), .A3(G214), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(G143), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n432), .B1(new_n433), .B2(new_n207), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n431), .B(new_n195), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(KEYINPUT18), .A3(G131), .ZN(new_n436));
  INV_X1    g250(.A(G140), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G125), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n365), .A2(G140), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(G146), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT86), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n188), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n434), .B(new_n436), .C1(new_n441), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n435), .A2(G131), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n432), .A2(new_n207), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT17), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n435), .A2(KEYINPUT17), .A3(G131), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT16), .ZN(new_n453));
  OR3_X1    g267(.A1(new_n365), .A2(KEYINPUT16), .A3(G140), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT75), .B1(new_n455), .B2(G146), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(KEYINPUT74), .A3(G146), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n453), .A2(new_n454), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT75), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n188), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n453), .A2(new_n454), .A3(G146), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT74), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n456), .A2(new_n457), .A3(new_n460), .A4(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n446), .B1(new_n452), .B2(new_n464), .ZN(new_n465));
  XOR2_X1   g279(.A(KEYINPUT87), .B(G104), .Z(new_n466));
  XNOR2_X1  g280(.A(G113), .B(G122), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n446), .A2(new_n468), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT76), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n461), .B(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n447), .A2(new_n448), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n443), .A2(new_n444), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT19), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(KEYINPUT19), .B2(new_n440), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n473), .B(new_n474), .C1(new_n477), .C2(G146), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(G475), .A2(G902), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n480), .B(KEYINPUT88), .Z(new_n481));
  NAND3_X1  g295(.A1(new_n470), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT20), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n465), .A2(new_n469), .B1(new_n471), .B2(new_n478), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT20), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n481), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n468), .A2(KEYINPUT89), .ZN(new_n487));
  AOI21_X1  g301(.A(G902), .B1(new_n465), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(new_n487), .B2(new_n465), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n483), .A2(new_n486), .B1(new_n489), .B2(G475), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n424), .A2(new_n429), .A3(new_n490), .ZN(new_n491));
  OR2_X1    g305(.A1(new_n378), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G469), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n193), .B1(new_n225), .B2(new_n196), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n197), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n194), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n320), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT10), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n252), .A2(new_n331), .A3(new_n329), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n320), .A2(new_n201), .A3(KEYINPUT10), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n499), .A2(new_n220), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(G110), .B(G140), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n414), .A2(G227), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n503), .B(new_n504), .Z(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n217), .A2(new_n219), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT79), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(KEYINPUT12), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n319), .A2(new_n194), .A3(new_n200), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n319), .B1(new_n194), .B2(new_n495), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n507), .B(new_n509), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n220), .B1(new_n497), .B2(new_n510), .ZN(new_n514));
  XOR2_X1   g328(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n515));
  OAI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n506), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n500), .A2(new_n501), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n512), .A2(KEYINPUT10), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n507), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n505), .B1(new_n520), .B2(new_n502), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n493), .B(new_n295), .C1(new_n517), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(G469), .A2(G902), .ZN(new_n523));
  INV_X1    g337(.A(new_n505), .ZN(new_n524));
  INV_X1    g338(.A(new_n502), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n524), .B1(new_n516), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n520), .A2(new_n502), .A3(new_n505), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(G469), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n522), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G221), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n530), .B1(new_n413), .B2(new_n295), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT80), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n492), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G217), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n537), .B1(G234), .B2(new_n295), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT22), .B(G137), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n414), .A2(G221), .A3(G234), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XOR2_X1   g355(.A(G119), .B(G128), .Z(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT24), .B(G110), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT23), .B1(new_n222), .B2(G119), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT72), .B1(new_n222), .B2(G119), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G119), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(G128), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT72), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT23), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(KEYINPUT73), .B(G110), .C1(new_n547), .C2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT73), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n545), .A2(new_n546), .B1(new_n549), .B2(new_n552), .ZN(new_n556));
  INV_X1    g370(.A(G110), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n544), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n557), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n542), .A2(new_n543), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n441), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n464), .A2(new_n559), .B1(new_n473), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n541), .B1(new_n563), .B2(KEYINPUT77), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n464), .A2(new_n559), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n473), .A2(new_n562), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT77), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(new_n568), .A3(new_n541), .ZN(new_n571));
  AOI21_X1  g385(.A(G902), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT25), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n538), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI211_X1 g388(.A(KEYINPUT25), .B(G902), .C1(new_n570), .C2(new_n571), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n570), .A2(new_n571), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n538), .A2(G902), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT78), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT78), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n577), .A2(new_n581), .A3(new_n578), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n308), .A2(new_n536), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G101), .ZN(G3));
  NAND2_X1  g400(.A1(new_n286), .A2(new_n295), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(G472), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n534), .B(new_n588), .C1(new_n288), .C2(new_n291), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n576), .A2(new_n583), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n376), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n592), .B1(new_n373), .B2(new_n374), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n429), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n419), .A2(new_n422), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n417), .B2(new_n418), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n406), .A2(new_n412), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n415), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n406), .A2(new_n412), .A3(new_n416), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(KEYINPUT33), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n422), .A2(G902), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n483), .A2(new_n486), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n489), .A2(G475), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n595), .A2(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n594), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n591), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT34), .B(G104), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G6));
  NAND2_X1  g425(.A1(new_n421), .A2(new_n423), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n490), .ZN(new_n613));
  NOR4_X1   g427(.A1(new_n589), .A2(new_n590), .A3(new_n594), .A4(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT35), .B(G107), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  INV_X1    g430(.A(new_n589), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT36), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n541), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n563), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n578), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n574), .B2(new_n575), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n492), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT37), .B(G110), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G12));
  NOR2_X1   g441(.A1(new_n533), .A2(KEYINPUT80), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT80), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n529), .B2(new_n532), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n622), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n613), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n426), .B(KEYINPUT93), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(G900), .B2(new_n428), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n308), .A2(new_n593), .A3(new_n632), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G128), .ZN(G30));
  NAND2_X1  g454(.A1(new_n301), .A2(new_n264), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n295), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n264), .B1(new_n297), .B2(new_n298), .ZN(new_n643));
  OAI21_X1  g457(.A(G472), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n292), .A2(new_n294), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT94), .ZN(new_n646));
  OR2_X1    g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n636), .B(KEYINPUT39), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n534), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT95), .B(KEYINPUT40), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n534), .A2(new_n648), .A3(new_n651), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n375), .B(KEYINPUT38), .ZN(new_n654));
  NOR4_X1   g468(.A1(new_n622), .A2(new_n592), .A3(new_n424), .A4(new_n490), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n645), .A2(new_n646), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n647), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT96), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n647), .A2(new_n657), .A3(KEYINPUT96), .A4(new_n658), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n195), .ZN(G45));
  NAND2_X1  g478(.A1(new_n603), .A2(new_n595), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n604), .A2(new_n605), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n666), .A3(new_n636), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT97), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT97), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n606), .A2(new_n669), .A3(new_n636), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n375), .A2(new_n376), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n631), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n308), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT98), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT98), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n308), .A2(new_n676), .A3(new_n673), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  OR2_X1    g493(.A1(new_n517), .A2(new_n521), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n295), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(G469), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n532), .A3(new_n522), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n308), .A2(new_n584), .A3(new_n608), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G15));
  NOR2_X1   g501(.A1(new_n672), .A2(new_n683), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n688), .A2(new_n429), .A3(new_n633), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n308), .A2(new_n584), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G116), .ZN(G18));
  AND2_X1   g505(.A1(new_n682), .A2(new_n522), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n593), .A3(new_n532), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n693), .A2(new_n491), .A3(new_n623), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n308), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G119), .ZN(G21));
  OAI21_X1  g510(.A(KEYINPUT102), .B1(new_n424), .B2(new_n490), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n612), .A2(new_n666), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n593), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT103), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n593), .A2(new_n697), .A3(new_n702), .A4(new_n699), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n287), .B(KEYINPUT99), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n299), .A2(KEYINPUT100), .A3(new_n270), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT100), .B1(new_n299), .B2(new_n270), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n707), .A2(new_n708), .A3(new_n264), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n266), .A2(new_n268), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n705), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(G902), .B1(new_n279), .B2(new_n285), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT101), .B(G472), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n584), .B(new_n711), .C1(new_n712), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n684), .A2(new_n429), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n704), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  NOR2_X1   g533(.A1(new_n708), .A2(new_n264), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n706), .ZN(new_n721));
  INV_X1    g535(.A(new_n710), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n587), .A2(new_n713), .B1(new_n723), .B2(new_n705), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n668), .A2(new_n670), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(new_n725), .A3(new_n688), .A4(new_n622), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n711), .B(new_n622), .C1(new_n712), .C2(new_n714), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n671), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(KEYINPUT104), .A3(new_n688), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n293), .A2(KEYINPUT32), .B1(G472), .B2(new_n306), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n286), .A2(new_n287), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n187), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n734), .B1(new_n738), .B2(new_n584), .ZN(new_n739));
  AOI211_X1 g553(.A(KEYINPUT108), .B(new_n590), .C1(new_n735), .C2(new_n737), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n529), .A2(new_n742), .A3(new_n532), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n742), .B1(new_n529), .B2(new_n532), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n373), .A2(KEYINPUT106), .A3(new_n374), .A4(new_n376), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n745), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT107), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n745), .A2(new_n748), .A3(new_n752), .A4(new_n749), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n725), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT42), .B1(new_n741), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n308), .A2(new_n584), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n671), .A2(KEYINPUT42), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n754), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n207), .ZN(G33));
  AND4_X1   g575(.A1(new_n308), .A2(new_n754), .A3(new_n584), .A4(new_n638), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n203), .ZN(G36));
  NAND3_X1  g577(.A1(new_n526), .A2(KEYINPUT45), .A3(new_n527), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n526), .A2(new_n527), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n764), .A2(G469), .A3(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n768), .A2(new_n523), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n769), .A2(KEYINPUT46), .ZN(new_n770));
  INV_X1    g584(.A(new_n522), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n769), .B2(KEYINPUT46), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n531), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n648), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n588), .B1(new_n288), .B2(new_n291), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n665), .A2(new_n490), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT43), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT43), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n623), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n748), .A2(new_n749), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n776), .A2(new_n782), .A3(KEYINPUT44), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n775), .A2(new_n785), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  NOR3_X1   g604(.A1(new_n786), .A2(new_n584), .A3(new_n671), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n292), .A3(new_n294), .A4(new_n307), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n792), .A2(KEYINPUT109), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(KEYINPUT109), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n773), .B(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT110), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT110), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n800), .B(new_n797), .C1(new_n793), .C2(new_n794), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(new_n437), .ZN(G42));
  AND3_X1   g617(.A1(new_n308), .A2(new_n676), .A3(new_n673), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n676), .B1(new_n308), .B2(new_n673), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n639), .B(new_n732), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n636), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n622), .A2(new_n533), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT113), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n645), .A2(new_n704), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT52), .B1(new_n806), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n732), .A2(new_n639), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n814), .A3(new_n678), .A4(new_n810), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT42), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n294), .A2(new_n307), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n293), .A2(KEYINPUT32), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n584), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT108), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n738), .A2(new_n734), .A3(new_n584), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n671), .B1(new_n751), .B2(new_n753), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n816), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AND4_X1   g638(.A1(new_n308), .A2(new_n754), .A3(new_n584), .A4(new_n758), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n824), .A2(new_n825), .A3(new_n762), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n685), .A2(new_n690), .A3(new_n695), .A4(new_n718), .ZN(new_n827));
  INV_X1    g641(.A(new_n776), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n607), .A2(new_n613), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n375), .A2(new_n829), .A3(new_n377), .A4(new_n429), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n828), .A2(new_n584), .A3(new_n534), .A4(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n585), .A2(new_n831), .A3(new_n625), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n754), .A2(new_n730), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n424), .A2(new_n490), .A3(new_n636), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT112), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n786), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n308), .A2(new_n632), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n827), .A2(new_n832), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n812), .A2(new_n815), .A3(new_n826), .A4(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n757), .A2(new_n638), .A3(new_n754), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT53), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n591), .A2(new_n830), .B1(new_n617), .B2(new_n624), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(new_n585), .A3(new_n833), .A4(new_n837), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n760), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n827), .B(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n848), .A2(new_n815), .A3(new_n850), .A4(new_n812), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n842), .A2(new_n843), .A3(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n826), .A2(new_n839), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(KEYINPUT53), .A3(new_n815), .A4(new_n812), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n843), .B1(new_n854), .B2(new_n842), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT115), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n842), .A2(new_n851), .A3(new_n843), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n635), .B1(new_n779), .B2(new_n781), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n724), .A3(new_n584), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT116), .B1(new_n684), .B2(new_n592), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n684), .A2(KEYINPUT116), .A3(new_n592), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n862), .A2(new_n863), .A3(new_n654), .A4(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT50), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n862), .A2(new_n786), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n692), .B(KEYINPUT111), .Z(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n532), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n867), .B1(new_n798), .B2(new_n869), .ZN(new_n870));
  OR3_X1    g684(.A1(new_n786), .A2(KEYINPUT117), .A3(new_n683), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT117), .B1(new_n786), .B2(new_n683), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n873), .A2(new_n861), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n622), .A3(new_n724), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n866), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n590), .B1(new_n647), .B2(new_n658), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n426), .B1(new_n871), .B2(new_n872), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n665), .A2(new_n666), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n876), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(KEYINPUT51), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n886));
  AOI211_X1 g700(.A(new_n886), .B(new_n876), .C1(new_n882), .C2(new_n883), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT48), .B1(new_n874), .B2(new_n822), .ZN(new_n888));
  OAI211_X1 g702(.A(G952), .B(new_n414), .C1(new_n862), .C2(new_n693), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n877), .A2(new_n606), .A3(new_n878), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n874), .A2(KEYINPUT48), .A3(new_n822), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OR3_X1    g707(.A1(new_n885), .A2(new_n887), .A3(new_n893), .ZN(new_n894));
  OAI22_X1  g708(.A1(new_n860), .A2(new_n894), .B1(G952), .B2(G953), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n778), .A2(new_n377), .A3(new_n532), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(new_n868), .B2(KEYINPUT49), .ZN(new_n897));
  AOI211_X1 g711(.A(new_n654), .B(new_n897), .C1(KEYINPUT49), .C2(new_n868), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n877), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n895), .A2(new_n899), .ZN(G75));
  AOI21_X1  g714(.A(new_n295), .B1(new_n842), .B2(new_n851), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT56), .B1(new_n901), .B2(G210), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n343), .A2(new_n348), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n354), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n902), .A2(new_n905), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n414), .A2(G952), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(G51));
  AOI211_X1 g723(.A(new_n295), .B(new_n768), .C1(new_n842), .C2(new_n851), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n523), .B(KEYINPUT57), .Z(new_n911));
  AOI21_X1  g725(.A(new_n843), .B1(new_n842), .B2(new_n851), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n911), .B1(new_n852), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n910), .B1(new_n913), .B2(new_n680), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT119), .B1(new_n914), .B2(new_n908), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n916));
  INV_X1    g730(.A(new_n908), .ZN(new_n917));
  INV_X1    g731(.A(new_n680), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n842), .A2(new_n851), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT54), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n857), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n918), .B1(new_n921), .B2(new_n911), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n916), .B(new_n917), .C1(new_n922), .C2(new_n910), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n915), .A2(new_n923), .ZN(G54));
  AND2_X1   g738(.A1(KEYINPUT58), .A2(G475), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n901), .A2(new_n484), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n484), .B1(new_n901), .B2(new_n925), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n908), .ZN(G60));
  INV_X1    g742(.A(new_n921), .ZN(new_n929));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT59), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n597), .A2(new_n601), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n917), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n860), .A2(new_n931), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n597), .A2(new_n601), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(G63));
  XNOR2_X1  g750(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n537), .A2(new_n295), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n919), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n577), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n908), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT61), .B1(new_n942), .B2(KEYINPUT122), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n620), .B(KEYINPUT121), .Z(new_n944));
  NAND3_X1  g758(.A1(new_n919), .A2(new_n939), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n942), .B(new_n945), .C1(KEYINPUT122), .C2(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(G66));
  INV_X1    g763(.A(new_n427), .ZN(new_n950));
  OAI21_X1  g764(.A(G953), .B1(new_n950), .B2(new_n351), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n827), .A2(new_n832), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n903), .B1(G898), .B2(new_n414), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G69));
  NAND2_X1  g769(.A1(new_n231), .A2(new_n254), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(new_n477), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n799), .A2(new_n801), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT123), .ZN(new_n960));
  INV_X1    g774(.A(new_n806), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n661), .A3(new_n662), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n959), .A2(KEYINPUT123), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n960), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n961), .A2(new_n661), .A3(new_n662), .A4(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n757), .A2(new_n649), .A3(new_n787), .A4(new_n829), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n789), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n967), .A2(new_n789), .A3(KEYINPUT124), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n958), .A2(new_n964), .A3(new_n966), .A4(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n957), .B1(new_n973), .B2(new_n414), .ZN(new_n974));
  INV_X1    g788(.A(new_n957), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(G900), .B2(G953), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n822), .A2(new_n775), .A3(new_n704), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n961), .A2(new_n826), .A3(new_n789), .A4(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n802), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n977), .B1(new_n980), .B2(new_n414), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT126), .B1(new_n974), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n802), .A2(new_n979), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n976), .B1(new_n984), .B2(G953), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n970), .B(new_n971), .C1(new_n799), .C2(new_n801), .ZN(new_n986));
  INV_X1    g800(.A(new_n966), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(G953), .B1(new_n988), .B2(new_n964), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n983), .B(new_n985), .C1(new_n989), .C2(new_n957), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n975), .A2(KEYINPUT125), .ZN(new_n991));
  AOI211_X1 g805(.A(new_n414), .B(new_n991), .C1(G227), .C2(G900), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n982), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n992), .B1(new_n982), .B2(new_n990), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(G72));
  NAND2_X1  g809(.A1(new_n980), .A2(new_n952), .ZN(new_n996));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT63), .Z(new_n998));
  AOI211_X1 g812(.A(new_n301), .B(new_n264), .C1(new_n996), .C2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n988), .A2(new_n952), .A3(new_n964), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n641), .B1(new_n1000), .B2(new_n998), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n302), .B(KEYINPUT127), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n265), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n998), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(new_n854), .B2(new_n842), .ZN(new_n1005));
  NOR4_X1   g819(.A1(new_n999), .A2(new_n1001), .A3(new_n908), .A4(new_n1005), .ZN(G57));
endmodule


