//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n638, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n467), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n465), .A2(G2105), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT70), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n473), .A2(G137), .B1(G101), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n469), .A2(new_n466), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n469), .B2(new_n466), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G125), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT68), .B1(new_n481), .B2(new_n482), .ZN(new_n486));
  NAND2_X1  g061(.A1(G113), .A2(G2104), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n477), .B1(new_n488), .B2(G2105), .ZN(G160));
  INV_X1    g064(.A(G136), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n472), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT71), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n494));
  XOR2_X1   g069(.A(new_n494), .B(KEYINPUT72), .Z(new_n495));
  NAND3_X1  g070(.A1(new_n467), .A2(G2105), .A3(new_n471), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n495), .B1(G124), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g074(.A(new_n499), .B(KEYINPUT73), .ZN(G162));
  INV_X1    g075(.A(KEYINPUT74), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n468), .B2(G114), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT74), .A3(G2105), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G126), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n496), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G138), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT4), .B1(new_n472), .B2(new_n511), .ZN(new_n512));
  NOR3_X1   g087(.A1(new_n511), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n513), .B1(new_n479), .B2(new_n480), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n510), .B1(new_n512), .B2(new_n514), .ZN(G164));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G62), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT78), .Z(new_n523));
  AOI21_X1  g098(.A(new_n516), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G50), .ZN(new_n525));
  AND2_X1   g100(.A1(KEYINPUT75), .A2(KEYINPUT6), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT75), .A2(KEYINPUT6), .ZN(new_n527));
  OAI21_X1  g102(.A(G651), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT76), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n530), .B(G651), .C1(new_n526), .C2(new_n527), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n516), .A2(KEYINPUT6), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n529), .A2(G543), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n529), .A2(new_n520), .A3(new_n531), .A4(new_n532), .ZN(new_n534));
  INV_X1    g109(.A(G88), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n525), .A2(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(KEYINPUT77), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(KEYINPUT77), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n524), .B1(new_n537), .B2(new_n538), .ZN(G166));
  XOR2_X1   g114(.A(KEYINPUT79), .B(KEYINPUT7), .Z(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(G63), .A2(G651), .ZN(new_n543));
  INV_X1    g118(.A(G51), .ZN(new_n544));
  OAI221_X1 g119(.A(new_n542), .B1(new_n519), .B2(new_n543), .C1(new_n533), .C2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n534), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n546), .A2(G89), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n545), .A2(new_n547), .ZN(G168));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G64), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n519), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n546), .A2(G90), .B1(G651), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n533), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G52), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n519), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G651), .ZN(new_n560));
  INV_X1    g135(.A(G81), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n534), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(G43), .B2(new_n553), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  AND3_X1   g139(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(G188));
  AND3_X1   g144(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n570), .A2(new_n571), .A3(G53), .A4(G543), .ZN(new_n572));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT80), .B1(new_n533), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(KEYINPUT9), .A3(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT81), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n534), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n532), .ZN(new_n578));
  OR2_X1    g153(.A1(KEYINPUT75), .A2(KEYINPUT6), .ZN(new_n579));
  NAND2_X1  g154(.A1(KEYINPUT75), .A2(KEYINPUT6), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n516), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n578), .B1(new_n581), .B2(new_n530), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n582), .A2(KEYINPUT81), .A3(new_n520), .A4(new_n529), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n577), .A2(G91), .A3(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n520), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(new_n516), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT9), .ZN(new_n587));
  OAI211_X1 g162(.A(KEYINPUT80), .B(new_n587), .C1(new_n533), .C2(new_n573), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n575), .A2(new_n584), .A3(new_n586), .A4(new_n588), .ZN(G299));
  INV_X1    g164(.A(G168), .ZN(G286));
  INV_X1    g165(.A(G166), .ZN(G303));
  AND2_X1   g166(.A1(new_n577), .A2(new_n583), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G87), .ZN(new_n593));
  INV_X1    g168(.A(G74), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n516), .B1(new_n519), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n570), .A2(KEYINPUT82), .A3(G49), .A4(G543), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT82), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n582), .A2(new_n529), .ZN(new_n598));
  NAND2_X1  g173(.A1(G49), .A2(G543), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n595), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n593), .A2(new_n601), .ZN(G288));
  NAND2_X1  g177(.A1(new_n592), .A2(G86), .ZN(new_n603));
  INV_X1    g178(.A(G61), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n519), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(G73), .A2(G543), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n605), .B2(new_n606), .ZN(new_n610));
  OAI21_X1  g185(.A(G651), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n553), .A2(G48), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n603), .A2(new_n611), .A3(new_n612), .ZN(G305));
  AOI22_X1  g188(.A1(G47), .A2(new_n553), .B1(new_n546), .B2(G85), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(KEYINPUT84), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(KEYINPUT84), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(G72), .A2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G60), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n519), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G651), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n617), .A2(new_n621), .ZN(G290));
  NAND2_X1  g197(.A1(G301), .A2(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(G79), .A2(G543), .ZN(new_n624));
  INV_X1    g199(.A(G66), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n519), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G651), .ZN(new_n627));
  INV_X1    g202(.A(G54), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n533), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n577), .A2(G92), .A3(new_n583), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT10), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g207(.A1(new_n577), .A2(new_n583), .A3(KEYINPUT10), .A4(G92), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n623), .B1(new_n634), .B2(G868), .ZN(G284));
  OAI21_X1  g210(.A(new_n623), .B1(new_n634), .B2(G868), .ZN(G321));
  NAND2_X1  g211(.A1(G286), .A2(G868), .ZN(new_n637));
  INV_X1    g212(.A(G299), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G868), .ZN(G297));
  OAI21_X1  g214(.A(new_n637), .B1(new_n638), .B2(G868), .ZN(G280));
  INV_X1    g215(.A(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n634), .B1(new_n641), .B2(G860), .ZN(G148));
  NAND2_X1  g217(.A1(new_n632), .A2(new_n633), .ZN(new_n643));
  INV_X1    g218(.A(new_n629), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(KEYINPUT85), .B1(new_n645), .B2(G559), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT85), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n634), .A2(new_n647), .A3(new_n641), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(G868), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n650), .A2(KEYINPUT86), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(KEYINPUT86), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n651), .B(new_n652), .C1(G868), .C2(new_n563), .ZN(G323));
  XNOR2_X1  g228(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g229(.A1(new_n479), .A2(new_n480), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(new_n475), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT12), .Z(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT13), .Z(new_n658));
  INV_X1    g233(.A(G2100), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  OR2_X1    g236(.A1(G99), .A2(G2105), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n662), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n663));
  INV_X1    g238(.A(G123), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n663), .B1(new_n496), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(G135), .B2(new_n473), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2096), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n660), .A2(new_n661), .A3(new_n667), .ZN(G156));
  XOR2_X1   g243(.A(G2451), .B(G2454), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT16), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1341), .B(G1348), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT14), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2427), .B(G2438), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2430), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT15), .B(G2435), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(new_n676), .B2(new_n675), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n672), .B(new_n678), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2443), .B(G2446), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(G14), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n682), .B2(new_n680), .ZN(G401));
  XOR2_X1   g259(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n685));
  XOR2_X1   g260(.A(G2084), .B(G2090), .Z(new_n686));
  XNOR2_X1  g261(.A(G2067), .B(G2678), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(KEYINPUT17), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n686), .A2(new_n687), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n685), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G2072), .B(G2078), .Z(new_n692));
  INV_X1    g267(.A(new_n685), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n692), .B1(new_n688), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n691), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G2096), .B(G2100), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G227));
  XOR2_X1   g272(.A(G1961), .B(G1966), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT88), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1956), .B(G2474), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1971), .B(G1976), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT19), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT20), .Z(new_n706));
  NOR2_X1   g281(.A1(new_n699), .A2(new_n701), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n708), .A2(new_n704), .A3(new_n702), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n706), .B(new_n709), .C1(new_n704), .C2(new_n708), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1991), .B(G1996), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1981), .B(G1986), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(G229));
  XOR2_X1   g291(.A(KEYINPUT89), .B(G29), .Z(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(G35), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G162), .B2(new_n718), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G2090), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT101), .Z(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G20), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT23), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n638), .B2(new_n724), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT102), .B(G1956), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT103), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(KEYINPUT103), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n655), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(new_n468), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT25), .Z(new_n736));
  INV_X1    g311(.A(G139), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n472), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT95), .Z(new_n740));
  MUX2_X1   g315(.A(G33), .B(new_n740), .S(G29), .Z(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(G2072), .Z(new_n742));
  NOR2_X1   g317(.A1(G171), .A2(new_n724), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G5), .B2(new_n724), .ZN(new_n744));
  INV_X1    g319(.A(G1961), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G34), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT96), .B(KEYINPUT24), .Z(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n718), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OAI22_X1  g326(.A1(new_n751), .A2(KEYINPUT97), .B1(new_n747), .B2(new_n749), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(KEYINPUT97), .B2(new_n751), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G160), .B2(G29), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n746), .B1(G2084), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G2084), .B2(new_n754), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n718), .A2(G27), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G164), .B2(new_n718), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2078), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n724), .A2(G21), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G168), .B2(new_n724), .ZN(new_n761));
  OAI22_X1  g336(.A1(new_n744), .A2(new_n745), .B1(G1966), .B2(new_n761), .ZN(new_n762));
  AOI211_X1 g337(.A(new_n759), .B(new_n762), .C1(G1966), .C2(new_n761), .ZN(new_n763));
  INV_X1    g338(.A(G29), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G32), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n497), .A2(G129), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT98), .Z(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT26), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n475), .A2(G105), .ZN(new_n770));
  AOI211_X1 g345(.A(new_n769), .B(new_n770), .C1(G141), .C2(new_n473), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n765), .B1(new_n772), .B2(new_n764), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT27), .B(G1996), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n773), .A2(new_n775), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n666), .A2(new_n718), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT31), .B(G11), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G28), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT99), .Z(new_n782));
  OAI211_X1 g357(.A(new_n782), .B(new_n764), .C1(new_n780), .C2(G28), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n778), .A2(new_n779), .A3(new_n783), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT100), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n717), .A2(G26), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT28), .ZN(new_n787));
  OR2_X1    g362(.A1(G104), .A2(G2105), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n788), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n789));
  INV_X1    g364(.A(G128), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n496), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G140), .B2(new_n473), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n787), .B1(new_n792), .B2(new_n764), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2067), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n776), .A2(new_n777), .A3(new_n785), .A4(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n742), .A2(new_n756), .A3(new_n763), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(G4), .A2(G16), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n634), .B2(G16), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G1348), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n721), .B2(G2090), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n798), .A2(G1348), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n724), .A2(G19), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT93), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n563), .B2(new_n724), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT94), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(G1341), .Z(new_n806));
  NOR4_X1   g381(.A1(new_n796), .A2(new_n800), .A3(new_n801), .A4(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n731), .A2(new_n732), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n724), .A2(G6), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n612), .A2(new_n611), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n592), .B2(G86), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n809), .B1(new_n811), .B2(new_n724), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT91), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT32), .B(G1981), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n724), .A2(G23), .ZN(new_n816));
  INV_X1    g391(.A(G288), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n724), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT33), .B(G1976), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n724), .A2(G22), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G166), .B2(new_n724), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1971), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n815), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT92), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT92), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n815), .A2(new_n827), .A3(new_n824), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT34), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n826), .A2(KEYINPUT34), .A3(new_n828), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n615), .A2(new_n616), .B1(G651), .B2(new_n620), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G16), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G16), .B2(G24), .ZN(new_n835));
  INV_X1    g410(.A(G1986), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n718), .A2(G25), .ZN(new_n839));
  INV_X1    g414(.A(G119), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n468), .A2(G107), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n496), .A2(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(G131), .B2(new_n473), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n839), .B1(new_n844), .B2(new_n718), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT35), .B(G1991), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT90), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n845), .B(new_n847), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n837), .A2(new_n838), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n831), .A2(new_n832), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT36), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(KEYINPUT36), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n808), .B1(new_n851), .B2(new_n853), .ZN(G311));
  AND3_X1   g429(.A1(new_n731), .A2(new_n732), .A3(new_n807), .ZN(new_n855));
  INV_X1    g430(.A(new_n851), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n852), .B2(new_n856), .ZN(G150));
  NAND2_X1  g432(.A1(new_n634), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT38), .ZN(new_n859));
  INV_X1    g434(.A(G93), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n861));
  OAI22_X1  g436(.A1(new_n534), .A2(new_n860), .B1(new_n861), .B2(new_n516), .ZN(new_n862));
  INV_X1    g437(.A(G55), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n533), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G43), .ZN(new_n867));
  OAI221_X1 g442(.A(new_n560), .B1(new_n534), .B2(new_n561), .C1(new_n867), .C2(new_n533), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n563), .A2(new_n865), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n859), .B(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n874));
  INV_X1    g449(.A(G860), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n865), .A2(new_n875), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(G145));
  XNOR2_X1  g455(.A(new_n740), .B(new_n772), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n497), .A2(G130), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n468), .A2(G118), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(G142), .B2(new_n473), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n657), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n881), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n512), .A2(new_n514), .ZN(new_n889));
  INV_X1    g464(.A(new_n510), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n792), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n844), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n888), .B(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(G160), .B(new_n666), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(G162), .ZN(new_n896));
  AOI21_X1  g471(.A(G37), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n896), .B2(new_n894), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n634), .B(G299), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT41), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n645), .A2(G299), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n584), .A2(new_n586), .A3(new_n588), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n634), .A2(new_n575), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(KEYINPUT105), .A3(KEYINPUT41), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT104), .B1(new_n902), .B2(new_n903), .ZN(new_n910));
  AND4_X1   g485(.A1(KEYINPUT104), .A2(new_n905), .A3(new_n903), .A4(new_n907), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n904), .B(new_n909), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n649), .B(new_n872), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n913), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT106), .B1(new_n913), .B2(new_n908), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n900), .B(new_n915), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n916), .B(KEYINPUT106), .C1(new_n913), .C2(new_n908), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n900), .B1(new_n921), .B2(new_n915), .ZN(new_n922));
  NAND2_X1  g497(.A1(G290), .A2(G166), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n833), .A2(G303), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n817), .A2(G305), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n811), .A2(G288), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n925), .B(new_n928), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n920), .A2(new_n922), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n928), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n925), .B(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n917), .A2(new_n918), .ZN(new_n933));
  INV_X1    g508(.A(new_n915), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT42), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n932), .B1(new_n935), .B2(new_n919), .ZN(new_n936));
  OAI21_X1  g511(.A(G868), .B1(new_n930), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n865), .A2(G868), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(G295));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n937), .A2(new_n941), .A3(new_n939), .ZN(new_n942));
  INV_X1    g517(.A(G868), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n929), .B1(new_n920), .B2(new_n922), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n935), .A2(new_n932), .A3(new_n919), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT107), .B1(new_n946), .B2(new_n938), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n942), .A2(new_n947), .ZN(G331));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n949));
  NAND2_X1  g524(.A1(G301), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n871), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(G286), .B1(G171), .B2(KEYINPUT108), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n869), .A2(new_n950), .A3(new_n870), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n953), .B1(new_n952), .B2(new_n954), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n912), .A2(new_n958), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n955), .A2(new_n956), .A3(new_n908), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(new_n929), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n902), .A2(new_n903), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n908), .A2(KEYINPUT41), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(new_n957), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n932), .B1(new_n966), .B2(new_n960), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  INV_X1    g543(.A(G37), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n962), .A2(new_n967), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT105), .B1(new_n908), .B2(KEYINPUT41), .ZN(new_n973));
  AOI211_X1 g548(.A(new_n901), .B(new_n903), .C1(new_n905), .C2(new_n907), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(new_n908), .B2(KEYINPUT41), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n902), .A2(KEYINPUT104), .A3(new_n903), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n957), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n932), .B1(new_n980), .B2(new_n960), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(new_n962), .A3(new_n969), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n960), .B1(new_n912), .B2(new_n958), .ZN(new_n984));
  AOI21_X1  g559(.A(G37), .B1(new_n984), .B2(new_n929), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n985), .A2(KEYINPUT109), .A3(new_n968), .A4(new_n967), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n972), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n985), .A2(KEYINPUT43), .A3(new_n967), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT43), .B1(new_n985), .B2(new_n981), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT44), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n989), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n990), .B1(new_n989), .B2(new_n993), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(G397));
  NAND3_X1  g571(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n998));
  INV_X1    g573(.A(G8), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n998), .B1(G166), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n891), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n891), .A2(KEYINPUT45), .A3(new_n1003), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1006), .A2(new_n1007), .A3(G160), .A4(G40), .ZN(new_n1008));
  INV_X1    g583(.A(G1971), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G40), .ZN(new_n1011));
  AOI211_X1 g586(.A(new_n1011), .B(new_n477), .C1(new_n488), .C2(G2105), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n891), .A2(new_n1013), .A3(new_n1003), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(new_n891), .B2(new_n1003), .ZN(new_n1016));
  NOR3_X1   g591(.A1(G164), .A2(KEYINPUT115), .A3(G1384), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1012), .B(new_n1014), .C1(new_n1018), .C2(new_n1013), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1010), .B1(new_n1019), .B2(G2090), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1020), .A2(KEYINPUT118), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT116), .B(G8), .Z(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n1020), .B2(KEYINPUT118), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1002), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT115), .B1(G164), .B2(G1384), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n891), .A2(new_n1015), .A3(new_n1003), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(new_n1027), .A3(new_n1013), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1004), .A2(KEYINPUT50), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(new_n1012), .A3(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1010), .B1(G2090), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G8), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(new_n1002), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1018), .A2(new_n1012), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n817), .A2(G1976), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(new_n1023), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT52), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n546), .A2(G86), .ZN(new_n1038));
  OAI21_X1  g613(.A(G1981), .B1(new_n810), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(G305), .B2(G1981), .ZN(new_n1040));
  NOR2_X1   g615(.A1(KEYINPUT117), .A2(KEYINPUT49), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI221_X1 g617(.A(new_n1039), .B1(KEYINPUT117), .B2(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1042), .A2(new_n1043), .A3(new_n1023), .A4(new_n1034), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n817), .B2(G1976), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1037), .B(new_n1044), .C1(new_n1036), .C2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1033), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1049), .B(new_n1012), .C1(new_n1018), .C2(KEYINPUT45), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT45), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G160), .A2(G40), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT119), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(G2078), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1050), .A2(new_n1053), .A3(new_n1007), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G2078), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1012), .A2(new_n1057), .A3(new_n1007), .A4(new_n1006), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1054), .A2(new_n1058), .B1(new_n1030), .B2(new_n745), .ZN(new_n1059));
  AOI21_X1  g634(.A(G301), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1025), .A2(new_n1048), .A3(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1030), .A2(G2084), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1050), .A2(new_n1053), .A3(new_n1007), .ZN(new_n1063));
  INV_X1    g638(.A(G1966), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(G168), .A2(new_n1022), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1067), .B1(new_n1065), .B2(new_n999), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT51), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1066), .A2(KEYINPUT51), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1065), .B2(new_n1022), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1068), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT62), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1061), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1065), .A2(new_n1022), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1077), .A2(new_n1071), .B1(new_n1069), .B2(KEYINPUT51), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1078), .A2(KEYINPUT62), .A3(new_n1068), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT126), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1033), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1034), .A2(new_n1023), .ZN(new_n1082));
  NOR2_X1   g657(.A1(G305), .A2(G1981), .ZN(new_n1083));
  NOR2_X1   g658(.A1(G288), .A2(G1976), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1083), .B1(new_n1044), .B2(new_n1084), .ZN(new_n1085));
  OAI22_X1  g660(.A1(new_n1081), .A2(new_n1047), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1348), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1030), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G2067), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1018), .A2(new_n1012), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(KEYINPUT60), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT124), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1088), .A2(new_n1093), .A3(KEYINPUT60), .A4(new_n1090), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n634), .A3(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1096), .A2(KEYINPUT60), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1091), .A2(KEYINPUT124), .A3(new_n645), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1008), .A2(G1996), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT58), .B(G1341), .Z(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n1018), .B2(new_n1012), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n563), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT59), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(new_n1105), .A3(KEYINPUT59), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1956), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1013), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1112));
  NAND3_X1  g687(.A1(G160), .A2(G40), .A3(new_n1014), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT56), .B(G2072), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT122), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1012), .A2(new_n1007), .A3(new_n1006), .A4(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n584), .A2(new_n586), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1120), .B2(KEYINPUT121), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(G299), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n638), .B(new_n1121), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1123), .A2(new_n1125), .A3(KEYINPUT61), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT61), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1099), .A2(new_n1110), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1123), .B1(new_n1096), .B2(new_n645), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1125), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1058), .A2(new_n1054), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1059), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(G171), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1132), .B1(new_n1135), .B2(new_n1060), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT125), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1138), .B(new_n1132), .C1(new_n1135), .C2(new_n1060), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1129), .A2(new_n1131), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1134), .A2(G171), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1056), .A2(new_n1059), .A3(G301), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1141), .A2(KEYINPUT54), .A3(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1025), .A2(new_n1143), .A3(new_n1048), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1073), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1086), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT62), .B1(new_n1078), .B2(new_n1068), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1061), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1076), .A2(G168), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT120), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1076), .A2(new_n1153), .A3(G168), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1032), .A2(new_n1002), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1048), .A2(KEYINPUT63), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1025), .A2(new_n1048), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1158), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1159));
  OAI22_X1  g734(.A1(new_n1155), .A2(new_n1157), .B1(new_n1159), .B2(KEYINPUT63), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1080), .A2(new_n1146), .A3(new_n1150), .A4(new_n1160), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n792), .A2(new_n1089), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n792), .A2(new_n1089), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT113), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1052), .A2(new_n1006), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT114), .ZN(new_n1168));
  INV_X1    g743(.A(new_n772), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1166), .A2(new_n1169), .A3(G1996), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1052), .A2(new_n1006), .A3(G1996), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1171), .B(KEYINPUT112), .Z(new_n1172));
  OAI211_X1 g747(.A(new_n1168), .B(new_n1170), .C1(new_n1169), .C2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n847), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n844), .B(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1173), .B1(new_n1166), .B2(new_n1175), .ZN(new_n1176));
  OR3_X1    g751(.A1(new_n833), .A2(KEYINPUT111), .A3(new_n836), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n833), .A2(new_n836), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT111), .B1(new_n833), .B2(new_n836), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1177), .B(new_n1166), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1176), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1161), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n844), .A2(new_n1174), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1163), .B1(new_n1173), .B2(new_n1184), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1185), .A2(new_n1166), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1166), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1172), .A2(KEYINPUT46), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1172), .A2(KEYINPUT46), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g765(.A(new_n1190), .B(KEYINPUT47), .Z(new_n1191));
  NAND2_X1  g766(.A1(new_n1179), .A2(new_n1166), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT48), .ZN(new_n1193));
  AOI211_X1 g768(.A(new_n1186), .B(new_n1191), .C1(new_n1176), .C2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1183), .A2(new_n1194), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g770(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1197));
  XOR2_X1   g771(.A(new_n1197), .B(KEYINPUT127), .Z(new_n1198));
  NOR2_X1   g772(.A1(G229), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g773(.A1(new_n898), .A2(new_n987), .A3(new_n1199), .ZN(G225));
  INV_X1    g774(.A(G225), .ZN(G308));
endmodule


