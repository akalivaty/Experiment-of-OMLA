

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745;

  NOR2_X2 U368 ( .A1(n650), .A2(n723), .ZN(n693) );
  OR2_X1 U369 ( .A1(n566), .A2(n557), .ZN(n364) );
  XNOR2_X1 U370 ( .A(n423), .B(G146), .ZN(n537) );
  INV_X1 U371 ( .A(G125), .ZN(n423) );
  XNOR2_X1 U372 ( .A(n529), .B(KEYINPUT76), .ZN(n553) );
  AND2_X2 U373 ( .A1(n689), .A2(n366), .ZN(n582) );
  XNOR2_X2 U374 ( .A(n732), .B(n482), .ZN(n527) );
  XNOR2_X2 U375 ( .A(n534), .B(n405), .ZN(n732) );
  INV_X1 U376 ( .A(n580), .ZN(n666) );
  INV_X4 U377 ( .A(G116), .ZN(n453) );
  INV_X2 U378 ( .A(G131), .ZN(n436) );
  NOR2_X1 U379 ( .A1(n666), .A2(n556), .ZN(n647) );
  XNOR2_X1 U380 ( .A(n401), .B(n400), .ZN(n554) );
  XNOR2_X1 U381 ( .A(n603), .B(n434), .ZN(n580) );
  XNOR2_X1 U382 ( .A(n528), .B(G472), .ZN(n675) );
  OR2_X1 U383 ( .A1(n706), .A2(G902), .ZN(n419) );
  XOR2_X1 U384 ( .A(n706), .B(n705), .Z(n708) );
  XNOR2_X1 U385 ( .A(n440), .B(n478), .ZN(n551) );
  OR2_X1 U386 ( .A1(n618), .A2(G902), .ZN(n440) );
  XNOR2_X1 U387 ( .A(n618), .B(n459), .ZN(n619) );
  XNOR2_X1 U388 ( .A(n386), .B(n476), .ZN(n618) );
  XNOR2_X1 U389 ( .A(n456), .B(n521), .ZN(n533) );
  XNOR2_X1 U390 ( .A(n532), .B(KEYINPUT16), .ZN(n451) );
  XNOR2_X1 U391 ( .A(G902), .B(KEYINPUT15), .ZN(n611) );
  AND2_X1 U392 ( .A1(n613), .A2(n433), .ZN(n395) );
  BUF_X2 U393 ( .A(n675), .Z(n345) );
  XNOR2_X1 U394 ( .A(n610), .B(KEYINPUT45), .ZN(n613) );
  XNOR2_X2 U395 ( .A(n375), .B(n369), .ZN(n366) );
  BUF_X1 U396 ( .A(n745), .Z(n346) );
  XNOR2_X1 U397 ( .A(n371), .B(n543), .ZN(n745) );
  XNOR2_X2 U398 ( .A(n541), .B(n380), .ZN(n378) );
  INV_X1 U399 ( .A(KEYINPUT48), .ZN(n410) );
  NOR2_X1 U400 ( .A1(n438), .A2(n611), .ZN(n433) );
  INV_X1 U401 ( .A(n651), .ZN(n438) );
  XNOR2_X1 U402 ( .A(n481), .B(n406), .ZN(n405) );
  XNOR2_X1 U403 ( .A(n435), .B(G134), .ZN(n406) );
  INV_X1 U404 ( .A(KEYINPUT67), .ZN(n435) );
  INV_X1 U405 ( .A(KEYINPUT6), .ZN(n367) );
  INV_X1 U406 ( .A(G146), .ZN(n482) );
  INV_X1 U407 ( .A(KEYINPUT1), .ZN(n434) );
  INV_X1 U408 ( .A(KEYINPUT107), .ZN(n448) );
  INV_X1 U409 ( .A(KEYINPUT44), .ZN(n429) );
  XNOR2_X1 U410 ( .A(KEYINPUT38), .B(KEYINPUT74), .ZN(n394) );
  XNOR2_X1 U411 ( .A(n494), .B(KEYINPUT20), .ZN(n503) );
  XNOR2_X1 U412 ( .A(G116), .B(KEYINPUT101), .ZN(n522) );
  XOR2_X1 U413 ( .A(G137), .B(KEYINPUT5), .Z(n523) );
  XNOR2_X1 U414 ( .A(n520), .B(n457), .ZN(n456) );
  INV_X1 U415 ( .A(KEYINPUT3), .ZN(n457) );
  INV_X1 U416 ( .A(KEYINPUT86), .ZN(n407) );
  INV_X1 U417 ( .A(n649), .ZN(n409) );
  INV_X1 U418 ( .A(n656), .ZN(n416) );
  INV_X1 U419 ( .A(KEYINPUT39), .ZN(n415) );
  XNOR2_X1 U420 ( .A(G128), .B(G119), .ZN(n507) );
  XNOR2_X1 U421 ( .A(G110), .B(KEYINPUT23), .ZN(n508) );
  XOR2_X1 U422 ( .A(KEYINPUT95), .B(KEYINPUT24), .Z(n509) );
  XOR2_X1 U423 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n469) );
  XNOR2_X1 U424 ( .A(n506), .B(n353), .ZN(n731) );
  XNOR2_X1 U425 ( .A(G134), .B(G122), .ZN(n463) );
  XOR2_X1 U426 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n464) );
  XOR2_X1 U427 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n466) );
  NOR2_X1 U428 ( .A1(G953), .A2(G237), .ZN(n525) );
  XNOR2_X1 U429 ( .A(n537), .B(n439), .ZN(n506) );
  XNOR2_X1 U430 ( .A(KEYINPUT10), .B(G140), .ZN(n439) );
  XNOR2_X1 U431 ( .A(n487), .B(n390), .ZN(n389) );
  XNOR2_X1 U432 ( .A(n486), .B(n485), .ZN(n487) );
  INV_X1 U433 ( .A(KEYINPUT94), .ZN(n485) );
  XNOR2_X1 U434 ( .A(G101), .B(G140), .ZN(n483) );
  INV_X1 U435 ( .A(KEYINPUT4), .ZN(n479) );
  XNOR2_X1 U436 ( .A(KEYINPUT79), .B(KEYINPUT78), .ZN(n535) );
  AND2_X1 U437 ( .A1(G224), .A2(n734), .ZN(n461) );
  XNOR2_X1 U438 ( .A(n365), .B(n425), .ZN(n566) );
  INV_X1 U439 ( .A(KEYINPUT110), .ZN(n425) );
  NOR2_X1 U440 ( .A1(n348), .A2(n639), .ZN(n365) );
  NOR2_X1 U441 ( .A1(n596), .A2(n666), .ZN(n588) );
  XNOR2_X1 U442 ( .A(n398), .B(KEYINPUT28), .ZN(n546) );
  NAND2_X1 U443 ( .A1(n399), .A2(n445), .ZN(n398) );
  INV_X1 U444 ( .A(n554), .ZN(n399) );
  NOR2_X1 U445 ( .A1(n449), .A2(n448), .ZN(n447) );
  INV_X1 U446 ( .A(n666), .ZN(n449) );
  NOR2_X1 U447 ( .A1(n446), .A2(n445), .ZN(n444) );
  NOR2_X1 U448 ( .A1(n666), .A2(KEYINPUT107), .ZN(n446) );
  XOR2_X1 U449 ( .A(n472), .B(n471), .Z(n560) );
  NOR2_X1 U450 ( .A1(n711), .A2(G902), .ZN(n471) );
  XNOR2_X1 U451 ( .A(KEYINPUT72), .B(G101), .ZN(n520) );
  INV_X1 U452 ( .A(KEYINPUT75), .ZN(n393) );
  NAND2_X1 U453 ( .A1(n609), .A2(n608), .ZN(n610) );
  OR2_X1 U454 ( .A1(G237), .A2(G902), .ZN(n542) );
  OR2_X2 U455 ( .A1(n656), .A2(n657), .ZN(n379) );
  NOR2_X1 U456 ( .A1(n587), .A2(n657), .ZN(n417) );
  INV_X1 U457 ( .A(KEYINPUT68), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n495), .B(n403), .ZN(n402) );
  NAND2_X1 U459 ( .A1(n503), .A2(G221), .ZN(n404) );
  INV_X1 U460 ( .A(KEYINPUT98), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n533), .B(n458), .ZN(n526) );
  XNOR2_X1 U462 ( .A(n524), .B(n355), .ZN(n458) );
  INV_X1 U463 ( .A(KEYINPUT85), .ZN(n427) );
  BUF_X1 U464 ( .A(n613), .Z(n652) );
  NOR2_X1 U465 ( .A1(n416), .A2(n415), .ZN(n414) );
  INV_X1 U466 ( .A(KEYINPUT0), .ZN(n369) );
  AND2_X1 U467 ( .A1(n596), .A2(n664), .ZN(n579) );
  AND2_X1 U468 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U469 ( .A(n557), .B(KEYINPUT19), .ZN(n577) );
  XNOR2_X1 U470 ( .A(n551), .B(n384), .ZN(n559) );
  INV_X1 U471 ( .A(KEYINPUT102), .ZN(n384) );
  XNOR2_X1 U472 ( .A(n363), .B(n731), .ZN(n717) );
  XNOR2_X1 U473 ( .A(n377), .B(n376), .ZN(n711) );
  XNOR2_X1 U474 ( .A(n420), .B(n465), .ZN(n376) );
  XNOR2_X1 U475 ( .A(n470), .B(n467), .ZN(n377) );
  XNOR2_X1 U476 ( .A(n350), .B(n506), .ZN(n386) );
  XNOR2_X1 U477 ( .A(n389), .B(n488), .ZN(n490) );
  NOR2_X1 U478 ( .A1(G952), .A2(n734), .ZN(n719) );
  XNOR2_X1 U479 ( .A(n549), .B(n548), .ZN(n743) );
  XNOR2_X1 U480 ( .A(n364), .B(KEYINPUT36), .ZN(n556) );
  XNOR2_X1 U481 ( .A(n594), .B(n593), .ZN(n381) );
  AND2_X1 U482 ( .A1(n441), .A2(n599), .ZN(n392) );
  AND2_X1 U483 ( .A1(n422), .A2(n444), .ZN(n443) );
  AND2_X1 U484 ( .A1(n560), .A2(n551), .ZN(n347) );
  OR2_X1 U485 ( .A1(n555), .A2(n554), .ZN(n348) );
  NOR2_X1 U486 ( .A1(n605), .A2(n368), .ZN(n349) );
  XOR2_X1 U487 ( .A(n481), .B(n477), .Z(n350) );
  XNOR2_X1 U488 ( .A(n362), .B(n513), .ZN(n670) );
  XOR2_X1 U489 ( .A(n507), .B(KEYINPUT96), .Z(n351) );
  AND2_X1 U490 ( .A1(G210), .A2(n542), .ZN(n352) );
  XNOR2_X1 U491 ( .A(G137), .B(KEYINPUT66), .ZN(n353) );
  XNOR2_X1 U492 ( .A(n404), .B(n402), .ZN(n671) );
  XOR2_X1 U493 ( .A(n493), .B(n492), .Z(n354) );
  AND2_X1 U494 ( .A1(n525), .A2(G210), .ZN(n355) );
  NAND2_X1 U495 ( .A1(n416), .A2(n415), .ZN(n356) );
  NOR2_X1 U496 ( .A1(n586), .A2(n599), .ZN(n664) );
  AND2_X1 U497 ( .A1(n347), .A2(n671), .ZN(n357) );
  XOR2_X1 U498 ( .A(KEYINPUT22), .B(KEYINPUT73), .Z(n358) );
  XOR2_X1 U499 ( .A(n623), .B(KEYINPUT62), .Z(n359) );
  AND2_X1 U500 ( .A1(n617), .A2(n616), .ZN(n360) );
  AND2_X2 U501 ( .A1(n617), .A2(n616), .ZN(n715) );
  NAND2_X1 U502 ( .A1(n361), .A2(n347), .ZN(n547) );
  XNOR2_X2 U503 ( .A(n379), .B(KEYINPUT111), .ZN(n361) );
  NAND2_X1 U504 ( .A1(n361), .A2(n660), .ZN(n661) );
  NOR2_X1 U505 ( .A1(n717), .A2(G902), .ZN(n362) );
  XNOR2_X1 U506 ( .A(n391), .B(n512), .ZN(n363) );
  AND2_X1 U507 ( .A1(n664), .A2(n366), .ZN(n601) );
  AND2_X2 U508 ( .A1(n366), .A2(n357), .ZN(n382) );
  XNOR2_X1 U509 ( .A(n675), .B(KEYINPUT106), .ZN(n587) );
  XNOR2_X1 U510 ( .A(n345), .B(n367), .ZN(n555) );
  INV_X1 U511 ( .A(n345), .ZN(n368) );
  NAND2_X1 U512 ( .A1(n426), .A2(n612), .ZN(n617) );
  XNOR2_X1 U513 ( .A(n370), .B(n410), .ZN(n396) );
  NAND2_X1 U514 ( .A1(n397), .A2(n383), .ZN(n370) );
  NAND2_X1 U515 ( .A1(n374), .A2(n561), .ZN(n371) );
  NAND2_X1 U516 ( .A1(n378), .A2(n611), .ZN(n428) );
  NAND2_X1 U517 ( .A1(n372), .A2(n431), .ZN(n430) );
  XNOR2_X1 U518 ( .A(n432), .B(KEYINPUT88), .ZN(n372) );
  INV_X1 U519 ( .A(n555), .ZN(n596) );
  XNOR2_X2 U520 ( .A(n421), .B(n581), .ZN(n689) );
  NAND2_X1 U521 ( .A1(n373), .A2(n395), .ZN(n388) );
  NAND2_X1 U522 ( .A1(n373), .A2(n615), .ZN(n650) );
  AND2_X1 U523 ( .A1(n373), .A2(n651), .ZN(n733) );
  XNOR2_X2 U524 ( .A(n408), .B(n407), .ZN(n373) );
  NAND2_X1 U525 ( .A1(n374), .A2(n644), .ZN(n651) );
  NAND2_X1 U526 ( .A1(n412), .A2(n411), .ZN(n374) );
  NAND2_X1 U527 ( .A1(n577), .A2(n578), .ZN(n375) );
  XNOR2_X1 U528 ( .A(n378), .B(n460), .ZN(n700) );
  XNOR2_X2 U529 ( .A(n387), .B(n394), .ZN(n656) );
  NAND2_X1 U530 ( .A1(n380), .A2(n726), .ZN(n727) );
  XNOR2_X2 U531 ( .A(n450), .B(n533), .ZN(n380) );
  NOR2_X2 U532 ( .A1(n631), .A2(n381), .ZN(n432) );
  XNOR2_X1 U533 ( .A(n381), .B(n744), .ZN(G21) );
  XNOR2_X2 U534 ( .A(n382), .B(n358), .ZN(n590) );
  AND2_X1 U535 ( .A1(n564), .A2(n565), .ZN(n383) );
  INV_X1 U536 ( .A(n587), .ZN(n445) );
  XNOR2_X1 U537 ( .A(n417), .B(KEYINPUT30), .ZN(n385) );
  XNOR2_X1 U538 ( .A(n550), .B(KEYINPUT46), .ZN(n397) );
  XNOR2_X1 U539 ( .A(n527), .B(n526), .ZN(n623) );
  NAND2_X1 U540 ( .A1(n385), .A2(n418), .ZN(n529) );
  NOR2_X1 U541 ( .A1(n545), .A2(n670), .ZN(n401) );
  AND2_X2 U542 ( .A1(n443), .A2(n392), .ZN(n631) );
  BUF_X1 U543 ( .A(n571), .Z(n387) );
  XNOR2_X1 U544 ( .A(n388), .B(n427), .ZN(n426) );
  XOR2_X1 U545 ( .A(G107), .B(G104), .Z(n484) );
  INV_X1 U546 ( .A(n531), .ZN(n390) );
  XNOR2_X1 U547 ( .A(n510), .B(n351), .ZN(n391) );
  NAND2_X1 U548 ( .A1(n442), .A2(n448), .ZN(n441) );
  XNOR2_X1 U549 ( .A(n537), .B(n461), .ZN(n538) );
  XNOR2_X2 U550 ( .A(n393), .B(G110), .ZN(n531) );
  XNOR2_X2 U551 ( .A(n530), .B(n531), .ZN(n452) );
  XNOR2_X2 U552 ( .A(n453), .B(G107), .ZN(n530) );
  NAND2_X1 U553 ( .A1(n396), .A2(n409), .ZN(n408) );
  XNOR2_X2 U554 ( .A(n436), .B(KEYINPUT65), .ZN(n481) );
  XNOR2_X2 U555 ( .A(n480), .B(n479), .ZN(n534) );
  XNOR2_X2 U556 ( .A(n437), .B(G128), .ZN(n480) );
  NAND2_X1 U557 ( .A1(n553), .A2(KEYINPUT39), .ZN(n411) );
  NOR2_X1 U558 ( .A1(n413), .A2(n414), .ZN(n412) );
  NOR2_X1 U559 ( .A1(n553), .A2(n356), .ZN(n413) );
  NAND2_X1 U560 ( .A1(n519), .A2(n518), .ZN(n418) );
  XNOR2_X2 U561 ( .A(n419), .B(n354), .ZN(n603) );
  XNOR2_X1 U562 ( .A(n707), .B(n708), .ZN(n709) );
  INV_X2 U563 ( .A(G143), .ZN(n437) );
  XNOR2_X2 U564 ( .A(n547), .B(KEYINPUT41), .ZN(n688) );
  XNOR2_X1 U565 ( .A(n530), .B(n466), .ZN(n420) );
  NAND2_X1 U566 ( .A1(n579), .A2(n580), .ZN(n421) );
  XNOR2_X2 U567 ( .A(n585), .B(KEYINPUT35), .ZN(n742) );
  XNOR2_X1 U568 ( .A(n430), .B(n429), .ZN(n609) );
  NAND2_X1 U569 ( .A1(n590), .A2(n447), .ZN(n422) );
  NAND2_X1 U570 ( .A1(n715), .A2(G475), .ZN(n620) );
  NOR2_X2 U571 ( .A1(n621), .A2(n719), .ZN(n622) );
  NOR2_X2 U572 ( .A1(n709), .A2(n719), .ZN(n710) );
  XNOR2_X1 U573 ( .A(n424), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U574 ( .A1(n702), .A2(n719), .ZN(n424) );
  NAND2_X1 U575 ( .A1(n715), .A2(G210), .ZN(n701) );
  NAND2_X2 U576 ( .A1(n571), .A2(n567), .ZN(n557) );
  XNOR2_X2 U577 ( .A(n428), .B(n352), .ZN(n571) );
  INV_X1 U578 ( .A(n742), .ZN(n431) );
  XNOR2_X2 U579 ( .A(G122), .B(G104), .ZN(n532) );
  INV_X1 U580 ( .A(n639), .ZN(n641) );
  NAND2_X1 U581 ( .A1(n590), .A2(n666), .ZN(n595) );
  INV_X1 U582 ( .A(n590), .ZN(n442) );
  XNOR2_X2 U583 ( .A(n452), .B(n451), .ZN(n450) );
  XNOR2_X1 U584 ( .A(n454), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U585 ( .A1(n455), .A2(n625), .ZN(n454) );
  XNOR2_X1 U586 ( .A(n624), .B(n359), .ZN(n455) );
  XNOR2_X1 U587 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U588 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U589 ( .A(KEYINPUT59), .B(KEYINPUT89), .ZN(n459) );
  XNOR2_X1 U590 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n460) );
  AND2_X1 U591 ( .A1(G214), .A2(n525), .ZN(n462) );
  XNOR2_X1 U592 ( .A(n475), .B(n462), .ZN(n476) );
  XNOR2_X1 U593 ( .A(KEYINPUT108), .B(KEYINPUT33), .ZN(n581) );
  XNOR2_X1 U594 ( .A(n538), .B(n539), .ZN(n540) );
  INV_X1 U595 ( .A(G469), .ZN(n492) );
  INV_X1 U596 ( .A(n693), .ZN(n616) );
  INV_X1 U597 ( .A(n719), .ZN(n625) );
  XNOR2_X1 U598 ( .A(KEYINPUT105), .B(G478), .ZN(n472) );
  XNOR2_X1 U599 ( .A(n464), .B(n463), .ZN(n467) );
  INV_X1 U600 ( .A(n480), .ZN(n465) );
  INV_X2 U601 ( .A(G953), .ZN(n734) );
  NAND2_X1 U602 ( .A1(G234), .A2(n734), .ZN(n468) );
  XNOR2_X1 U603 ( .A(n469), .B(n468), .ZN(n511) );
  NAND2_X1 U604 ( .A1(G217), .A2(n511), .ZN(n470) );
  XOR2_X1 U605 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n474) );
  XNOR2_X1 U606 ( .A(G143), .B(G113), .ZN(n473) );
  XNOR2_X1 U607 ( .A(n474), .B(n473), .ZN(n475) );
  INV_X1 U608 ( .A(n532), .ZN(n477) );
  XNOR2_X1 U609 ( .A(KEYINPUT13), .B(G475), .ZN(n478) );
  XNOR2_X1 U610 ( .A(n484), .B(n483), .ZN(n488) );
  NAND2_X1 U611 ( .A1(G227), .A2(n734), .ZN(n486) );
  INV_X1 U612 ( .A(n353), .ZN(n489) );
  XNOR2_X1 U613 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U614 ( .A(n527), .B(n491), .ZN(n706) );
  XNOR2_X1 U615 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n493) );
  XOR2_X1 U616 ( .A(KEYINPUT99), .B(KEYINPUT21), .Z(n495) );
  NAND2_X1 U617 ( .A1(n611), .A2(G234), .ZN(n494) );
  NAND2_X1 U618 ( .A1(G234), .A2(G237), .ZN(n496) );
  XNOR2_X1 U619 ( .A(n496), .B(KEYINPUT14), .ZN(n498) );
  NAND2_X1 U620 ( .A1(G952), .A2(n498), .ZN(n687) );
  NOR2_X1 U621 ( .A1(n687), .A2(G953), .ZN(n497) );
  XOR2_X1 U622 ( .A(n497), .B(KEYINPUT90), .Z(n572) );
  NAND2_X1 U623 ( .A1(n498), .A2(G902), .ZN(n499) );
  XNOR2_X1 U624 ( .A(n499), .B(KEYINPUT92), .ZN(n573) );
  NOR2_X1 U625 ( .A1(n573), .A2(G900), .ZN(n500) );
  NAND2_X1 U626 ( .A1(G953), .A2(n500), .ZN(n501) );
  NAND2_X1 U627 ( .A1(n572), .A2(n501), .ZN(n502) );
  NAND2_X1 U628 ( .A1(n671), .A2(n502), .ZN(n544) );
  NOR2_X1 U629 ( .A1(n603), .A2(n544), .ZN(n517) );
  XOR2_X1 U630 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n505) );
  NAND2_X1 U631 ( .A1(n503), .A2(G217), .ZN(n504) );
  XNOR2_X1 U632 ( .A(n505), .B(n504), .ZN(n513) );
  XNOR2_X1 U633 ( .A(n509), .B(n508), .ZN(n510) );
  NAND2_X1 U634 ( .A1(G221), .A2(n511), .ZN(n512) );
  NAND2_X1 U635 ( .A1(n517), .A2(n670), .ZN(n514) );
  NAND2_X1 U636 ( .A1(n514), .A2(KEYINPUT77), .ZN(n519) );
  INV_X1 U637 ( .A(KEYINPUT77), .ZN(n515) );
  AND2_X1 U638 ( .A1(n670), .A2(n515), .ZN(n516) );
  NAND2_X1 U639 ( .A1(n517), .A2(n516), .ZN(n518) );
  NAND2_X1 U640 ( .A1(G214), .A2(n542), .ZN(n567) );
  INV_X1 U641 ( .A(n567), .ZN(n657) );
  XOR2_X1 U642 ( .A(G119), .B(G113), .Z(n521) );
  XNOR2_X1 U643 ( .A(n523), .B(n522), .ZN(n524) );
  NOR2_X1 U644 ( .A1(n623), .A2(G902), .ZN(n528) );
  XOR2_X1 U645 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n536) );
  XNOR2_X1 U646 ( .A(n536), .B(n535), .ZN(n539) );
  XNOR2_X1 U647 ( .A(n534), .B(n540), .ZN(n541) );
  INV_X1 U648 ( .A(KEYINPUT40), .ZN(n543) );
  XOR2_X1 U649 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n549) );
  XOR2_X1 U650 ( .A(n544), .B(KEYINPUT69), .Z(n545) );
  NOR2_X1 U651 ( .A1(n603), .A2(n546), .ZN(n558) );
  NAND2_X1 U652 ( .A1(n558), .A2(n688), .ZN(n548) );
  NOR2_X2 U653 ( .A1(n745), .A2(n743), .ZN(n550) );
  NOR2_X1 U654 ( .A1(n560), .A2(n551), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n387), .A2(n583), .ZN(n552) );
  NOR2_X1 U656 ( .A1(n553), .A2(n552), .ZN(n637) );
  XNOR2_X1 U657 ( .A(KEYINPUT83), .B(n637), .ZN(n565) );
  XNOR2_X1 U658 ( .A(n561), .B(KEYINPUT109), .ZN(n639) );
  NAND2_X1 U659 ( .A1(n577), .A2(n558), .ZN(n638) );
  NOR2_X1 U660 ( .A1(n560), .A2(n559), .ZN(n644) );
  NOR2_X1 U661 ( .A1(n561), .A2(n644), .ZN(n659) );
  NOR2_X1 U662 ( .A1(n638), .A2(n659), .ZN(n562) );
  XOR2_X1 U663 ( .A(KEYINPUT47), .B(n562), .Z(n563) );
  NOR2_X1 U664 ( .A1(n647), .A2(n563), .ZN(n564) );
  NOR2_X1 U665 ( .A1(n580), .A2(n566), .ZN(n568) );
  NAND2_X1 U666 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U667 ( .A(KEYINPUT43), .B(n569), .Z(n570) );
  NOR2_X1 U668 ( .A1(n387), .A2(n570), .ZN(n649) );
  INV_X1 U669 ( .A(n572), .ZN(n575) );
  XNOR2_X1 U670 ( .A(G898), .B(KEYINPUT91), .ZN(n722) );
  NAND2_X1 U671 ( .A1(G953), .A2(n722), .ZN(n726) );
  NOR2_X1 U672 ( .A1(n573), .A2(n726), .ZN(n574) );
  NOR2_X1 U673 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U674 ( .A(KEYINPUT93), .B(n576), .ZN(n578) );
  INV_X1 U675 ( .A(n671), .ZN(n586) );
  INV_X1 U676 ( .A(n670), .ZN(n599) );
  XNOR2_X1 U677 ( .A(n582), .B(KEYINPUT34), .ZN(n584) );
  NAND2_X1 U678 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U679 ( .A1(n599), .A2(n588), .ZN(n589) );
  XNOR2_X1 U680 ( .A(n589), .B(KEYINPUT81), .ZN(n591) );
  NAND2_X1 U681 ( .A1(n591), .A2(n590), .ZN(n594) );
  XOR2_X1 U682 ( .A(KEYINPUT32), .B(KEYINPUT80), .Z(n592) );
  XNOR2_X1 U683 ( .A(KEYINPUT64), .B(n592), .ZN(n593) );
  NOR2_X1 U684 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U685 ( .A(n597), .B(KEYINPUT87), .ZN(n598) );
  NOR2_X1 U686 ( .A1(n599), .A2(n598), .ZN(n626) );
  NOR2_X1 U687 ( .A1(n345), .A2(n666), .ZN(n665) );
  INV_X1 U688 ( .A(n664), .ZN(n667) );
  NAND2_X1 U689 ( .A1(n665), .A2(n601), .ZN(n600) );
  XNOR2_X1 U690 ( .A(n600), .B(KEYINPUT31), .ZN(n645) );
  INV_X1 U691 ( .A(n601), .ZN(n602) );
  NOR2_X1 U692 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U693 ( .A(KEYINPUT100), .B(n604), .Z(n605) );
  NOR2_X1 U694 ( .A1(n645), .A2(n349), .ZN(n606) );
  NOR2_X1 U695 ( .A1(n659), .A2(n606), .ZN(n607) );
  NOR2_X1 U696 ( .A1(n626), .A2(n607), .ZN(n608) );
  INV_X1 U697 ( .A(KEYINPUT2), .ZN(n694) );
  OR2_X1 U698 ( .A1(n611), .A2(n694), .ZN(n612) );
  INV_X1 U699 ( .A(n652), .ZN(n723) );
  NAND2_X1 U700 ( .A1(KEYINPUT2), .A2(n651), .ZN(n614) );
  XOR2_X1 U701 ( .A(KEYINPUT82), .B(n614), .Z(n615) );
  XNOR2_X1 U702 ( .A(n622), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U703 ( .A1(n360), .A2(G472), .ZN(n624) );
  XOR2_X1 U704 ( .A(G101), .B(n626), .Z(G3) );
  NAND2_X1 U705 ( .A1(n641), .A2(n349), .ZN(n627) );
  XNOR2_X1 U706 ( .A(n627), .B(G104), .ZN(G6) );
  XOR2_X1 U707 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n629) );
  NAND2_X1 U708 ( .A1(n349), .A2(n644), .ZN(n628) );
  XNOR2_X1 U709 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U710 ( .A(G107), .B(n630), .ZN(G9) );
  XNOR2_X1 U711 ( .A(n631), .B(G110), .ZN(n632) );
  XNOR2_X1 U712 ( .A(n632), .B(KEYINPUT113), .ZN(G12) );
  INV_X1 U713 ( .A(n644), .ZN(n633) );
  NOR2_X1 U714 ( .A1(n633), .A2(n638), .ZN(n635) );
  XNOR2_X1 U715 ( .A(KEYINPUT29), .B(KEYINPUT114), .ZN(n634) );
  XNOR2_X1 U716 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U717 ( .A(G128), .B(n636), .ZN(G30) );
  XOR2_X1 U718 ( .A(n637), .B(G143), .Z(G45) );
  NOR2_X1 U719 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U720 ( .A(G146), .B(n640), .Z(G48) );
  XOR2_X1 U721 ( .A(G113), .B(KEYINPUT115), .Z(n643) );
  NAND2_X1 U722 ( .A1(n641), .A2(n645), .ZN(n642) );
  XNOR2_X1 U723 ( .A(n643), .B(n642), .ZN(G15) );
  NAND2_X1 U724 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U725 ( .A(n646), .B(G116), .ZN(G18) );
  XNOR2_X1 U726 ( .A(n647), .B(G125), .ZN(n648) );
  XNOR2_X1 U727 ( .A(n648), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U728 ( .A(G134), .B(n651), .ZN(G36) );
  XOR2_X1 U729 ( .A(G140), .B(n649), .Z(G42) );
  INV_X1 U730 ( .A(n650), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n652), .A2(n733), .ZN(n653) );
  NOR2_X1 U732 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U733 ( .A1(G953), .A2(n655), .ZN(n698) );
  NAND2_X1 U734 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U735 ( .A1(n658), .A2(n347), .ZN(n662) );
  INV_X1 U736 ( .A(n659), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U738 ( .A1(n689), .A2(n663), .ZN(n683) );
  NAND2_X1 U739 ( .A1(n665), .A2(n664), .ZN(n678) );
  XOR2_X1 U740 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n669) );
  NAND2_X1 U741 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U742 ( .A(n669), .B(n668), .ZN(n674) );
  NOR2_X1 U743 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U744 ( .A(KEYINPUT49), .B(n672), .Z(n673) );
  NOR2_X1 U745 ( .A1(n674), .A2(n673), .ZN(n676) );
  NAND2_X1 U746 ( .A1(n676), .A2(n345), .ZN(n677) );
  NAND2_X1 U747 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U748 ( .A(n679), .B(KEYINPUT51), .ZN(n680) );
  XNOR2_X1 U749 ( .A(n680), .B(KEYINPUT117), .ZN(n681) );
  NAND2_X1 U750 ( .A1(n681), .A2(n688), .ZN(n682) );
  NAND2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U752 ( .A(n684), .B(KEYINPUT52), .ZN(n685) );
  XOR2_X1 U753 ( .A(KEYINPUT118), .B(n685), .Z(n686) );
  NOR2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n691) );
  AND2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U757 ( .A(n692), .B(KEYINPUT119), .ZN(n696) );
  NOR2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U759 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U760 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U761 ( .A(KEYINPUT53), .B(n699), .Z(G75) );
  XOR2_X1 U762 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n704) );
  XNOR2_X1 U763 ( .A(KEYINPUT121), .B(KEYINPUT120), .ZN(n703) );
  XNOR2_X1 U764 ( .A(n704), .B(n703), .ZN(n705) );
  NAND2_X1 U765 ( .A1(n715), .A2(G469), .ZN(n707) );
  XNOR2_X1 U766 ( .A(n710), .B(KEYINPUT122), .ZN(G54) );
  XOR2_X1 U767 ( .A(n711), .B(KEYINPUT123), .Z(n713) );
  NAND2_X1 U768 ( .A1(n360), .A2(G478), .ZN(n712) );
  XNOR2_X1 U769 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U770 ( .A1(n719), .A2(n714), .ZN(G63) );
  NAND2_X1 U771 ( .A1(G217), .A2(n360), .ZN(n716) );
  XNOR2_X1 U772 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U773 ( .A1(n719), .A2(n718), .ZN(G66) );
  NAND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n720) );
  XOR2_X1 U775 ( .A(KEYINPUT61), .B(n720), .Z(n721) );
  NOR2_X1 U776 ( .A1(n722), .A2(n721), .ZN(n725) );
  NOR2_X1 U777 ( .A1(G953), .A2(n723), .ZN(n724) );
  NOR2_X1 U778 ( .A1(n725), .A2(n724), .ZN(n730) );
  XOR2_X1 U779 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n728) );
  XNOR2_X1 U780 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U781 ( .A(n730), .B(n729), .ZN(G69) );
  XNOR2_X1 U782 ( .A(n732), .B(n731), .ZN(n736) );
  XOR2_X1 U783 ( .A(n733), .B(n736), .Z(n735) );
  NAND2_X1 U784 ( .A1(n735), .A2(n734), .ZN(n740) );
  XNOR2_X1 U785 ( .A(G227), .B(n736), .ZN(n737) );
  NAND2_X1 U786 ( .A1(n737), .A2(G900), .ZN(n738) );
  NAND2_X1 U787 ( .A1(G953), .A2(n738), .ZN(n739) );
  NAND2_X1 U788 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U789 ( .A(KEYINPUT126), .B(n741), .ZN(G72) );
  XOR2_X1 U790 ( .A(n742), .B(G122), .Z(G24) );
  XOR2_X1 U791 ( .A(n743), .B(G137), .Z(G39) );
  XNOR2_X1 U792 ( .A(G119), .B(KEYINPUT127), .ZN(n744) );
  XOR2_X1 U793 ( .A(G131), .B(n346), .Z(G33) );
endmodule

