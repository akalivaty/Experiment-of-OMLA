

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U560 ( .A(G2104), .ZN(n592) );
  NOR2_X1 U561 ( .A1(n671), .A2(n968), .ZN(n616) );
  NOR2_X1 U562 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U563 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U564 ( .A1(G1966), .A2(n717), .ZN(n687) );
  OR2_X1 U565 ( .A1(n690), .A2(n689), .ZN(n691) );
  INV_X1 U566 ( .A(KEYINPUT103), .ZN(n693) );
  AND2_X1 U567 ( .A1(n606), .A2(n722), .ZN(n657) );
  INV_X1 U568 ( .A(n657), .ZN(n671) );
  NOR2_X1 U569 ( .A1(G164), .A2(G1384), .ZN(n605) );
  XNOR2_X1 U570 ( .A(n605), .B(KEYINPUT64), .ZN(n722) );
  INV_X1 U571 ( .A(G2105), .ZN(n591) );
  NOR2_X1 U572 ( .A1(n711), .A2(n710), .ZN(n720) );
  NAND2_X1 U573 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U574 ( .A1(n577), .A2(G651), .ZN(n810) );
  XNOR2_X1 U575 ( .A(n596), .B(KEYINPUT67), .ZN(n776) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n577) );
  INV_X1 U577 ( .A(G651), .ZN(n531) );
  NOR2_X1 U578 ( .A1(n577), .A2(n531), .ZN(n809) );
  NAND2_X1 U579 ( .A1(G73), .A2(n809), .ZN(n529) );
  XNOR2_X1 U580 ( .A(n529), .B(KEYINPUT82), .ZN(n530) );
  XNOR2_X1 U581 ( .A(n530), .B(KEYINPUT2), .ZN(n534) );
  NOR2_X1 U582 ( .A1(G543), .A2(n531), .ZN(n532) );
  XOR2_X1 U583 ( .A(KEYINPUT1), .B(n532), .Z(n805) );
  NAND2_X1 U584 ( .A1(G61), .A2(n805), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n538) );
  NOR2_X1 U586 ( .A1(G543), .A2(G651), .ZN(n806) );
  NAND2_X1 U587 ( .A1(G86), .A2(n806), .ZN(n536) );
  NAND2_X1 U588 ( .A1(G48), .A2(n810), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U590 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U591 ( .A(KEYINPUT83), .B(n539), .ZN(G305) );
  NAND2_X1 U592 ( .A1(G65), .A2(n805), .ZN(n541) );
  NAND2_X1 U593 ( .A1(G53), .A2(n810), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n541), .A2(n540), .ZN(n545) );
  NAND2_X1 U595 ( .A1(G91), .A2(n806), .ZN(n543) );
  NAND2_X1 U596 ( .A1(G78), .A2(n809), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n544) );
  OR2_X1 U598 ( .A1(n545), .A2(n544), .ZN(G299) );
  NAND2_X1 U599 ( .A1(G64), .A2(n805), .ZN(n547) );
  NAND2_X1 U600 ( .A1(G52), .A2(n810), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n552) );
  NAND2_X1 U602 ( .A1(G90), .A2(n806), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G77), .A2(n809), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U605 ( .A(KEYINPUT9), .B(n550), .Z(n551) );
  NOR2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U607 ( .A(KEYINPUT69), .B(n553), .Z(G171) );
  XNOR2_X1 U608 ( .A(KEYINPUT6), .B(KEYINPUT78), .ZN(n557) );
  NAND2_X1 U609 ( .A1(G63), .A2(n805), .ZN(n555) );
  NAND2_X1 U610 ( .A1(G51), .A2(n810), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U612 ( .A(n557), .B(n556), .ZN(n564) );
  NAND2_X1 U613 ( .A1(n806), .A2(G89), .ZN(n558) );
  XNOR2_X1 U614 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G76), .A2(n809), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U617 ( .A(KEYINPUT77), .B(n561), .ZN(n562) );
  XNOR2_X1 U618 ( .A(KEYINPUT5), .B(n562), .ZN(n563) );
  NOR2_X1 U619 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U620 ( .A(KEYINPUT7), .B(n565), .Z(G168) );
  NAND2_X1 U621 ( .A1(G88), .A2(n806), .ZN(n567) );
  NAND2_X1 U622 ( .A1(G75), .A2(n809), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n567), .A2(n566), .ZN(n572) );
  NAND2_X1 U624 ( .A1(G50), .A2(n810), .ZN(n568) );
  XNOR2_X1 U625 ( .A(n568), .B(KEYINPUT84), .ZN(n570) );
  NAND2_X1 U626 ( .A1(n805), .A2(G62), .ZN(n569) );
  NAND2_X1 U627 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U628 ( .A1(n572), .A2(n571), .ZN(G166) );
  INV_X1 U629 ( .A(G166), .ZN(G303) );
  XOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U631 ( .A1(G49), .A2(n810), .ZN(n574) );
  NAND2_X1 U632 ( .A1(G74), .A2(G651), .ZN(n573) );
  NAND2_X1 U633 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U634 ( .A1(n805), .A2(n575), .ZN(n576) );
  XOR2_X1 U635 ( .A(KEYINPUT81), .B(n576), .Z(n579) );
  NAND2_X1 U636 ( .A1(n577), .A2(G87), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n579), .A2(n578), .ZN(G288) );
  NAND2_X1 U638 ( .A1(G85), .A2(n806), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G72), .A2(n809), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U641 ( .A1(G60), .A2(n805), .ZN(n583) );
  NAND2_X1 U642 ( .A1(G47), .A2(n810), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U644 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U645 ( .A(KEYINPUT68), .B(n586), .Z(G290) );
  NOR2_X1 U646 ( .A1(G2104), .A2(n591), .ZN(n598) );
  BUF_X1 U647 ( .A(n598), .Z(n892) );
  NAND2_X1 U648 ( .A1(G125), .A2(n892), .ZN(n587) );
  XNOR2_X1 U649 ( .A(n587), .B(KEYINPUT66), .ZN(n590) );
  AND2_X1 U650 ( .A1(n591), .A2(G2104), .ZN(n887) );
  NAND2_X1 U651 ( .A1(G101), .A2(n887), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT23), .B(n588), .Z(n589) );
  AND2_X1 U653 ( .A1(n590), .A2(n589), .ZN(n775) );
  AND2_X1 U654 ( .A1(G40), .A2(n775), .ZN(n597) );
  XNOR2_X2 U655 ( .A(n593), .B(KEYINPUT17), .ZN(n886) );
  NAND2_X1 U656 ( .A1(n886), .A2(G137), .ZN(n595) );
  AND2_X1 U657 ( .A1(G2104), .A2(G2105), .ZN(n890) );
  NAND2_X1 U658 ( .A1(n890), .A2(G113), .ZN(n594) );
  NAND2_X1 U659 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n597), .A2(n776), .ZN(n721) );
  INV_X1 U661 ( .A(n721), .ZN(n606) );
  NAND2_X1 U662 ( .A1(n886), .A2(G138), .ZN(n604) );
  NAND2_X1 U663 ( .A1(G114), .A2(n890), .ZN(n600) );
  NAND2_X1 U664 ( .A1(G126), .A2(n598), .ZN(n599) );
  AND2_X1 U665 ( .A1(n600), .A2(n599), .ZN(n602) );
  NAND2_X1 U666 ( .A1(G102), .A2(n887), .ZN(n601) );
  AND2_X1 U667 ( .A1(n602), .A2(n601), .ZN(n603) );
  AND2_X1 U668 ( .A1(n604), .A2(n603), .ZN(G164) );
  NAND2_X1 U669 ( .A1(G8), .A2(n671), .ZN(n607) );
  XOR2_X2 U670 ( .A(KEYINPUT97), .B(n607), .Z(n717) );
  NOR2_X1 U671 ( .A1(G1981), .A2(G305), .ZN(n608) );
  XOR2_X1 U672 ( .A(n608), .B(KEYINPUT24), .Z(n609) );
  NOR2_X1 U673 ( .A1(n717), .A2(n609), .ZN(n711) );
  XNOR2_X1 U674 ( .A(n657), .B(KEYINPUT99), .ZN(n641) );
  INV_X1 U675 ( .A(G2072), .ZN(n951) );
  NOR2_X1 U676 ( .A1(n641), .A2(n951), .ZN(n611) );
  XNOR2_X1 U677 ( .A(KEYINPUT27), .B(KEYINPUT100), .ZN(n610) );
  XNOR2_X1 U678 ( .A(n611), .B(n610), .ZN(n613) );
  NAND2_X1 U679 ( .A1(n641), .A2(G1956), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U681 ( .A(n614), .B(KEYINPUT101), .Z(n652) );
  OR2_X1 U682 ( .A1(G299), .A2(n652), .ZN(n650) );
  INV_X1 U683 ( .A(G1996), .ZN(n968) );
  INV_X1 U684 ( .A(KEYINPUT26), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n616), .B(n615), .ZN(n629) );
  AND2_X1 U686 ( .A1(n671), .A2(G1341), .ZN(n627) );
  XOR2_X1 U687 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n618) );
  NAND2_X1 U688 ( .A1(G56), .A2(n805), .ZN(n617) );
  XNOR2_X1 U689 ( .A(n618), .B(n617), .ZN(n624) );
  NAND2_X1 U690 ( .A1(n806), .A2(G81), .ZN(n619) );
  XNOR2_X1 U691 ( .A(n619), .B(KEYINPUT12), .ZN(n621) );
  NAND2_X1 U692 ( .A1(G68), .A2(n809), .ZN(n620) );
  NAND2_X1 U693 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U694 ( .A(KEYINPUT13), .B(n622), .Z(n623) );
  NOR2_X1 U695 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n810), .A2(G43), .ZN(n625) );
  NAND2_X1 U697 ( .A1(n626), .A2(n625), .ZN(n997) );
  NOR2_X1 U698 ( .A1(n627), .A2(n997), .ZN(n628) );
  AND2_X1 U699 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U700 ( .A(KEYINPUT65), .B(n630), .ZN(n646) );
  XNOR2_X1 U701 ( .A(KEYINPUT76), .B(KEYINPUT15), .ZN(n640) );
  NAND2_X1 U702 ( .A1(G92), .A2(n806), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n631), .B(KEYINPUT74), .ZN(n638) );
  NAND2_X1 U704 ( .A1(G66), .A2(n805), .ZN(n633) );
  NAND2_X1 U705 ( .A1(G54), .A2(n810), .ZN(n632) );
  NAND2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U707 ( .A1(G79), .A2(n809), .ZN(n634) );
  XNOR2_X1 U708 ( .A(KEYINPUT75), .B(n634), .ZN(n635) );
  NOR2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U711 ( .A(n640), .B(n639), .ZN(n802) );
  INV_X1 U712 ( .A(n802), .ZN(n986) );
  OR2_X1 U713 ( .A1(n646), .A2(n986), .ZN(n645) );
  INV_X1 U714 ( .A(n641), .ZN(n659) );
  NAND2_X1 U715 ( .A1(n659), .A2(G2067), .ZN(n643) );
  NAND2_X1 U716 ( .A1(G1348), .A2(n671), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U719 ( .A1(n986), .A2(n646), .ZN(n647) );
  NAND2_X1 U720 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U722 ( .A(KEYINPUT102), .B(n651), .Z(n655) );
  NAND2_X1 U723 ( .A1(G299), .A2(n652), .ZN(n653) );
  XOR2_X1 U724 ( .A(KEYINPUT28), .B(n653), .Z(n654) );
  XNOR2_X1 U725 ( .A(KEYINPUT29), .B(n656), .ZN(n663) );
  NOR2_X1 U726 ( .A1(n657), .A2(G1961), .ZN(n658) );
  XOR2_X1 U727 ( .A(KEYINPUT98), .B(n658), .Z(n661) );
  XNOR2_X1 U728 ( .A(G2078), .B(KEYINPUT25), .ZN(n967) );
  NAND2_X1 U729 ( .A1(n659), .A2(n967), .ZN(n660) );
  NAND2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n667) );
  NAND2_X1 U731 ( .A1(n667), .A2(G171), .ZN(n662) );
  NAND2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n685) );
  NOR2_X1 U733 ( .A1(G2084), .A2(n671), .ZN(n686) );
  NOR2_X1 U734 ( .A1(n687), .A2(n686), .ZN(n664) );
  NAND2_X1 U735 ( .A1(G8), .A2(n664), .ZN(n665) );
  XNOR2_X1 U736 ( .A(KEYINPUT30), .B(n665), .ZN(n666) );
  NOR2_X1 U737 ( .A1(G168), .A2(n666), .ZN(n669) );
  NOR2_X1 U738 ( .A1(G171), .A2(n667), .ZN(n668) );
  XOR2_X1 U739 ( .A(KEYINPUT31), .B(n670), .Z(n684) );
  INV_X1 U740 ( .A(G8), .ZN(n676) );
  NOR2_X1 U741 ( .A1(G2090), .A2(n671), .ZN(n673) );
  NOR2_X1 U742 ( .A1(G1971), .A2(n717), .ZN(n672) );
  NOR2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U744 ( .A1(n674), .A2(G303), .ZN(n675) );
  OR2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n678) );
  AND2_X1 U746 ( .A1(n684), .A2(n678), .ZN(n677) );
  NAND2_X1 U747 ( .A1(n685), .A2(n677), .ZN(n682) );
  INV_X1 U748 ( .A(n678), .ZN(n680) );
  AND2_X1 U749 ( .A1(G286), .A2(G8), .ZN(n679) );
  OR2_X1 U750 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U751 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U752 ( .A(n683), .B(KEYINPUT32), .ZN(n692) );
  AND2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n690) );
  AND2_X1 U754 ( .A1(G8), .A2(n686), .ZN(n688) );
  OR2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U756 ( .A1(n692), .A2(n691), .ZN(n694) );
  XNOR2_X1 U757 ( .A(n694), .B(n693), .ZN(n712) );
  NOR2_X1 U758 ( .A1(G1976), .A2(G288), .ZN(n993) );
  NOR2_X1 U759 ( .A1(G1971), .A2(G303), .ZN(n695) );
  NOR2_X1 U760 ( .A1(n993), .A2(n695), .ZN(n697) );
  INV_X1 U761 ( .A(KEYINPUT33), .ZN(n696) );
  AND2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U763 ( .A1(n712), .A2(n698), .ZN(n708) );
  INV_X1 U764 ( .A(n717), .ZN(n699) );
  NAND2_X1 U765 ( .A1(G1976), .A2(G288), .ZN(n994) );
  AND2_X1 U766 ( .A1(n699), .A2(n994), .ZN(n700) );
  NOR2_X1 U767 ( .A1(KEYINPUT33), .A2(n700), .ZN(n706) );
  NAND2_X1 U768 ( .A1(KEYINPUT33), .A2(n993), .ZN(n701) );
  XNOR2_X1 U769 ( .A(KEYINPUT104), .B(n701), .ZN(n702) );
  NOR2_X1 U770 ( .A1(n717), .A2(n702), .ZN(n703) );
  XNOR2_X1 U771 ( .A(KEYINPUT105), .B(n703), .ZN(n704) );
  XOR2_X1 U772 ( .A(G1981), .B(G305), .Z(n1005) );
  NAND2_X1 U773 ( .A1(n704), .A2(n1005), .ZN(n705) );
  NOR2_X1 U774 ( .A1(n706), .A2(n705), .ZN(n707) );
  AND2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U776 ( .A(n709), .B(KEYINPUT106), .ZN(n710) );
  INV_X1 U777 ( .A(n712), .ZN(n715) );
  NAND2_X1 U778 ( .A1(G8), .A2(G166), .ZN(n713) );
  NOR2_X1 U779 ( .A1(G2090), .A2(n713), .ZN(n714) );
  NOR2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U781 ( .A(KEYINPUT107), .B(n716), .ZN(n718) );
  NAND2_X1 U782 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U783 ( .A1(n720), .A2(n719), .ZN(n759) );
  XNOR2_X1 U784 ( .A(G1986), .B(G290), .ZN(n999) );
  NOR2_X1 U785 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U786 ( .A(n723), .B(KEYINPUT88), .ZN(n769) );
  NAND2_X1 U787 ( .A1(n999), .A2(n769), .ZN(n757) );
  XOR2_X1 U788 ( .A(G2067), .B(KEYINPUT37), .Z(n767) );
  NAND2_X1 U789 ( .A1(G140), .A2(n886), .ZN(n725) );
  NAND2_X1 U790 ( .A1(G104), .A2(n887), .ZN(n724) );
  NAND2_X1 U791 ( .A1(n725), .A2(n724), .ZN(n727) );
  XOR2_X1 U792 ( .A(KEYINPUT89), .B(KEYINPUT34), .Z(n726) );
  XNOR2_X1 U793 ( .A(n727), .B(n726), .ZN(n733) );
  NAND2_X1 U794 ( .A1(n892), .A2(G128), .ZN(n728) );
  XNOR2_X1 U795 ( .A(n728), .B(KEYINPUT90), .ZN(n730) );
  NAND2_X1 U796 ( .A1(G116), .A2(n890), .ZN(n729) );
  NAND2_X1 U797 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U798 ( .A(KEYINPUT35), .B(n731), .Z(n732) );
  NOR2_X1 U799 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U800 ( .A(KEYINPUT36), .B(n734), .Z(n912) );
  NAND2_X1 U801 ( .A1(n767), .A2(n912), .ZN(n735) );
  XNOR2_X1 U802 ( .A(KEYINPUT91), .B(n735), .ZN(n960) );
  NAND2_X1 U803 ( .A1(n769), .A2(n960), .ZN(n736) );
  XNOR2_X1 U804 ( .A(n736), .B(KEYINPUT92), .ZN(n765) );
  NAND2_X1 U805 ( .A1(G141), .A2(n886), .ZN(n737) );
  XNOR2_X1 U806 ( .A(n737), .B(KEYINPUT94), .ZN(n744) );
  NAND2_X1 U807 ( .A1(G117), .A2(n890), .ZN(n739) );
  NAND2_X1 U808 ( .A1(G129), .A2(n892), .ZN(n738) );
  NAND2_X1 U809 ( .A1(n739), .A2(n738), .ZN(n742) );
  NAND2_X1 U810 ( .A1(n887), .A2(G105), .ZN(n740) );
  XOR2_X1 U811 ( .A(KEYINPUT38), .B(n740), .Z(n741) );
  NOR2_X1 U812 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U813 ( .A1(n744), .A2(n743), .ZN(n901) );
  NAND2_X1 U814 ( .A1(G1996), .A2(n901), .ZN(n753) );
  NAND2_X1 U815 ( .A1(G107), .A2(n890), .ZN(n746) );
  NAND2_X1 U816 ( .A1(G119), .A2(n892), .ZN(n745) );
  NAND2_X1 U817 ( .A1(n746), .A2(n745), .ZN(n749) );
  NAND2_X1 U818 ( .A1(G131), .A2(n886), .ZN(n747) );
  XNOR2_X1 U819 ( .A(KEYINPUT93), .B(n747), .ZN(n748) );
  NOR2_X1 U820 ( .A1(n749), .A2(n748), .ZN(n751) );
  NAND2_X1 U821 ( .A1(n887), .A2(G95), .ZN(n750) );
  NAND2_X1 U822 ( .A1(n751), .A2(n750), .ZN(n902) );
  NAND2_X1 U823 ( .A1(G1991), .A2(n902), .ZN(n752) );
  NAND2_X1 U824 ( .A1(n753), .A2(n752), .ZN(n947) );
  NAND2_X1 U825 ( .A1(n947), .A2(n769), .ZN(n754) );
  XNOR2_X1 U826 ( .A(n754), .B(KEYINPUT95), .ZN(n762) );
  XOR2_X1 U827 ( .A(n762), .B(KEYINPUT96), .Z(n755) );
  AND2_X1 U828 ( .A1(n765), .A2(n755), .ZN(n756) );
  AND2_X1 U829 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U830 ( .A1(n759), .A2(n758), .ZN(n772) );
  NOR2_X1 U831 ( .A1(G1996), .A2(n901), .ZN(n940) );
  NOR2_X1 U832 ( .A1(G1991), .A2(n902), .ZN(n943) );
  NOR2_X1 U833 ( .A1(G1986), .A2(G290), .ZN(n760) );
  NOR2_X1 U834 ( .A1(n943), .A2(n760), .ZN(n761) );
  NOR2_X1 U835 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U836 ( .A1(n940), .A2(n763), .ZN(n764) );
  XNOR2_X1 U837 ( .A(KEYINPUT39), .B(n764), .ZN(n766) );
  NAND2_X1 U838 ( .A1(n766), .A2(n765), .ZN(n768) );
  OR2_X1 U839 ( .A1(n767), .A2(n912), .ZN(n948) );
  NAND2_X1 U840 ( .A1(n768), .A2(n948), .ZN(n770) );
  NAND2_X1 U841 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U842 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U843 ( .A(n773), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U844 ( .A1(n776), .A2(n775), .ZN(G160) );
  AND2_X1 U845 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U846 ( .A(G57), .ZN(G237) );
  INV_X1 U847 ( .A(G132), .ZN(G219) );
  INV_X1 U848 ( .A(G82), .ZN(G220) );
  NAND2_X1 U849 ( .A1(G7), .A2(G661), .ZN(n777) );
  XNOR2_X1 U850 ( .A(n777), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U851 ( .A(KEYINPUT71), .B(KEYINPUT11), .Z(n779) );
  INV_X1 U852 ( .A(G223), .ZN(n843) );
  NAND2_X1 U853 ( .A1(G567), .A2(n843), .ZN(n778) );
  XNOR2_X1 U854 ( .A(n779), .B(n778), .ZN(n780) );
  XOR2_X1 U855 ( .A(KEYINPUT70), .B(n780), .Z(G234) );
  INV_X1 U856 ( .A(G860), .ZN(n804) );
  NOR2_X1 U857 ( .A1(n804), .A2(n997), .ZN(n781) );
  XNOR2_X1 U858 ( .A(n781), .B(KEYINPUT73), .ZN(G153) );
  INV_X1 U859 ( .A(G171), .ZN(G301) );
  NAND2_X1 U860 ( .A1(G868), .A2(G301), .ZN(n783) );
  INV_X1 U861 ( .A(G868), .ZN(n824) );
  NAND2_X1 U862 ( .A1(n986), .A2(n824), .ZN(n782) );
  NAND2_X1 U863 ( .A1(n783), .A2(n782), .ZN(G284) );
  NOR2_X1 U864 ( .A1(G286), .A2(n824), .ZN(n785) );
  NOR2_X1 U865 ( .A1(G868), .A2(G299), .ZN(n784) );
  NOR2_X1 U866 ( .A1(n785), .A2(n784), .ZN(G297) );
  NAND2_X1 U867 ( .A1(G559), .A2(n804), .ZN(n786) );
  XOR2_X1 U868 ( .A(KEYINPUT79), .B(n786), .Z(n787) );
  NAND2_X1 U869 ( .A1(n802), .A2(n787), .ZN(n788) );
  XNOR2_X1 U870 ( .A(n788), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U871 ( .A1(G868), .A2(n997), .ZN(n791) );
  NAND2_X1 U872 ( .A1(n802), .A2(G868), .ZN(n789) );
  NOR2_X1 U873 ( .A1(G559), .A2(n789), .ZN(n790) );
  NOR2_X1 U874 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U875 ( .A(KEYINPUT80), .B(n792), .ZN(G282) );
  NAND2_X1 U876 ( .A1(G123), .A2(n892), .ZN(n793) );
  XNOR2_X1 U877 ( .A(n793), .B(KEYINPUT18), .ZN(n795) );
  NAND2_X1 U878 ( .A1(n890), .A2(G111), .ZN(n794) );
  NAND2_X1 U879 ( .A1(n795), .A2(n794), .ZN(n799) );
  NAND2_X1 U880 ( .A1(G135), .A2(n886), .ZN(n797) );
  NAND2_X1 U881 ( .A1(G99), .A2(n887), .ZN(n796) );
  NAND2_X1 U882 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U883 ( .A1(n799), .A2(n798), .ZN(n942) );
  XNOR2_X1 U884 ( .A(n942), .B(G2096), .ZN(n801) );
  INV_X1 U885 ( .A(G2100), .ZN(n800) );
  NAND2_X1 U886 ( .A1(n801), .A2(n800), .ZN(G156) );
  NAND2_X1 U887 ( .A1(n802), .A2(G559), .ZN(n803) );
  XOR2_X1 U888 ( .A(n997), .B(n803), .Z(n821) );
  NAND2_X1 U889 ( .A1(n804), .A2(n821), .ZN(n815) );
  NAND2_X1 U890 ( .A1(G67), .A2(n805), .ZN(n808) );
  NAND2_X1 U891 ( .A1(G93), .A2(n806), .ZN(n807) );
  NAND2_X1 U892 ( .A1(n808), .A2(n807), .ZN(n814) );
  NAND2_X1 U893 ( .A1(G80), .A2(n809), .ZN(n812) );
  NAND2_X1 U894 ( .A1(G55), .A2(n810), .ZN(n811) );
  NAND2_X1 U895 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U896 ( .A1(n814), .A2(n813), .ZN(n823) );
  XOR2_X1 U897 ( .A(n815), .B(n823), .Z(G145) );
  XNOR2_X1 U898 ( .A(G166), .B(n823), .ZN(n819) );
  XNOR2_X1 U899 ( .A(G288), .B(KEYINPUT19), .ZN(n817) );
  XOR2_X1 U900 ( .A(G290), .B(G299), .Z(n816) );
  XNOR2_X1 U901 ( .A(n817), .B(n816), .ZN(n818) );
  XNOR2_X1 U902 ( .A(n819), .B(n818), .ZN(n820) );
  XNOR2_X1 U903 ( .A(n820), .B(G305), .ZN(n917) );
  XOR2_X1 U904 ( .A(n917), .B(n821), .Z(n822) );
  NOR2_X1 U905 ( .A1(n824), .A2(n822), .ZN(n826) );
  AND2_X1 U906 ( .A1(n824), .A2(n823), .ZN(n825) );
  NOR2_X1 U907 ( .A1(n826), .A2(n825), .ZN(G295) );
  XOR2_X1 U908 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n830) );
  NAND2_X1 U909 ( .A1(G2078), .A2(G2084), .ZN(n827) );
  XOR2_X1 U910 ( .A(KEYINPUT20), .B(n827), .Z(n828) );
  NAND2_X1 U911 ( .A1(n828), .A2(G2090), .ZN(n829) );
  XNOR2_X1 U912 ( .A(n830), .B(n829), .ZN(n831) );
  NAND2_X1 U913 ( .A1(G2072), .A2(n831), .ZN(G158) );
  XNOR2_X1 U914 ( .A(KEYINPUT86), .B(G44), .ZN(n832) );
  XNOR2_X1 U915 ( .A(n832), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U916 ( .A1(G220), .A2(G219), .ZN(n833) );
  XOR2_X1 U917 ( .A(KEYINPUT22), .B(n833), .Z(n834) );
  NOR2_X1 U918 ( .A1(G218), .A2(n834), .ZN(n835) );
  NAND2_X1 U919 ( .A1(G96), .A2(n835), .ZN(n848) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n848), .ZN(n839) );
  NAND2_X1 U921 ( .A1(G69), .A2(G120), .ZN(n836) );
  NOR2_X1 U922 ( .A1(G237), .A2(n836), .ZN(n837) );
  NAND2_X1 U923 ( .A1(G108), .A2(n837), .ZN(n847) );
  NAND2_X1 U924 ( .A1(G567), .A2(n847), .ZN(n838) );
  NAND2_X1 U925 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U926 ( .A(KEYINPUT87), .B(n840), .ZN(G319) );
  INV_X1 U927 ( .A(G319), .ZN(n842) );
  NAND2_X1 U928 ( .A1(G661), .A2(G483), .ZN(n841) );
  NOR2_X1 U929 ( .A1(n842), .A2(n841), .ZN(n846) );
  NAND2_X1 U930 ( .A1(n846), .A2(G36), .ZN(G176) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U933 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n845) );
  NAND2_X1 U935 ( .A1(n846), .A2(n845), .ZN(G188) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(G69), .ZN(G235) );
  NOR2_X1 U940 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U941 ( .A(n849), .B(KEYINPUT110), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U943 ( .A(G1986), .B(KEYINPUT41), .ZN(n859) );
  XOR2_X1 U944 ( .A(G1976), .B(G1971), .Z(n851) );
  XNOR2_X1 U945 ( .A(G1961), .B(G1956), .ZN(n850) );
  XNOR2_X1 U946 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U947 ( .A(G1981), .B(G1966), .Z(n853) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U949 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U950 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U951 ( .A(G2474), .B(KEYINPUT112), .ZN(n856) );
  XNOR2_X1 U952 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U953 ( .A(n859), .B(n858), .ZN(G229) );
  XOR2_X1 U954 ( .A(KEYINPUT111), .B(G2084), .Z(n861) );
  XNOR2_X1 U955 ( .A(G2090), .B(G2072), .ZN(n860) );
  XNOR2_X1 U956 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U957 ( .A(n862), .B(G2100), .Z(n864) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2078), .ZN(n863) );
  XNOR2_X1 U959 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U960 ( .A(G2096), .B(G2678), .Z(n866) );
  XNOR2_X1 U961 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n865) );
  XNOR2_X1 U962 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U963 ( .A(n868), .B(n867), .Z(G227) );
  NAND2_X1 U964 ( .A1(G124), .A2(n892), .ZN(n869) );
  XOR2_X1 U965 ( .A(KEYINPUT44), .B(n869), .Z(n870) );
  XNOR2_X1 U966 ( .A(n870), .B(KEYINPUT113), .ZN(n872) );
  NAND2_X1 U967 ( .A1(G136), .A2(n886), .ZN(n871) );
  NAND2_X1 U968 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U969 ( .A(KEYINPUT114), .B(n873), .ZN(n877) );
  NAND2_X1 U970 ( .A1(G112), .A2(n890), .ZN(n875) );
  NAND2_X1 U971 ( .A1(G100), .A2(n887), .ZN(n874) );
  NAND2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n876) );
  NOR2_X1 U973 ( .A1(n877), .A2(n876), .ZN(G162) );
  NAND2_X1 U974 ( .A1(G118), .A2(n890), .ZN(n879) );
  NAND2_X1 U975 ( .A1(G130), .A2(n892), .ZN(n878) );
  NAND2_X1 U976 ( .A1(n879), .A2(n878), .ZN(n884) );
  NAND2_X1 U977 ( .A1(G142), .A2(n886), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G106), .A2(n887), .ZN(n880) );
  NAND2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U980 ( .A(KEYINPUT45), .B(n882), .Z(n883) );
  NOR2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(n885), .B(G162), .Z(n900) );
  NAND2_X1 U983 ( .A1(G139), .A2(n886), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G103), .A2(n887), .ZN(n888) );
  NAND2_X1 U985 ( .A1(n889), .A2(n888), .ZN(n898) );
  NAND2_X1 U986 ( .A1(n890), .A2(G115), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n891), .B(KEYINPUT116), .ZN(n894) );
  NAND2_X1 U988 ( .A1(G127), .A2(n892), .ZN(n893) );
  NAND2_X1 U989 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U990 ( .A(KEYINPUT47), .B(n895), .ZN(n896) );
  XNOR2_X1 U991 ( .A(KEYINPUT117), .B(n896), .ZN(n897) );
  NOR2_X1 U992 ( .A1(n898), .A2(n897), .ZN(n950) );
  XNOR2_X1 U993 ( .A(G160), .B(n950), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n900), .B(n899), .ZN(n905) );
  XNOR2_X1 U995 ( .A(n942), .B(n901), .ZN(n903) );
  XNOR2_X1 U996 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U997 ( .A(n905), .B(n904), .Z(n910) );
  XOR2_X1 U998 ( .A(KEYINPUT115), .B(KEYINPUT118), .Z(n907) );
  XNOR2_X1 U999 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1001 ( .A(G164), .B(n908), .ZN(n909) );
  XNOR2_X1 U1002 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1003 ( .A(n912), .B(n911), .Z(n913) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n913), .ZN(n914) );
  XOR2_X1 U1005 ( .A(KEYINPUT119), .B(n914), .Z(G395) );
  XNOR2_X1 U1006 ( .A(n997), .B(KEYINPUT120), .ZN(n916) );
  XNOR2_X1 U1007 ( .A(G171), .B(n986), .ZN(n915) );
  XNOR2_X1 U1008 ( .A(n916), .B(n915), .ZN(n919) );
  XNOR2_X1 U1009 ( .A(G286), .B(n917), .ZN(n918) );
  XNOR2_X1 U1010 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n920), .ZN(n921) );
  XOR2_X1 U1012 ( .A(KEYINPUT121), .B(n921), .Z(G397) );
  XNOR2_X1 U1013 ( .A(G2446), .B(KEYINPUT108), .ZN(n931) );
  XOR2_X1 U1014 ( .A(KEYINPUT109), .B(G2427), .Z(n923) );
  XNOR2_X1 U1015 ( .A(G2435), .B(G2438), .ZN(n922) );
  XNOR2_X1 U1016 ( .A(n923), .B(n922), .ZN(n927) );
  XOR2_X1 U1017 ( .A(G2454), .B(G2430), .Z(n925) );
  XNOR2_X1 U1018 ( .A(G1348), .B(G1341), .ZN(n924) );
  XNOR2_X1 U1019 ( .A(n925), .B(n924), .ZN(n926) );
  XOR2_X1 U1020 ( .A(n927), .B(n926), .Z(n929) );
  XNOR2_X1 U1021 ( .A(G2443), .B(G2451), .ZN(n928) );
  XNOR2_X1 U1022 ( .A(n929), .B(n928), .ZN(n930) );
  XNOR2_X1 U1023 ( .A(n931), .B(n930), .ZN(n932) );
  NAND2_X1 U1024 ( .A1(n932), .A2(G14), .ZN(n938) );
  NAND2_X1 U1025 ( .A1(G319), .A2(n938), .ZN(n935) );
  NOR2_X1 U1026 ( .A1(G229), .A2(G227), .ZN(n933) );
  XNOR2_X1 U1027 ( .A(KEYINPUT49), .B(n933), .ZN(n934) );
  NOR2_X1 U1028 ( .A1(n935), .A2(n934), .ZN(n937) );
  NOR2_X1 U1029 ( .A1(G395), .A2(G397), .ZN(n936) );
  NAND2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(G225) );
  INV_X1 U1031 ( .A(G225), .ZN(G308) );
  INV_X1 U1032 ( .A(G108), .ZN(G238) );
  INV_X1 U1033 ( .A(n938), .ZN(G401) );
  XOR2_X1 U1034 ( .A(G2090), .B(G162), .Z(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1036 ( .A(KEYINPUT51), .B(n941), .Z(n958) );
  XNOR2_X1 U1037 ( .A(G160), .B(G2084), .ZN(n945) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n949) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n956) );
  XOR2_X1 U1042 ( .A(G164), .B(G2078), .Z(n953) );
  XNOR2_X1 U1043 ( .A(n951), .B(n950), .ZN(n952) );
  NOR2_X1 U1044 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1045 ( .A(KEYINPUT50), .B(n954), .Z(n955) );
  NOR2_X1 U1046 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1047 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1048 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1049 ( .A(KEYINPUT52), .B(n961), .ZN(n962) );
  INV_X1 U1050 ( .A(KEYINPUT55), .ZN(n982) );
  NAND2_X1 U1051 ( .A1(n962), .A2(n982), .ZN(n963) );
  NAND2_X1 U1052 ( .A1(n963), .A2(G29), .ZN(n1042) );
  XNOR2_X1 U1053 ( .A(G2090), .B(G35), .ZN(n977) );
  XOR2_X1 U1054 ( .A(G1991), .B(G25), .Z(n964) );
  NAND2_X1 U1055 ( .A1(n964), .A2(G28), .ZN(n974) );
  XNOR2_X1 U1056 ( .A(G2067), .B(G26), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(G33), .B(G2072), .ZN(n965) );
  NOR2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n972) );
  XOR2_X1 U1059 ( .A(n967), .B(G27), .Z(n970) );
  XOR2_X1 U1060 ( .A(n968), .B(G32), .Z(n969) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1063 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(KEYINPUT53), .B(n975), .ZN(n976) );
  NOR2_X1 U1065 ( .A1(n977), .A2(n976), .ZN(n980) );
  XOR2_X1 U1066 ( .A(G2084), .B(G34), .Z(n978) );
  XNOR2_X1 U1067 ( .A(KEYINPUT54), .B(n978), .ZN(n979) );
  NAND2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1069 ( .A(n982), .B(n981), .ZN(n984) );
  INV_X1 U1070 ( .A(G29), .ZN(n983) );
  NAND2_X1 U1071 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1072 ( .A1(G11), .A2(n985), .ZN(n1040) );
  XNOR2_X1 U1073 ( .A(G16), .B(KEYINPUT56), .ZN(n1012) );
  XNOR2_X1 U1074 ( .A(G171), .B(G1961), .ZN(n992) );
  XOR2_X1 U1075 ( .A(G1348), .B(n986), .Z(n988) );
  XOR2_X1 U1076 ( .A(G299), .B(G1956), .Z(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(G1971), .B(G303), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n1003) );
  INV_X1 U1081 ( .A(n993), .ZN(n995) );
  NAND2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(n996), .B(KEYINPUT123), .ZN(n1001) );
  XNOR2_X1 U1084 ( .A(G1341), .B(n997), .ZN(n998) );
  NOR2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1087 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1088 ( .A(KEYINPUT124), .B(n1004), .ZN(n1010) );
  XNOR2_X1 U1089 ( .A(G1966), .B(G168), .ZN(n1006) );
  NAND2_X1 U1090 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1091 ( .A(n1007), .B(KEYINPUT57), .ZN(n1008) );
  XNOR2_X1 U1092 ( .A(KEYINPUT122), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1093 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1094 ( .A1(n1012), .A2(n1011), .ZN(n1038) );
  INV_X1 U1095 ( .A(G16), .ZN(n1036) );
  XOR2_X1 U1096 ( .A(G1971), .B(G22), .Z(n1015) );
  XOR2_X1 U1097 ( .A(G23), .B(KEYINPUT126), .Z(n1013) );
  XNOR2_X1 U1098 ( .A(n1013), .B(G1976), .ZN(n1014) );
  NAND2_X1 U1099 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  XNOR2_X1 U1100 ( .A(G24), .B(G1986), .ZN(n1016) );
  NOR2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1102 ( .A(KEYINPUT58), .B(n1018), .Z(n1033) );
  XOR2_X1 U1103 ( .A(G1961), .B(G5), .Z(n1028) );
  XNOR2_X1 U1104 ( .A(G1348), .B(KEYINPUT59), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(n1019), .B(G4), .ZN(n1023) );
  XNOR2_X1 U1106 ( .A(G1341), .B(G19), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(G1981), .B(G6), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1025) );
  XNOR2_X1 U1110 ( .A(G20), .B(G1956), .ZN(n1024) );
  NOR2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1112 ( .A(KEYINPUT60), .B(n1026), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1030) );
  XNOR2_X1 U1114 ( .A(G21), .B(G1966), .ZN(n1029) );
  NOR2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1116 ( .A(KEYINPUT125), .B(n1031), .ZN(n1032) );
  NOR2_X1 U1117 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1118 ( .A(KEYINPUT61), .B(n1034), .ZN(n1035) );
  NAND2_X1 U1119 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1120 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NOR2_X1 U1121 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  NAND2_X1 U1122 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  XNOR2_X1 U1123 ( .A(n1043), .B(KEYINPUT62), .ZN(n1044) );
  XNOR2_X1 U1124 ( .A(KEYINPUT127), .B(n1044), .ZN(G311) );
  INV_X1 U1125 ( .A(G311), .ZN(G150) );
endmodule

