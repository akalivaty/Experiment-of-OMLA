//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT73), .Z(new_n189));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n191), .B1(KEYINPUT0), .B2(G128), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n192), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT64), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT0), .A2(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n190), .B1(new_n197), .B2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(G143), .B(G146), .ZN(new_n203));
  AND2_X1   g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n204), .B1(KEYINPUT64), .B2(new_n198), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n195), .A2(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n193), .A2(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n206), .A2(KEYINPUT65), .A3(new_n209), .A4(new_n192), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n202), .A2(new_n205), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT70), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT70), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n202), .A2(new_n213), .A3(new_n210), .A4(new_n205), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  OR2_X1    g030(.A1(KEYINPUT66), .A2(G134), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT66), .A2(G134), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(G137), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G134), .ZN(new_n220));
  INV_X1    g034(.A(G137), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n216), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n217), .A2(new_n218), .ZN(new_n224));
  NOR3_X1   g038(.A1(new_n224), .A2(KEYINPUT11), .A3(G137), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT67), .B(G131), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n223), .B2(new_n225), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n215), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n220), .A2(KEYINPUT68), .A3(G137), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n224), .B2(G137), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT68), .B1(new_n220), .B2(G137), .ZN(new_n235));
  OAI21_X1  g049(.A(G131), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT1), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n203), .A2(new_n237), .A3(G128), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n196), .A2(KEYINPUT1), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n238), .B(new_n239), .C1(G128), .C2(new_n203), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n230), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n232), .A2(KEYINPUT30), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G119), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G116), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT69), .B(G116), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(new_n243), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT2), .B(G113), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT30), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n211), .B1(new_n227), .B2(new_n230), .ZN(new_n250));
  INV_X1    g064(.A(new_n241), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n242), .A2(new_n248), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n251), .B1(new_n215), .B2(new_n231), .ZN(new_n254));
  XOR2_X1   g068(.A(new_n246), .B(new_n247), .Z(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G101), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT27), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT71), .B(G237), .ZN(new_n259));
  INV_X1    g073(.A(G953), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n258), .B1(new_n261), .B2(G210), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT26), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(new_n258), .A3(G210), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n264), .B1(new_n263), .B2(new_n265), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n257), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n268), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(G101), .A3(new_n266), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n253), .A2(new_n256), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT72), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n253), .A2(new_n272), .A3(new_n275), .A4(new_n256), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n274), .A2(KEYINPUT31), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT31), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n256), .A2(KEYINPUT28), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n254), .A2(new_n282), .A3(new_n255), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n272), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n189), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n187), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n286), .B1(new_n277), .B2(new_n279), .ZN(new_n291));
  OAI211_X1 g105(.A(KEYINPUT74), .B(KEYINPUT32), .C1(new_n291), .C2(new_n189), .ZN(new_n292));
  OR2_X1    g106(.A1(new_n254), .A2(new_n255), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n254), .A2(new_n282), .A3(new_n255), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n282), .B1(new_n254), .B2(new_n255), .ZN(new_n295));
  OAI211_X1 g109(.A(KEYINPUT29), .B(new_n293), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n272), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT75), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n254), .A2(new_n255), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n299), .B1(new_n281), .B2(new_n283), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT29), .A4(new_n272), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n298), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n284), .A2(new_n285), .A3(new_n272), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n253), .A2(new_n256), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n297), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n298), .A2(new_n302), .A3(KEYINPUT76), .A4(new_n303), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n306), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n290), .A2(new_n292), .B1(G472), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G128), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT23), .A3(G119), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT23), .B1(new_n315), .B2(G119), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n315), .A2(G119), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n243), .A2(G128), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT78), .A3(KEYINPUT23), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G110), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n322), .A2(new_n323), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT24), .B(G110), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n332), .A2(KEYINPUT80), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(KEYINPUT80), .ZN(new_n334));
  XNOR2_X1  g148(.A(G125), .B(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n195), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G140), .ZN(new_n338));
  MUX2_X1   g152(.A(new_n338), .B(new_n335), .S(KEYINPUT16), .Z(new_n339));
  OR2_X1    g153(.A1(new_n339), .A2(new_n195), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n333), .A2(new_n334), .A3(new_n336), .A4(new_n340), .ZN(new_n341));
  OR2_X1    g155(.A1(new_n326), .A2(new_n327), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n339), .B(new_n195), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n343), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n329), .A2(new_n330), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n344), .A2(new_n345), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(KEYINPUT22), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(G137), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n341), .A2(new_n348), .A3(new_n352), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n303), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT25), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n354), .A2(KEYINPUT25), .A3(new_n303), .A4(new_n355), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G217), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(G234), .B2(new_n303), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n364));
  INV_X1    g178(.A(new_n355), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n352), .B1(new_n341), .B2(new_n348), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n362), .A2(G902), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n354), .A2(KEYINPUT81), .A3(new_n355), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT82), .B1(new_n363), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n362), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(new_n358), .B2(new_n359), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n374), .A2(new_n370), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n314), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G469), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G104), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT3), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n382), .A2(G104), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n381), .A2(new_n387), .A3(new_n382), .A4(G104), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n384), .A2(new_n257), .A3(new_n386), .A4(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G104), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(G107), .ZN(new_n391));
  OAI21_X1  g205(.A(G101), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n240), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n380), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n380), .A3(new_n394), .ZN(new_n397));
  INV_X1    g211(.A(new_n393), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n396), .A2(new_n397), .B1(KEYINPUT10), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n384), .A2(new_n386), .A3(new_n388), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G101), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT4), .A3(new_n389), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n403), .A3(G101), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(new_n212), .B2(new_n214), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n231), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n399), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n240), .B1(new_n389), .B2(new_n392), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n231), .B1(new_n398), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT12), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n411), .B(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G140), .ZN(new_n414));
  INV_X1    g228(.A(G227), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(G953), .ZN(new_n416));
  XOR2_X1   g230(.A(new_n414), .B(new_n416), .Z(new_n417));
  AND3_X1   g231(.A1(new_n409), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n397), .ZN(new_n419));
  OAI22_X1  g233(.A1(new_n419), .A2(new_n395), .B1(new_n394), .B2(new_n393), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n231), .B1(new_n420), .B2(new_n406), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n417), .B1(new_n409), .B2(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n379), .B(new_n303), .C1(new_n418), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(G469), .A2(G902), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n409), .A2(new_n413), .ZN(new_n425));
  INV_X1    g239(.A(new_n417), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n409), .A2(new_n421), .A3(new_n417), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(G469), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n423), .A2(new_n424), .A3(new_n429), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT9), .B(G234), .Z(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G221), .B1(new_n432), .B2(G902), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G214), .B1(G237), .B2(G902), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT85), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n436), .B1(new_n405), .B2(new_n255), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT5), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n243), .A3(G116), .ZN(new_n439));
  OAI211_X1 g253(.A(G113), .B(new_n439), .C1(new_n246), .C2(new_n438), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(new_n246), .B2(new_n247), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n389), .A2(new_n392), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  XOR2_X1   g257(.A(G110), .B(G122), .Z(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n248), .A2(new_n402), .A3(KEYINPUT85), .A4(new_n404), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n437), .A2(new_n443), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n211), .A2(new_n337), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n240), .A2(new_n337), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n260), .A2(G224), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT86), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT7), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n449), .A2(KEYINPUT7), .A3(new_n454), .A4(new_n450), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n441), .B(new_n442), .Z(new_n459));
  XOR2_X1   g273(.A(KEYINPUT88), .B(KEYINPUT8), .Z(new_n460));
  XNOR2_X1  g274(.A(new_n444), .B(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n458), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT89), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n448), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n458), .B(KEYINPUT89), .C1(new_n459), .C2(new_n462), .ZN(new_n466));
  AOI21_X1  g280(.A(G902), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n437), .A2(new_n443), .A3(new_n446), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n444), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(KEYINPUT6), .A3(new_n447), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n451), .B(new_n454), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(new_n472), .A3(new_n444), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n470), .A2(KEYINPUT87), .A3(new_n471), .A4(new_n473), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n467), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G210), .B1(G237), .B2(G902), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(KEYINPUT90), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n467), .A2(new_n476), .A3(new_n480), .A4(new_n477), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n434), .A2(new_n435), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n259), .A2(G214), .A3(new_n260), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n193), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n259), .A2(G143), .A3(G214), .A4(new_n260), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n228), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT91), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT17), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT91), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n488), .A2(new_n492), .A3(new_n228), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n486), .A2(new_n487), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n229), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n490), .A2(new_n491), .A3(new_n493), .A4(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n345), .B1(new_n496), .B2(KEYINPUT92), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n492), .B1(new_n488), .B2(new_n228), .ZN(new_n498));
  AOI211_X1 g312(.A(KEYINPUT91), .B(new_n229), .C1(new_n486), .C2(new_n487), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT17), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n498), .A2(new_n499), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT92), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n501), .A2(new_n502), .A3(new_n491), .A4(new_n495), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n497), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(G113), .B(G122), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(new_n390), .ZN(new_n506));
  NAND2_X1  g320(.A1(KEYINPUT18), .A2(G131), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n494), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n335), .B(G146), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n504), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n506), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n335), .B(KEYINPUT19), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n340), .B1(new_n515), .B2(G146), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(new_n501), .B2(new_n495), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n513), .B1(new_n510), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(G475), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n520), .A3(new_n303), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT20), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n519), .A2(KEYINPUT20), .A3(new_n520), .A4(new_n303), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT93), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n504), .A2(new_n511), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n527), .B1(new_n528), .B2(new_n513), .ZN(new_n529));
  AOI211_X1 g343(.A(KEYINPUT93), .B(new_n506), .C1(new_n504), .C2(new_n511), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n512), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n303), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G475), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n260), .A2(G952), .ZN(new_n534));
  NAND2_X1  g348(.A1(G234), .A2(G237), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g350(.A(KEYINPUT21), .B(G898), .Z(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(G902), .A3(G953), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G122), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n245), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(G116), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G107), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n382), .B(new_n542), .C1(new_n245), .C2(new_n540), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n315), .A2(G143), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n547), .A2(KEYINPUT13), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(KEYINPUT13), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n315), .A2(G143), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G134), .ZN(new_n552));
  INV_X1    g366(.A(new_n547), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n550), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n224), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n546), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n546), .A2(KEYINPUT94), .A3(new_n552), .A4(new_n556), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT14), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n541), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n542), .A2(KEYINPUT96), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT95), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n541), .B2(new_n562), .ZN(new_n567));
  OAI211_X1 g381(.A(KEYINPUT95), .B(KEYINPUT14), .C1(new_n245), .C2(new_n540), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n541), .A2(KEYINPUT96), .A3(new_n562), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n565), .A2(new_n567), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(G107), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n554), .A2(new_n217), .A3(new_n218), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n556), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(new_n545), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n561), .A2(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n432), .A2(new_n361), .A3(G953), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n561), .A2(new_n574), .A3(new_n576), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n303), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(KEYINPUT97), .A3(new_n303), .ZN(new_n584));
  INV_X1    g398(.A(G478), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n586));
  AOI211_X1 g400(.A(KEYINPUT15), .B(new_n585), .C1(new_n582), .C2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n583), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n585), .A2(KEYINPUT15), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n581), .A2(new_n586), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n526), .A2(new_n533), .A3(new_n539), .A4(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n484), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n378), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  INV_X1    g409(.A(KEYINPUT103), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n476), .A2(new_n477), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT100), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n479), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n479), .A2(new_n598), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n597), .A2(new_n467), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n478), .A2(new_n598), .A3(new_n479), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n526), .A2(new_n533), .ZN(new_n604));
  INV_X1    g418(.A(new_n579), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n576), .B1(new_n561), .B2(new_n574), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT101), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT33), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n578), .B(new_n579), .C1(KEYINPUT101), .C2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(G478), .B(new_n303), .C1(new_n610), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT102), .ZN(new_n615));
  INV_X1    g429(.A(new_n583), .ZN(new_n616));
  INV_X1    g430(.A(new_n584), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n585), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n580), .B(KEYINPUT33), .C1(new_n608), .C2(new_n606), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n612), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT102), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n620), .A2(new_n621), .A3(G478), .A4(new_n303), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n615), .A2(new_n618), .A3(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n603), .A2(new_n604), .A3(new_n435), .A4(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n539), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n596), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n520), .B1(new_n531), .B2(new_n303), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n623), .B1(new_n627), .B2(new_n525), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n601), .A2(new_n602), .A3(new_n435), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(KEYINPUT103), .A3(new_n539), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(G472), .B1(new_n291), .B2(G902), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n633), .A2(KEYINPUT99), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(KEYINPUT99), .ZN(new_n635));
  INV_X1    g449(.A(new_n288), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .A4(new_n434), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n377), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  NOR3_X1   g455(.A1(new_n637), .A2(new_n377), .A3(new_n625), .ZN(new_n642));
  INV_X1    g456(.A(new_n591), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n526), .A2(new_n533), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n629), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  AND2_X1   g462(.A1(new_n634), .A2(new_n635), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n353), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n349), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n368), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n363), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n649), .A2(new_n593), .A3(new_n636), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT104), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT37), .B(G110), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  NAND2_X1  g471(.A1(new_n290), .A2(new_n292), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n313), .A2(G472), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n260), .A2(G900), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(G902), .A3(new_n535), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(new_n536), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n644), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n434), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n629), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n660), .A2(new_n653), .A3(new_n668), .A4(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n653), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n658), .B2(new_n659), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n675), .A2(KEYINPUT106), .A3(new_n668), .A4(new_n670), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  INV_X1    g492(.A(new_n435), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n666), .B(KEYINPUT108), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT39), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n434), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n674), .B1(new_n683), .B2(KEYINPUT40), .ZN(new_n684));
  AOI211_X1 g498(.A(new_n679), .B(new_n684), .C1(KEYINPUT40), .C2(new_n683), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n482), .A2(new_n483), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT38), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n604), .A2(new_n643), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n274), .A2(new_n276), .ZN(new_n690));
  INV_X1    g504(.A(new_n256), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n297), .B1(new_n691), .B2(new_n299), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n693), .A2(KEYINPUT107), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n303), .B1(new_n693), .B2(KEYINPUT107), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n658), .A2(new_n696), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n685), .A2(new_n689), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(new_n193), .ZN(G45));
  OAI211_X1 g513(.A(new_n623), .B(new_n666), .C1(new_n627), .C2(new_n525), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n660), .A2(new_n653), .A3(new_n670), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  OAI21_X1  g517(.A(new_n303), .B1(new_n418), .B2(new_n422), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n433), .A3(new_n423), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n314), .A2(new_n377), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT103), .B1(new_n630), .B2(new_n539), .ZN(new_n708));
  NOR4_X1   g522(.A1(new_n628), .A2(new_n629), .A3(new_n596), .A4(new_n625), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT41), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G113), .ZN(G15));
  INV_X1    g526(.A(new_n377), .ZN(new_n713));
  INV_X1    g527(.A(new_n706), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n539), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n660), .A2(new_n713), .A3(new_n645), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  INV_X1    g532(.A(new_n592), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n629), .A2(new_n706), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n675), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT109), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  NOR2_X1   g537(.A1(new_n688), .A2(new_n629), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n633), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n374), .A2(new_n370), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n280), .B1(new_n272), .B2(new_n300), .ZN(new_n728));
  INV_X1    g542(.A(new_n189), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(KEYINPUT110), .B(G472), .C1(new_n291), .C2(G902), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n726), .A2(new_n727), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n716), .B(new_n724), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  AND4_X1   g551(.A1(new_n653), .A2(new_n726), .A3(new_n730), .A4(new_n731), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n701), .A3(new_n720), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  INV_X1    g554(.A(new_n727), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n313), .A2(G472), .B1(KEYINPUT32), .B2(new_n288), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n636), .A2(new_n187), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n686), .A2(new_n435), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n700), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(new_n746), .A3(KEYINPUT42), .A4(new_n434), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n686), .A2(new_n434), .A3(new_n435), .ZN(new_n749));
  NOR4_X1   g563(.A1(new_n314), .A2(new_n377), .A3(new_n700), .A4(new_n749), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n747), .B(new_n748), .C1(new_n750), .C2(KEYINPUT42), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n749), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n660), .A2(new_n713), .A3(new_n701), .A4(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n748), .B1(new_n756), .B2(new_n747), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G131), .ZN(G33));
  NAND4_X1  g573(.A1(new_n660), .A2(new_n713), .A3(new_n668), .A4(new_n753), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  INV_X1    g575(.A(new_n623), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n604), .A2(new_n762), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n763), .A2(KEYINPUT43), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(KEYINPUT43), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n766), .A2(KEYINPUT114), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n649), .A2(new_n636), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(KEYINPUT114), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n767), .A2(new_n768), .A3(new_n653), .A4(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n745), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(new_n770), .B2(new_n771), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n427), .A2(new_n428), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT45), .ZN(new_n776));
  OAI21_X1  g590(.A(G469), .B1(new_n776), .B2(G902), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(KEYINPUT113), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(KEYINPUT113), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n779), .A2(new_n423), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n433), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n681), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n772), .A2(new_n774), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n221), .ZN(G39));
  XNOR2_X1  g601(.A(new_n783), .B(KEYINPUT47), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AND4_X1   g603(.A1(new_n314), .A2(new_n789), .A3(new_n377), .A4(new_n746), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(G140), .Z(G42));
  NAND2_X1  g605(.A1(new_n705), .A2(new_n423), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n792), .A2(KEYINPUT49), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(KEYINPUT49), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n687), .A2(new_n727), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n763), .A2(new_n433), .ZN(new_n796));
  OR4_X1    g610(.A1(new_n679), .A2(new_n795), .A3(new_n697), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n697), .A2(new_n536), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n745), .A2(new_n706), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n713), .A3(new_n799), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n800), .A2(new_n628), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n800), .A2(new_n604), .A3(new_n623), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n766), .A2(new_n536), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n734), .A2(new_n735), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n805), .A2(new_n714), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n679), .A3(new_n687), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n806), .A2(KEYINPUT50), .A3(new_n679), .A4(new_n687), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n802), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n803), .A2(new_n738), .A3(new_n799), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n805), .A2(new_n773), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n792), .A2(new_n433), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n813), .B1(new_n789), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n811), .A2(KEYINPUT51), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n803), .A2(new_n744), .A3(new_n799), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n803), .A2(KEYINPUT120), .A3(new_n744), .A4(new_n799), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(KEYINPUT48), .A3(new_n820), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n821), .B(new_n534), .C1(KEYINPUT48), .C2(new_n819), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(new_n720), .B2(new_n805), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n816), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n814), .B(KEYINPUT119), .Z(new_n826));
  OAI21_X1  g640(.A(new_n813), .B1(new_n789), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n811), .A2(new_n827), .A3(new_n812), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n824), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n702), .A2(new_n739), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n673), .B2(new_n676), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n674), .A2(new_n434), .A3(new_n666), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT116), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n697), .A3(new_n724), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n830), .ZN(new_n836));
  AND4_X1   g650(.A1(KEYINPUT52), .A2(new_n677), .A3(new_n836), .A4(new_n834), .ZN(new_n837));
  OR3_X1    g651(.A1(new_n835), .A2(new_n837), .A3(KEYINPUT117), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n738), .A2(KEYINPUT115), .A3(new_n701), .A4(new_n753), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n760), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n726), .A2(new_n653), .A3(new_n730), .A4(new_n731), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n700), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT115), .B1(new_n843), .B2(new_n753), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n604), .A2(new_n643), .A3(new_n667), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n660), .A2(new_n653), .A3(new_n845), .A4(new_n753), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n841), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n594), .A2(new_n654), .A3(new_n721), .A4(new_n717), .ZN(new_n848));
  AOI211_X1 g662(.A(new_n679), .B(new_n686), .C1(new_n628), .C2(new_n644), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n632), .A2(new_n707), .B1(new_n642), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n847), .A2(new_n736), .A3(new_n848), .A4(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n752), .A2(new_n757), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n837), .A2(KEYINPUT117), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n838), .A2(new_n839), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n638), .A2(new_n539), .A3(new_n849), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n736), .A2(new_n856), .A3(new_n710), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n738), .A2(new_n701), .A3(new_n753), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n675), .A2(new_n753), .A3(new_n845), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n760), .A3(new_n861), .A4(new_n840), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n594), .A2(new_n654), .A3(new_n721), .A4(new_n717), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n857), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n758), .B(new_n864), .C1(new_n835), .C2(new_n837), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT53), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n855), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT54), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n756), .A2(new_n747), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n851), .A2(new_n839), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n838), .A2(new_n854), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n677), .A2(new_n836), .A3(new_n834), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT52), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n831), .A2(KEYINPUT52), .A3(new_n834), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI211_X1 g693(.A(new_n874), .B(KEYINPUT53), .C1(new_n853), .C2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT118), .B1(new_n865), .B2(new_n839), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n872), .B(new_n873), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n801), .A2(new_n829), .A3(new_n869), .A4(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(G952), .A2(G953), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n797), .B1(new_n883), .B2(new_n884), .ZN(G75));
  OAI21_X1  g699(.A(new_n872), .B1(new_n880), .B2(new_n881), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(G210), .A3(G902), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT56), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT121), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n887), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n470), .A2(new_n473), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(new_n471), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT55), .Z(new_n895));
  AND3_X1   g709(.A1(new_n890), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n895), .B1(new_n890), .B2(new_n892), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n260), .A2(G952), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(G51));
  NAND2_X1  g713(.A1(new_n886), .A2(KEYINPUT54), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(KEYINPUT122), .A3(new_n882), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n886), .A2(new_n902), .A3(KEYINPUT54), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n424), .B(KEYINPUT57), .Z(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT123), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n418), .A2(new_n422), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n901), .A2(new_n908), .A3(new_n903), .A4(new_n904), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n886), .A2(G902), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n911), .A2(G469), .A3(new_n776), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n898), .B1(new_n910), .B2(new_n912), .ZN(G54));
  NAND3_X1  g727(.A1(new_n911), .A2(KEYINPUT58), .A3(G475), .ZN(new_n914));
  INV_X1    g728(.A(new_n519), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n916), .A2(new_n917), .A3(new_n898), .ZN(G60));
  INV_X1    g732(.A(new_n898), .ZN(new_n919));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT59), .Z(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n869), .B2(new_n882), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n919), .B1(new_n922), .B2(new_n620), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n901), .A2(new_n903), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n921), .B1(new_n619), .B2(new_n612), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(G63));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT125), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT60), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n886), .A2(new_n651), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n886), .A2(new_n929), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n367), .A2(new_n369), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n919), .B(new_n930), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT124), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT61), .ZN(G66));
  NAND2_X1  g750(.A1(new_n537), .A2(G224), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(G953), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n848), .A2(new_n850), .A3(new_n736), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n938), .B1(new_n940), .B2(G953), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n893), .B1(G898), .B2(new_n260), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(G69));
  NOR2_X1   g757(.A1(new_n786), .A2(new_n790), .ZN(new_n944));
  INV_X1    g758(.A(new_n698), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n831), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT62), .Z(new_n947));
  NAND2_X1  g761(.A1(new_n628), .A2(new_n644), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n378), .A2(new_n682), .A3(new_n753), .A4(new_n948), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n944), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(G953), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n831), .A2(new_n760), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n784), .A2(new_n724), .A3(new_n744), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n944), .A2(new_n758), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n661), .B1(new_n954), .B2(new_n260), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n242), .A2(new_n252), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(new_n515), .ZN(new_n957));
  MUX2_X1   g771(.A(new_n951), .B(new_n955), .S(new_n957), .Z(new_n958));
  AOI21_X1  g772(.A(new_n260), .B1(G227), .B2(G900), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT126), .Z(new_n960));
  XNOR2_X1  g774(.A(new_n958), .B(new_n960), .ZN(G72));
  NAND2_X1  g775(.A1(G472), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT63), .Z(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n954), .B2(new_n939), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n309), .A2(new_n272), .ZN(new_n967));
  OAI211_X1 g781(.A(KEYINPUT127), .B(new_n963), .C1(new_n954), .C2(new_n939), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n950), .A2(new_n940), .ZN(new_n970));
  INV_X1    g784(.A(new_n963), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n272), .B(new_n309), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n690), .B2(new_n310), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n868), .A2(new_n973), .ZN(new_n974));
  AND4_X1   g788(.A1(new_n919), .A2(new_n969), .A3(new_n972), .A4(new_n974), .ZN(G57));
endmodule


