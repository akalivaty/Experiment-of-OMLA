//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT95), .A3(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(G143), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G122), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G116), .ZN(new_n197));
  INV_X1    g011(.A(G116), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G122), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n200), .B(G107), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT13), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT96), .B1(new_n192), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT96), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n189), .A2(new_n191), .A3(new_n204), .A4(KEYINPUT13), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n192), .A2(new_n202), .ZN(new_n206));
  AND4_X1   g020(.A1(new_n194), .A2(new_n203), .A3(new_n205), .A4(new_n206), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n195), .B(new_n201), .C1(new_n207), .C2(new_n193), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n200), .A2(G107), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n192), .A2(new_n194), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G134), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n209), .B1(new_n211), .B2(new_n195), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n200), .A2(KEYINPUT14), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT14), .ZN(new_n214));
  OAI21_X1  g028(.A(G107), .B1(new_n199), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT97), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G107), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n196), .A2(G116), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(KEYINPUT14), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT97), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n219), .B(new_n220), .C1(KEYINPUT14), .C2(new_n200), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT98), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n212), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n223), .B1(new_n212), .B2(new_n222), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n208), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT99), .ZN(new_n227));
  XOR2_X1   g041(.A(KEYINPUT9), .B(G234), .Z(new_n228));
  XNOR2_X1  g042(.A(new_n228), .B(KEYINPUT82), .ZN(new_n229));
  INV_X1    g043(.A(G953), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(G217), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT99), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n208), .B(new_n232), .C1(new_n224), .C2(new_n225), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n227), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G902), .ZN(new_n235));
  INV_X1    g049(.A(new_n231), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n226), .A2(KEYINPUT99), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT100), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G478), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(KEYINPUT15), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n234), .A2(KEYINPUT100), .A3(new_n235), .A4(new_n237), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT101), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT101), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n240), .A2(new_n246), .A3(new_n242), .A4(new_n243), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n242), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n234), .A2(new_n235), .A3(new_n249), .A4(new_n237), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT102), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G475), .ZN(new_n254));
  INV_X1    g068(.A(G237), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(new_n230), .A3(G214), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n256), .B(new_n190), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G131), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT17), .ZN(new_n259));
  OR2_X1    g073(.A1(new_n256), .A2(new_n190), .ZN(new_n260));
  INV_X1    g074(.A(G131), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n256), .A2(new_n190), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n258), .A2(new_n259), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G146), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT16), .ZN(new_n266));
  INV_X1    g080(.A(G140), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(G125), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT77), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G125), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n267), .B1(new_n271), .B2(KEYINPUT76), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT76), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(G125), .A3(G140), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n266), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n265), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n268), .B(KEYINPUT77), .ZN(new_n277));
  INV_X1    g091(.A(new_n275), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(new_n278), .A3(G146), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n257), .A2(KEYINPUT17), .A3(G131), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n264), .A2(new_n276), .A3(new_n279), .A4(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n257), .A2(KEYINPUT18), .A3(G131), .ZN(new_n282));
  XNOR2_X1  g096(.A(G125), .B(G140), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n265), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n272), .A2(new_n274), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n284), .B1(new_n285), .B2(new_n265), .ZN(new_n286));
  NAND2_X1  g100(.A1(KEYINPUT18), .A2(G131), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n260), .A2(new_n262), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n282), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n281), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(G113), .B(G122), .ZN(new_n291));
  INV_X1    g105(.A(G104), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n281), .A2(new_n293), .A3(new_n289), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n254), .B1(new_n297), .B2(new_n235), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n258), .A2(new_n263), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT19), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n283), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n301), .B(new_n265), .C1(new_n300), .C2(new_n285), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n279), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(KEYINPUT94), .A3(new_n289), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n294), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT94), .B1(new_n303), .B2(new_n289), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n296), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(G475), .A2(G902), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT20), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT20), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n307), .A2(new_n311), .A3(new_n308), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n298), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n230), .A2(G952), .ZN(new_n314));
  INV_X1    g128(.A(G234), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(new_n255), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  AOI211_X1 g131(.A(new_n235), .B(new_n230), .C1(G234), .C2(G237), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT21), .B(G898), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n313), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G214), .B1(G237), .B2(G902), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G210), .B1(G237), .B2(G902), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  AND2_X1   g141(.A1(KEYINPUT0), .A2(G128), .ZN(new_n328));
  XNOR2_X1  g142(.A(G143), .B(G146), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT64), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n265), .A2(G143), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n190), .A2(G146), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(KEYINPUT0), .A2(G128), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n328), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n336), .A3(KEYINPUT64), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n271), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  OR2_X1    g152(.A1(new_n338), .A2(KEYINPUT91), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n190), .A2(G146), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n265), .A2(G143), .ZN(new_n342));
  OAI211_X1 g156(.A(G128), .B(new_n340), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n332), .B(new_n333), .C1(KEYINPUT1), .C2(new_n188), .ZN(new_n344));
  AOI21_X1  g158(.A(G125), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT91), .B1(new_n338), .B2(new_n345), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n339), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G224), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(G953), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(KEYINPUT92), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n347), .B(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT2), .ZN(new_n352));
  INV_X1    g166(.A(G113), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT66), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT66), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(KEYINPUT2), .B2(G113), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n354), .A2(new_n356), .B1(KEYINPUT2), .B2(G113), .ZN(new_n357));
  XNOR2_X1  g171(.A(G116), .B(G119), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(KEYINPUT5), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n198), .A2(KEYINPUT5), .A3(G119), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(new_n353), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n359), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  AND2_X1   g177(.A1(KEYINPUT84), .A2(G101), .ZN(new_n364));
  NOR2_X1   g178(.A1(KEYINPUT84), .A2(G101), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT3), .B1(new_n292), .B2(G107), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n217), .A3(G104), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n292), .A2(G107), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n366), .A2(new_n367), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n217), .A2(G104), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n370), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n372), .B1(new_n374), .B2(G101), .ZN(new_n375));
  INV_X1    g189(.A(G101), .ZN(new_n376));
  AOI211_X1 g190(.A(KEYINPUT85), .B(new_n376), .C1(new_n373), .C2(new_n370), .ZN(new_n377));
  OAI211_X1 g191(.A(KEYINPUT86), .B(new_n371), .C1(new_n375), .C2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G104), .B(G107), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT85), .B1(new_n380), .B2(new_n376), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n374), .A2(new_n372), .A3(G101), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT86), .B1(new_n383), .B2(new_n371), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n363), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n357), .A2(new_n358), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n359), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G101), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT4), .A3(new_n371), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(new_n391), .A3(G101), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n387), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n385), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(G110), .B(G122), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(KEYINPUT90), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n385), .A2(new_n393), .A3(new_n395), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n394), .A2(KEYINPUT6), .A3(new_n396), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n351), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n395), .B(KEYINPUT8), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n357), .A2(new_n358), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT93), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n360), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n362), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n360), .A2(new_n406), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n383), .A2(new_n371), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT86), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n410), .B1(new_n413), .B2(new_n378), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n363), .B1(new_n371), .B2(new_n383), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n404), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n338), .A2(new_n345), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT7), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n350), .A2(new_n418), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n339), .A2(new_n346), .A3(new_n419), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n416), .A2(new_n398), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n235), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n327), .B1(new_n403), .B2(new_n423), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n347), .A2(new_n350), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n347), .A2(new_n350), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n398), .A2(KEYINPUT6), .B1(new_n394), .B2(new_n396), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n394), .A2(KEYINPUT6), .A3(new_n396), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n425), .B(new_n426), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n398), .A2(new_n420), .A3(new_n421), .ZN(new_n430));
  AOI21_X1  g244(.A(G902), .B1(new_n430), .B2(new_n416), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(new_n326), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n325), .B1(new_n424), .B2(new_n432), .ZN(new_n433));
  AND4_X1   g247(.A1(new_n248), .A2(new_n253), .A3(new_n323), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n230), .A2(G227), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT83), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G140), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT11), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n439), .B1(new_n193), .B2(G137), .ZN(new_n440));
  INV_X1    g254(.A(G137), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT11), .A3(G134), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n193), .A2(G137), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G131), .ZN(new_n445));
  AOI21_X1  g259(.A(G131), .B1(new_n193), .B2(G137), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n440), .A2(new_n446), .A3(new_n442), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n343), .A2(new_n344), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n379), .A2(new_n384), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n371), .A3(new_n383), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n448), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT12), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n343), .A2(new_n344), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n413), .A2(new_n456), .A3(new_n378), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n451), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(KEYINPUT12), .A3(new_n448), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT10), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n392), .A2(new_n331), .A3(new_n337), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n461), .A2(new_n451), .B1(new_n462), .B2(new_n390), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n456), .A2(new_n461), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n379), .B2(new_n384), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n440), .A2(new_n442), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n466), .A2(new_n446), .B1(new_n444), .B2(G131), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n463), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT87), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n463), .A2(new_n465), .A3(new_n470), .A4(new_n467), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n460), .A2(KEYINPUT88), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT88), .B1(new_n460), .B2(new_n472), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n438), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n438), .B1(new_n469), .B2(new_n471), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n463), .A2(new_n465), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n448), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(G902), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G469), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT89), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n438), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT88), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n469), .A2(new_n471), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT12), .B1(new_n458), .B2(new_n448), .ZN(new_n486));
  AOI211_X1 g300(.A(new_n454), .B(new_n467), .C1(new_n457), .C2(new_n451), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n484), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n460), .A2(KEYINPUT88), .A3(new_n472), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n483), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n479), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n235), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT89), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(G469), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n476), .A2(new_n460), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n483), .B1(new_n472), .B2(new_n478), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n481), .B(new_n235), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n482), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G217), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(G234), .B2(new_n235), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(G902), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT81), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT22), .B(G137), .ZN(new_n504));
  INV_X1    g318(.A(G221), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n505), .A2(new_n315), .A3(G953), .ZN(new_n506));
  XOR2_X1   g320(.A(new_n504), .B(new_n506), .Z(new_n507));
  NAND2_X1  g321(.A1(new_n276), .A2(new_n279), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT23), .ZN(new_n509));
  INV_X1    g323(.A(G119), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(G128), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n188), .A2(KEYINPUT23), .A3(G119), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n511), .B(new_n512), .C1(G119), .C2(new_n188), .ZN(new_n513));
  XNOR2_X1  g327(.A(G119), .B(G128), .ZN(new_n514));
  XOR2_X1   g328(.A(KEYINPUT24), .B(G110), .Z(new_n515));
  AOI22_X1  g329(.A1(new_n513), .A2(G110), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  OAI22_X1  g331(.A1(new_n513), .A2(G110), .B1(new_n514), .B2(new_n515), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n279), .A2(new_n518), .A3(new_n284), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT78), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n517), .A2(KEYINPUT78), .A3(new_n519), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n507), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n507), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n517), .B2(new_n519), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n503), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n524), .A2(KEYINPUT81), .A3(new_n527), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n502), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n235), .B1(new_n524), .B2(new_n527), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT79), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(KEYINPUT80), .B2(KEYINPUT25), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n501), .ZN(new_n537));
  OAI211_X1 g351(.A(KEYINPUT79), .B(new_n235), .C1(new_n524), .C2(new_n527), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT25), .B1(new_n538), .B2(KEYINPUT80), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n531), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n541));
  INV_X1    g355(.A(G210), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n542), .A2(G237), .A3(G953), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n541), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT26), .B(G101), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT28), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT67), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n331), .A2(new_n337), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n549), .B1(new_n467), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n448), .A2(KEYINPUT67), .A3(new_n331), .A4(new_n337), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n359), .A2(new_n386), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n440), .A2(new_n446), .A3(new_n442), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n441), .A2(G134), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n261), .B1(new_n556), .B2(new_n443), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT68), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n193), .A2(G137), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n441), .A2(G134), .ZN(new_n560));
  OAI21_X1  g374(.A(G131), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT68), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n447), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n558), .A2(new_n449), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT69), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT69), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n558), .A2(new_n449), .A3(new_n566), .A4(new_n563), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n553), .A2(new_n554), .A3(new_n565), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n561), .A2(new_n447), .ZN(new_n569));
  OAI22_X1  g383(.A1(new_n467), .A2(new_n550), .B1(new_n569), .B2(new_n456), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n387), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n548), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n448), .A2(new_n331), .A3(new_n337), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n564), .A2(new_n573), .A3(new_n554), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n548), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT72), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n574), .A2(KEYINPUT72), .A3(new_n548), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n547), .B1(new_n572), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT73), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n565), .A2(new_n567), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n571), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT28), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n574), .A2(KEYINPUT72), .A3(new_n548), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT72), .B1(new_n574), .B2(new_n548), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(KEYINPUT73), .A3(new_n547), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n582), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n553), .A2(KEYINPUT30), .A3(new_n565), .A4(new_n567), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT65), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n331), .A2(new_n337), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n561), .A2(new_n447), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n595), .A2(new_n448), .B1(new_n449), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n594), .B1(new_n597), .B2(KEYINPUT30), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT30), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n570), .A2(KEYINPUT65), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n593), .A2(new_n601), .A3(new_n387), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT31), .ZN(new_n603));
  INV_X1    g417(.A(new_n583), .ZN(new_n604));
  INV_X1    g418(.A(new_n584), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n547), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n602), .A2(new_n603), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n602), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT31), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT71), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n603), .B1(new_n602), .B2(new_n606), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT71), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n592), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(G472), .A2(G902), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT32), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n586), .A2(new_n589), .A3(new_n546), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT75), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n602), .A2(new_n568), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n547), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT29), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT75), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n586), .A2(new_n589), .A3(new_n624), .A4(new_n546), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n620), .A2(new_n622), .A3(new_n623), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n551), .A2(new_n552), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n387), .B1(new_n583), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n548), .B1(new_n628), .B2(new_n568), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(new_n579), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n547), .A2(new_n623), .ZN(new_n631));
  AOI21_X1  g445(.A(G902), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n614), .A2(new_n618), .B1(new_n633), .B2(G472), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT73), .B1(new_n590), .B2(new_n547), .ZN(new_n635));
  AOI211_X1 g449(.A(new_n581), .B(new_n546), .C1(new_n586), .C2(new_n589), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n613), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n602), .A2(new_n603), .A3(new_n606), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n638), .B1(new_n612), .B2(KEYINPUT71), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n615), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT74), .B(KEYINPUT32), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n540), .B1(new_n634), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n505), .B1(new_n229), .B2(new_n235), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n434), .A2(new_n499), .A3(new_n644), .A4(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(new_n366), .Z(G3));
  INV_X1    g462(.A(new_n498), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n493), .A2(G469), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n649), .B1(new_n650), .B2(KEYINPUT89), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n645), .B1(new_n651), .B2(new_n495), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n241), .A2(G902), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n231), .A2(KEYINPUT104), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n226), .B(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT33), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT33), .B1(new_n234), .B2(new_n237), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n654), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n653), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n313), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n326), .B1(new_n429), .B2(new_n431), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n325), .B1(new_n664), .B2(KEYINPUT103), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n424), .A2(new_n666), .A3(new_n432), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n663), .A2(new_n668), .A3(new_n320), .ZN(new_n669));
  INV_X1    g483(.A(G472), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n614), .B2(new_n235), .ZN(new_n671));
  AOI211_X1 g485(.A(new_n610), .B(new_n603), .C1(new_n602), .C2(new_n606), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n582), .B2(new_n591), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n616), .B1(new_n673), .B2(new_n611), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n671), .A2(new_n674), .A3(new_n540), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n652), .A2(new_n669), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT34), .B(G104), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  AOI21_X1  g492(.A(new_n252), .B1(new_n245), .B2(new_n247), .ZN(new_n679));
  NOR4_X1   g493(.A1(new_n679), .A2(new_n668), .A3(new_n320), .A4(new_n662), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n652), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT35), .B(G107), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G9));
  NAND2_X1  g497(.A1(new_n522), .A2(new_n523), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n526), .A2(KEYINPUT36), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n684), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n502), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n536), .A2(new_n501), .ZN(new_n690));
  INV_X1    g504(.A(new_n539), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n671), .A2(new_n674), .A3(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n434), .A2(new_n499), .A3(new_n646), .A4(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT37), .B(G110), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G12));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n692), .B1(new_n634), .B2(new_n643), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n665), .A2(new_n667), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n499), .A2(new_n698), .A3(new_n646), .A4(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(G900), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n317), .B1(new_n318), .B2(new_n701), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n679), .A2(new_n662), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n697), .B1(new_n700), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n688), .B1(new_n537), .B2(new_n539), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n633), .A2(G472), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n618), .B1(new_n637), .B2(new_n639), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n641), .B1(new_n614), .B2(new_n615), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n706), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n668), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n652), .A2(new_n712), .A3(KEYINPUT105), .A4(new_n703), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G128), .ZN(G30));
  NAND2_X1  g529(.A1(new_n628), .A2(new_n568), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n670), .B1(new_n716), .B2(new_n547), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n717), .A2(new_n608), .B1(G472), .B2(G902), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n718), .B(KEYINPUT106), .Z(new_n719));
  NAND3_X1  g533(.A1(new_n643), .A2(new_n708), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT107), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n424), .A2(new_n432), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n722), .B(KEYINPUT38), .Z(new_n723));
  NAND3_X1  g537(.A1(new_n692), .A2(new_n662), .A3(new_n324), .ZN(new_n724));
  NOR4_X1   g538(.A1(new_n721), .A2(new_n679), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  XOR2_X1   g539(.A(new_n702), .B(KEYINPUT39), .Z(new_n726));
  NAND2_X1  g540(.A1(new_n652), .A2(new_n726), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n727), .A2(KEYINPUT40), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(KEYINPUT40), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n725), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G143), .ZN(G45));
  INV_X1    g545(.A(new_n702), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n661), .A2(new_n662), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n700), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n265), .ZN(G48));
  NAND2_X1  g549(.A1(new_n472), .A2(new_n478), .ZN(new_n736));
  AOI22_X1  g550(.A1(new_n736), .A2(new_n438), .B1(new_n476), .B2(new_n460), .ZN(new_n737));
  OAI21_X1  g551(.A(G469), .B1(new_n737), .B2(G902), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n646), .A3(new_n498), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n644), .A2(new_n669), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT41), .B(G113), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G15));
  NAND3_X1  g557(.A1(new_n680), .A2(new_n644), .A3(new_n740), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G116), .ZN(G18));
  NAND4_X1  g559(.A1(new_n679), .A2(new_n740), .A3(new_n699), .A4(new_n323), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT108), .B1(new_n746), .B2(new_n711), .ZN(new_n747));
  AOI211_X1 g561(.A(new_n322), .B(new_n252), .C1(new_n245), .C2(new_n247), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n668), .A2(new_n739), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n698), .A2(new_n748), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  NOR2_X1   g567(.A1(new_n607), .A2(new_n612), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n547), .B1(new_n629), .B2(new_n579), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n616), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n671), .A2(new_n540), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n665), .A2(new_n667), .A3(new_n662), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n679), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n759), .A3(new_n321), .A4(new_n740), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G122), .ZN(G24));
  NOR3_X1   g575(.A1(new_n733), .A2(new_n668), .A3(new_n739), .ZN(new_n762));
  INV_X1    g576(.A(new_n756), .ZN(new_n763));
  AOI21_X1  g577(.A(G902), .B1(new_n673), .B2(new_n611), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n706), .B(new_n763), .C1(new_n764), .C2(new_n670), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT109), .B1(new_n762), .B2(new_n766), .ZN(new_n767));
  AOI211_X1 g581(.A(new_n702), .B(new_n313), .C1(new_n653), .C2(new_n660), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n740), .A3(new_n699), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n769), .A2(new_n765), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n271), .ZN(G27));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n708), .B(new_n707), .C1(new_n674), .C2(new_n641), .ZN(new_n775));
  INV_X1    g589(.A(new_n540), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n498), .B1(new_n480), .B2(new_n481), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n645), .A2(new_n325), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n424), .A2(new_n432), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n775), .A2(new_n776), .A3(new_n777), .A4(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n774), .B1(new_n781), .B2(new_n733), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n649), .B1(new_n493), .B2(G469), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n783), .A2(new_n733), .A3(new_n779), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n640), .A2(new_n617), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n540), .B1(new_n634), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(KEYINPUT42), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G131), .ZN(G33));
  OR2_X1    g603(.A1(new_n781), .A2(new_n704), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  NAND3_X1  g605(.A1(new_n424), .A2(new_n324), .A3(new_n432), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n640), .B1(new_n764), .B2(new_n670), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n706), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n797));
  XNOR2_X1  g611(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n662), .B1(new_n653), .B2(new_n660), .ZN(new_n799));
  MUX2_X1   g613(.A(new_n797), .B(new_n798), .S(new_n799), .Z(new_n800));
  NAND2_X1  g614(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n792), .B1(new_n802), .B2(KEYINPUT44), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n804), .B1(new_n491), .B2(new_n492), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n475), .A2(KEYINPUT45), .A3(new_n479), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n806), .A3(G469), .ZN(new_n807));
  NAND2_X1  g621(.A1(G469), .A2(G902), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT46), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n649), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(KEYINPUT46), .A3(new_n808), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n645), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n726), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n813), .A2(KEYINPUT110), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(KEYINPUT110), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT44), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n801), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n803), .A2(new_n814), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  XOR2_X1   g632(.A(KEYINPUT113), .B(G137), .Z(new_n819));
  XNOR2_X1  g633(.A(new_n818), .B(new_n819), .ZN(G39));
  XOR2_X1   g634(.A(KEYINPUT114), .B(KEYINPUT47), .Z(new_n821));
  NOR2_X1   g635(.A1(new_n812), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n822), .B1(new_n812), .B2(new_n823), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n775), .A2(new_n733), .A3(new_n776), .A4(new_n792), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G140), .ZN(G42));
  NAND4_X1  g641(.A1(new_n723), .A2(new_n799), .A3(new_n776), .A4(new_n778), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n738), .A2(new_n498), .ZN(new_n829));
  XOR2_X1   g643(.A(new_n829), .B(KEYINPUT115), .Z(new_n830));
  AOI21_X1  g644(.A(new_n828), .B1(new_n830), .B2(KEYINPUT49), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n831), .B(new_n721), .C1(KEYINPUT49), .C2(new_n830), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n792), .A2(new_n662), .A3(new_n702), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n679), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n711), .A2(new_n835), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n652), .A2(new_n836), .B1(new_n766), .B2(new_n784), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n788), .A2(new_n837), .A3(new_n790), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n752), .A2(new_n741), .A3(new_n744), .A4(new_n760), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n647), .A2(new_n694), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n499), .A2(new_n675), .A3(new_n646), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n663), .B1(new_n679), .B2(new_n662), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n433), .A2(new_n321), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT116), .B1(new_n841), .B2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n652), .A2(new_n675), .A3(new_n843), .A4(new_n844), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n647), .A4(new_n694), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n840), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT117), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n840), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  INV_X1    g671(.A(new_n772), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n692), .A2(new_n646), .A3(new_n732), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n720), .A2(new_n759), .A3(new_n777), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n700), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n861), .B1(new_n862), .B2(new_n768), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n857), .A2(new_n714), .A3(new_n858), .A4(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(KEYINPUT118), .B(KEYINPUT52), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n772), .B1(new_n705), .B2(new_n713), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n865), .B1(new_n866), .B2(new_n863), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT53), .B1(new_n856), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n869), .A2(KEYINPUT119), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n857), .B1(new_n866), .B2(new_n863), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n840), .A2(new_n854), .A3(new_n851), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n854), .B1(new_n840), .B2(new_n851), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n869), .A2(KEYINPUT119), .B1(new_n876), .B2(KEYINPUT53), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n833), .B1(new_n870), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  INV_X1    g693(.A(new_n830), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n824), .B1(new_n645), .B2(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n800), .A2(new_n317), .A3(new_n757), .ZN(new_n882));
  INV_X1    g696(.A(new_n792), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n800), .A2(new_n317), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n757), .A2(new_n325), .A3(new_n723), .A4(new_n740), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT50), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n739), .A2(new_n316), .A3(new_n792), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n800), .A2(new_n766), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n721), .A2(new_n776), .A3(new_n890), .ZN(new_n892));
  OR3_X1    g706(.A1(new_n892), .A2(new_n662), .A3(new_n661), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n889), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n879), .B1(new_n885), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n882), .A2(new_n750), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n896), .B(new_n314), .C1(new_n663), .C2(new_n892), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n800), .A2(new_n786), .A3(new_n890), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT48), .Z(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n885), .A2(new_n879), .A3(new_n894), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n714), .A2(new_n858), .A3(new_n863), .ZN(new_n905));
  INV_X1    g719(.A(new_n865), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n866), .A2(new_n857), .A3(new_n863), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n840), .A2(new_n851), .A3(KEYINPUT53), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n904), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n840), .A2(KEYINPUT53), .A3(new_n851), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n868), .A2(new_n912), .A3(KEYINPUT120), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT53), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n875), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(KEYINPUT54), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n878), .A2(new_n903), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(G952), .A2(G953), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n832), .B1(new_n919), .B2(new_n920), .ZN(G75));
  NOR2_X1   g735(.A1(new_n230), .A2(G952), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n917), .A2(G902), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n924), .A2(new_n542), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n427), .A2(new_n428), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n351), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n429), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT55), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n929), .A2(KEYINPUT56), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n923), .B1(new_n925), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n924), .B2(new_n542), .ZN(new_n933));
  AOI22_X1  g747(.A1(new_n911), .A2(new_n913), .B1(new_n875), .B2(new_n915), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(new_n235), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(KEYINPUT121), .A3(G210), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT56), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n933), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n931), .B1(new_n929), .B2(new_n938), .ZN(G51));
  NOR2_X1   g753(.A1(new_n934), .A2(new_n833), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n918), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n808), .B(KEYINPUT57), .ZN(new_n942));
  OAI22_X1  g756(.A1(new_n941), .A2(new_n942), .B1(new_n497), .B2(new_n496), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n924), .A2(new_n807), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n922), .B1(new_n943), .B2(new_n944), .ZN(G54));
  NAND3_X1  g759(.A1(new_n935), .A2(KEYINPUT58), .A3(G475), .ZN(new_n946));
  INV_X1    g760(.A(new_n307), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n948), .A2(new_n949), .A3(new_n922), .ZN(G60));
  NOR2_X1   g764(.A1(new_n658), .A2(new_n659), .ZN(new_n951));
  NAND2_X1  g765(.A1(G478), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT59), .Z(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n918), .B2(new_n940), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n923), .ZN(new_n956));
  INV_X1    g770(.A(new_n953), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n878), .B2(new_n918), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n956), .B1(new_n951), .B2(new_n958), .ZN(G63));
  XNOR2_X1  g773(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n500), .A2(new_n235), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n911), .A2(new_n913), .ZN(new_n963));
  AOI21_X1  g777(.A(KEYINPUT53), .B1(new_n856), .B2(new_n872), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n529), .A2(new_n530), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n922), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  AND4_X1   g782(.A1(KEYINPUT123), .A2(new_n917), .A3(new_n687), .A4(new_n962), .ZN(new_n969));
  INV_X1    g783(.A(new_n962), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n914), .B2(new_n916), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT123), .B1(new_n971), .B2(new_n687), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n968), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n968), .B(KEYINPUT61), .C1(new_n969), .C2(new_n972), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(G66));
  INV_X1    g791(.A(new_n839), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n851), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n230), .ZN(new_n980));
  OAI21_X1  g794(.A(G953), .B1(new_n319), .B2(new_n348), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n926), .B1(G898), .B2(new_n230), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(G69));
  NAND2_X1  g798(.A1(new_n593), .A2(new_n601), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n301), .B1(new_n285), .B2(new_n300), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n230), .A2(G900), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n788), .A2(new_n790), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(new_n824), .B2(new_n825), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n814), .A2(new_n759), .A3(new_n786), .A4(new_n815), .ZN(new_n991));
  AOI211_X1 g805(.A(new_n734), .B(new_n772), .C1(new_n705), .C2(new_n713), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n990), .A2(new_n818), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n988), .B1(new_n993), .B2(new_n230), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT124), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n994), .A2(new_n995), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n987), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(G227), .ZN(new_n999));
  OAI21_X1  g813(.A(G953), .B1(new_n999), .B2(new_n701), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT125), .ZN(new_n1001));
  OR2_X1    g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n992), .A2(new_n730), .ZN(new_n1003));
  OR2_X1    g817(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n843), .A2(new_n644), .A3(new_n883), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n727), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1007), .B1(new_n824), .B2(new_n825), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1004), .A2(new_n818), .A3(new_n1005), .A4(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n987), .A2(G953), .ZN(new_n1010));
  AOI22_X1  g824(.A1(new_n1009), .A2(new_n1010), .B1(new_n1001), .B2(new_n1000), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n998), .A2(new_n1002), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1002), .B1(new_n998), .B2(new_n1011), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1012), .A2(new_n1013), .ZN(G72));
  NAND2_X1  g828(.A1(G472), .A2(G902), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1015), .B(KEYINPUT63), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1017), .B1(new_n1009), .B2(new_n979), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n621), .B(KEYINPUT126), .Z(new_n1019));
  NAND3_X1  g833(.A1(new_n1018), .A2(new_n546), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1017), .B1(new_n993), .B2(new_n979), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1019), .A2(new_n546), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n922), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n870), .A2(new_n877), .ZN(new_n1025));
  OR2_X1    g839(.A1(new_n622), .A2(KEYINPUT127), .ZN(new_n1026));
  AOI22_X1  g840(.A1(new_n622), .A2(KEYINPUT127), .B1(new_n602), .B2(new_n606), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1016), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1024), .B1(new_n1025), .B2(new_n1028), .ZN(G57));
endmodule


