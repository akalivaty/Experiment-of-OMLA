//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1207,
    new_n1208, new_n1209, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT64), .Z(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n210), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n213), .B(new_n218), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G226), .B(G232), .Z(new_n228));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT67), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  XNOR2_X1  g0044(.A(KEYINPUT3), .B(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G1698), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G222), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G223), .A2(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n250));
  OAI211_X1 g0050(.A(new_n249), .B(new_n250), .C1(G77), .C2(new_n245), .ZN(new_n251));
  AND2_X1   g0051(.A1(G1), .A2(G13), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(G274), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G226), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n251), .B(new_n258), .C1(new_n259), .C2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G169), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n207), .A2(G20), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT68), .ZN(new_n266));
  NAND3_X1  g0066(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n267), .A2(new_n216), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G50), .ZN(new_n272));
  INV_X1    g0072(.A(new_n269), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n201), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n208), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G150), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI22_X1  g0079(.A1(new_n275), .A2(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(G20), .B2(new_n204), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n272), .B(new_n274), .C1(new_n268), .C2(new_n281), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n264), .B(new_n282), .C1(G179), .C2(new_n262), .ZN(new_n283));
  XNOR2_X1  g0083(.A(new_n282), .B(KEYINPUT9), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT10), .ZN(new_n285));
  INV_X1    g0085(.A(G190), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n262), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n287), .B1(G200), .B2(new_n262), .ZN(new_n288));
  AND3_X1   g0088(.A1(new_n284), .A2(new_n285), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n285), .B1(new_n284), .B2(new_n288), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n283), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n275), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(new_n269), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(new_n271), .B2(new_n292), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n202), .A2(new_n203), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G58), .A2(G68), .ZN(new_n297));
  OAI21_X1  g0097(.A(G20), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G159), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(new_n279), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT3), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(G33), .ZN(new_n302));
  INV_X1    g0102(.A(G33), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(KEYINPUT3), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n208), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n203), .B1(new_n305), .B2(KEYINPUT7), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(KEYINPUT3), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n301), .A2(G33), .ZN(new_n308));
  AOI21_X1  g0108(.A(G20), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n310));
  NOR2_X1   g0110(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n300), .B1(new_n306), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n268), .B1(new_n314), .B2(KEYINPUT16), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT16), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT75), .B1(new_n301), .B2(G33), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT75), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(new_n303), .A3(KEYINPUT3), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n319), .A3(new_n308), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT7), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(G20), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n312), .B1(new_n245), .B2(G20), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n203), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n316), .B1(new_n325), .B2(new_n300), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n295), .B1(new_n315), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G232), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n258), .B1(new_n261), .B2(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(G223), .A2(G1698), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n259), .A2(G1698), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n307), .A2(new_n330), .A3(new_n308), .A4(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G33), .A2(G87), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n254), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(new_n263), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n329), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT18), .B1(new_n327), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n323), .A2(new_n324), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G68), .ZN(new_n342));
  XNOR2_X1  g0142(.A(G58), .B(G68), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n343), .A2(G20), .B1(G159), .B2(new_n278), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT16), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(G68), .B1(new_n309), .B2(new_n321), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n307), .A2(new_n308), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n347), .A2(new_n312), .A3(new_n208), .ZN(new_n348));
  OAI211_X1 g0148(.A(KEYINPUT16), .B(new_n344), .C1(new_n346), .C2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n268), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n294), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n336), .A2(new_n338), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT18), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(KEYINPUT76), .A2(KEYINPUT17), .ZN(new_n356));
  INV_X1    g0156(.A(G200), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n335), .A2(new_n357), .ZN(new_n358));
  NOR3_X1   g0158(.A1(new_n329), .A2(new_n334), .A3(new_n286), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n356), .B1(new_n327), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n326), .A2(new_n350), .A3(new_n349), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n363));
  AND4_X1   g0163(.A1(new_n362), .A2(new_n360), .A3(new_n294), .A4(new_n363), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n340), .B(new_n355), .C1(new_n361), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G238), .A2(G1698), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n245), .B(new_n366), .C1(new_n328), .C2(G1698), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n367), .B(new_n250), .C1(G107), .C2(new_n245), .ZN(new_n368));
  INV_X1    g0168(.A(new_n261), .ZN(new_n369));
  INV_X1    g0169(.A(G274), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n252), .B2(new_n253), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n369), .A2(G244), .B1(new_n257), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT69), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n368), .A2(new_n372), .A3(KEYINPUT69), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(new_n357), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n286), .B1(new_n375), .B2(new_n376), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g0180(.A(KEYINPUT15), .B(G87), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n276), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n382), .A2(new_n383), .B1(G20), .B2(G77), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n292), .A2(new_n278), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n268), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G77), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n273), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT70), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n271), .A2(G77), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n389), .B1(new_n388), .B2(new_n390), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n380), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n377), .A2(new_n337), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n375), .A2(new_n263), .A3(new_n376), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n388), .A2(new_n390), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n291), .A2(new_n365), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT12), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n271), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n203), .A2(G20), .ZN(new_n403));
  OAI221_X1 g0203(.A(new_n403), .B1(new_n276), .B2(new_n387), .C1(new_n279), .C2(new_n201), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(KEYINPUT11), .A3(new_n350), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n350), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT11), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G13), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n401), .A2(new_n409), .A3(G1), .ZN(new_n410));
  INV_X1    g0210(.A(new_n403), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n410), .A2(new_n411), .B1(new_n401), .B2(new_n269), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n402), .A2(new_n405), .A3(new_n408), .A4(new_n412), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT73), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT14), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n254), .A2(G238), .A3(new_n260), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n258), .A2(new_n416), .A3(KEYINPUT72), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT72), .B1(new_n258), .B2(new_n416), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n259), .A2(new_n246), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n328), .A2(G1698), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n307), .A2(new_n420), .A3(new_n308), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G97), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT71), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT71), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n422), .A2(new_n426), .A3(new_n423), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n427), .A3(new_n250), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n419), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n429), .B1(new_n419), .B2(new_n428), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n415), .B(G169), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n419), .A2(new_n428), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT13), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(G179), .A3(new_n430), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n430), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n415), .B1(new_n438), .B2(G169), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n414), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  XOR2_X1   g0240(.A(new_n413), .B(KEYINPUT73), .Z(new_n441));
  NAND3_X1  g0241(.A1(new_n435), .A2(G190), .A3(new_n430), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n438), .A2(G200), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n400), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT21), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n255), .A2(KEYINPUT5), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n207), .B(G45), .C1(new_n255), .C2(KEYINPUT5), .ZN(new_n451));
  OAI211_X1 g0251(.A(G270), .B(new_n254), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n451), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n453), .A2(new_n371), .A3(new_n449), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT79), .B(G303), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n250), .B1(new_n245), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G264), .A2(G1698), .ZN(new_n457));
  INV_X1    g0257(.A(G257), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n457), .B1(new_n458), .B2(G1698), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n347), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n452), .B(new_n454), .C1(new_n456), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G169), .ZN(new_n462));
  INV_X1    g0262(.A(G116), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n273), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n207), .A2(G33), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n269), .A2(new_n465), .A3(new_n216), .A4(new_n267), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n464), .B1(new_n466), .B2(new_n463), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n267), .A2(new_n216), .B1(G20), .B2(new_n463), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  INV_X1    g0269(.A(G97), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n469), .B(new_n208), .C1(G33), .C2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT20), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n468), .A2(KEYINPUT20), .A3(new_n471), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n448), .B1(new_n462), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n466), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G116), .ZN(new_n478));
  INV_X1    g0278(.A(new_n474), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n478), .B(new_n464), .C1(new_n479), .C2(new_n472), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n480), .A2(KEYINPUT21), .A3(G169), .A4(new_n461), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n461), .A2(new_n337), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n480), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n476), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n461), .A2(new_n286), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n480), .B1(G200), .B2(new_n461), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n307), .A2(new_n308), .A3(new_n208), .A4(G87), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT22), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT22), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n245), .A2(new_n490), .A3(new_n208), .A4(G87), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT24), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT23), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n208), .B2(G107), .ZN(new_n495));
  INV_X1    g0295(.A(G107), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(KEYINPUT23), .A3(G20), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n383), .A2(G116), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n492), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n493), .B1(new_n492), .B2(new_n498), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n350), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OR3_X1    g0301(.A1(new_n269), .A2(KEYINPUT80), .A3(G107), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT80), .B1(new_n269), .B2(G107), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT25), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT25), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n502), .A2(new_n506), .A3(new_n503), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n505), .A2(new_n507), .B1(G107), .B2(new_n477), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n501), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n307), .A2(new_n308), .A3(G250), .A4(new_n246), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G294), .ZN(new_n511));
  AND2_X1   g0311(.A1(G257), .A2(G1698), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n307), .A2(new_n308), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n250), .ZN(new_n515));
  OAI211_X1 g0315(.A(G264), .B(new_n254), .C1(new_n450), .C2(new_n451), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n454), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n263), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n515), .A2(new_n337), .A3(new_n454), .A4(new_n516), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n509), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n516), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n250), .B2(new_n514), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(G190), .A3(new_n454), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n517), .A2(G200), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n501), .A2(new_n524), .A3(new_n508), .A4(new_n525), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n381), .A2(new_n273), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n307), .A2(new_n308), .A3(new_n208), .A4(G68), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT19), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n276), .B2(new_n470), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n208), .B1(new_n423), .B2(new_n530), .ZN(new_n533));
  INV_X1    g0333(.A(G87), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(new_n470), .A3(new_n496), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT78), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n533), .A2(KEYINPUT78), .A3(new_n535), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n532), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n528), .B1(new_n540), .B2(new_n268), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n466), .A2(new_n534), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n207), .A2(new_n370), .A3(G45), .ZN(new_n544));
  INV_X1    g0344(.A(G250), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n256), .B2(G1), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n254), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(G238), .A2(G1698), .ZN(new_n548));
  INV_X1    g0348(.A(G244), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(G1698), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(new_n245), .B1(G33), .B2(G116), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n547), .B1(new_n551), .B2(new_n254), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G200), .ZN(new_n553));
  OAI211_X1 g0353(.A(G190), .B(new_n547), .C1(new_n551), .C2(new_n254), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n263), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n337), .B(new_n547), .C1(new_n551), .C2(new_n254), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI221_X1 g0358(.A(new_n528), .B1(new_n381), .B2(new_n466), .C1(new_n540), .C2(new_n268), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n543), .A2(new_n555), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(G257), .B(new_n254), .C1(new_n450), .C2(new_n451), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n454), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(KEYINPUT77), .A2(KEYINPUT4), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n549), .A2(G1698), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n563), .B1(new_n347), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n245), .B(new_n564), .C1(KEYINPUT77), .C2(KEYINPUT4), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n245), .A2(G250), .A3(G1698), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n469), .A4(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n562), .B1(new_n569), .B2(new_n250), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n263), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT6), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n573), .A2(new_n470), .A3(G107), .ZN(new_n574));
  XNOR2_X1  g0374(.A(G97), .B(G107), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n574), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n576), .A2(new_n208), .B1(new_n387), .B2(new_n279), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n496), .B1(new_n323), .B2(new_n324), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n350), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n273), .A2(new_n470), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n466), .B2(new_n470), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n570), .A2(new_n337), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n572), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n341), .A2(G107), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n575), .A2(new_n573), .ZN(new_n587));
  INV_X1    g0387(.A(new_n574), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n589), .A2(G20), .B1(G77), .B2(new_n278), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n581), .B1(new_n591), .B2(new_n350), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n570), .A2(G190), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n592), .B(new_n593), .C1(new_n357), .C2(new_n570), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n560), .A2(new_n585), .A3(new_n594), .ZN(new_n595));
  AND4_X1   g0395(.A1(new_n447), .A2(new_n487), .A3(new_n527), .A4(new_n595), .ZN(G372));
  NAND3_X1  g0396(.A1(new_n360), .A2(new_n362), .A3(new_n294), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(KEYINPUT76), .B2(KEYINPUT17), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n327), .A2(new_n363), .A3(new_n360), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n398), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n444), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n601), .B1(new_n603), .B2(new_n440), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT82), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n327), .A2(KEYINPUT18), .A3(new_n339), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n354), .B1(new_n352), .B2(new_n353), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n340), .A2(KEYINPUT82), .A3(new_n355), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  OAI22_X1  g0411(.A1(new_n604), .A2(new_n611), .B1(new_n290), .B2(new_n289), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n283), .ZN(new_n613));
  XNOR2_X1  g0413(.A(new_n613), .B(KEYINPUT83), .ZN(new_n614));
  INV_X1    g0414(.A(new_n585), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n543), .A2(new_n555), .ZN(new_n616));
  XOR2_X1   g0416(.A(KEYINPUT81), .B(KEYINPUT26), .Z(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n594), .A2(new_n616), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n476), .A2(new_n481), .A3(new_n483), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n501), .A2(new_n508), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n524), .A2(new_n525), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n521), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n621), .B1(new_n625), .B2(new_n615), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n619), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n558), .A2(new_n559), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n614), .B1(new_n446), .B2(new_n631), .ZN(G369));
  NAND3_X1  g0432(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(G213), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G343), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(new_n475), .ZN(new_n640));
  MUX2_X1   g0440(.A(new_n487), .B(new_n484), .S(new_n640), .Z(new_n641));
  AND2_X1   g0441(.A1(new_n641), .A2(G330), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n527), .B1(new_n623), .B2(new_n639), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n521), .B2(new_n639), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n518), .A2(new_n519), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n501), .B2(new_n508), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n639), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n622), .A2(new_n638), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n527), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n645), .A2(new_n648), .A3(new_n650), .ZN(G399));
  NOR2_X1   g0451(.A1(new_n631), .A2(new_n638), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT29), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n615), .A2(KEYINPUT26), .A3(new_n616), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n526), .B1(new_n647), .B2(new_n484), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n620), .B1(new_n656), .B2(new_n585), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n655), .B1(new_n657), .B2(new_n618), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n638), .B1(new_n658), .B2(new_n629), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(new_n653), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n595), .A2(new_n527), .A3(new_n487), .A4(new_n639), .ZN(new_n661));
  INV_X1    g0461(.A(new_n552), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n570), .A2(new_n482), .A3(new_n523), .A4(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT30), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n662), .A2(new_n523), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n666), .A2(new_n570), .A3(KEYINPUT30), .A4(new_n482), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n517), .A2(new_n337), .A3(new_n461), .A4(new_n552), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n570), .ZN(new_n670));
  OAI211_X1 g0470(.A(KEYINPUT31), .B(new_n638), .C1(new_n668), .C2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT85), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT84), .B1(new_n669), .B2(new_n570), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n552), .A2(new_n461), .A3(new_n337), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT84), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n571), .A2(new_n674), .A3(new_n675), .A4(new_n517), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n665), .A2(new_n667), .A3(new_n673), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n638), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT31), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n672), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  AOI211_X1 g0480(.A(KEYINPUT85), .B(KEYINPUT31), .C1(new_n677), .C2(new_n638), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n661), .B(new_n671), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n654), .A2(new_n660), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n207), .ZN(new_n686));
  INV_X1    g0486(.A(new_n211), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G41), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n535), .A2(G116), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G1), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n214), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n686), .A2(new_n693), .ZN(G364));
  NOR2_X1   g0494(.A1(G13), .A2(G33), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G20), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n641), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n216), .B1(G20), .B2(new_n263), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G190), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n702), .A2(new_n286), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n704), .A2(new_n203), .B1(new_n706), .B2(new_n201), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n208), .A2(new_n286), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(new_n337), .A3(G200), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n208), .A2(G190), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n337), .A2(G200), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n710), .A2(G87), .B1(new_n714), .B2(G77), .ZN(new_n715));
  INV_X1    g0515(.A(new_n711), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n716), .A2(G179), .A3(new_n357), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n715), .B(new_n245), .C1(new_n496), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n708), .A2(new_n712), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT89), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n720), .A2(new_n721), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI211_X1 g0526(.A(new_n707), .B(new_n719), .C1(G58), .C2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n337), .A2(new_n357), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT90), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n716), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n299), .ZN(new_n732));
  XOR2_X1   g0532(.A(KEYINPUT91), .B(KEYINPUT32), .Z(new_n733));
  OAI21_X1  g0533(.A(G20), .B1(new_n729), .B2(new_n286), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n732), .A2(new_n733), .B1(G97), .B2(new_n734), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n727), .B(new_n735), .C1(new_n732), .C2(new_n733), .ZN(new_n736));
  INV_X1    g0536(.A(G326), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n706), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G283), .ZN(new_n739));
  INV_X1    g0539(.A(G311), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n718), .A2(new_n739), .B1(new_n713), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(KEYINPUT33), .B(G317), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n738), .B(new_n741), .C1(new_n703), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n734), .A2(G294), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n726), .A2(G322), .B1(new_n730), .B2(G329), .ZN(new_n745));
  INV_X1    g0545(.A(G303), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n347), .B1(new_n709), .B2(new_n746), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT92), .Z(new_n748));
  NAND4_X1  g0548(.A1(new_n743), .A2(new_n744), .A3(new_n745), .A4(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n701), .B1(new_n736), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n409), .A2(G20), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G45), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n689), .A2(G1), .A3(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n211), .A2(new_n245), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n755), .B(KEYINPUT86), .Z(new_n756));
  XOR2_X1   g0556(.A(G355), .B(KEYINPUT87), .Z(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(G116), .B2(new_n211), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n687), .A2(new_n245), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(new_n215), .B2(new_n256), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT88), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n763), .A2(KEYINPUT88), .B1(G45), .B2(new_n240), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n759), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n697), .A2(new_n700), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n754), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n699), .A2(new_n750), .A3(new_n769), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n641), .A2(G330), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n642), .A2(new_n754), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(G396));
  NOR2_X1   g0574(.A1(new_n398), .A2(new_n638), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n397), .A2(new_n638), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n394), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n775), .B1(new_n777), .B2(new_n398), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n652), .B(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n754), .B1(new_n779), .B2(new_n684), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n684), .B2(new_n779), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n700), .A2(new_n695), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n754), .B1(G77), .B2(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n730), .A2(G311), .B1(G87), .B2(new_n717), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT93), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n347), .B1(new_n713), .B2(new_n463), .C1(new_n709), .C2(new_n496), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n704), .A2(new_n739), .B1(new_n706), .B2(new_n746), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n787), .B(new_n788), .C1(new_n726), .C2(G294), .ZN(new_n789));
  INV_X1    g0589(.A(new_n734), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n786), .B(new_n789), .C1(new_n470), .C2(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n714), .A2(G159), .B1(G150), .B2(new_n703), .ZN(new_n792));
  INV_X1    g0592(.A(G137), .ZN(new_n793));
  INV_X1    g0593(.A(G143), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n792), .B1(new_n793), .B2(new_n706), .C1(new_n725), .C2(new_n794), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT34), .Z(new_n796));
  OAI22_X1  g0596(.A1(new_n718), .A2(new_n203), .B1(new_n201), .B2(new_n709), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT94), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n347), .B1(new_n730), .B2(G132), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(new_n202), .C2(new_n790), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n791), .B1(new_n796), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n784), .B1(new_n801), .B2(new_n700), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n778), .B2(new_n696), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT95), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n781), .A2(new_n804), .ZN(G384));
  OR2_X1    g0605(.A1(new_n589), .A2(KEYINPUT35), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n589), .A2(KEYINPUT35), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n806), .A2(G116), .A3(new_n217), .A4(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT96), .B(KEYINPUT36), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n296), .A2(new_n214), .A3(new_n387), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT97), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n812), .A2(KEYINPUT97), .B1(new_n201), .B2(G68), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n207), .B(G13), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT101), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT99), .ZN(new_n818));
  OR3_X1    g0618(.A1(new_n440), .A2(new_n818), .A3(new_n638), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n440), .B2(new_n638), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT39), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT38), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT37), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n352), .A2(new_n353), .ZN(new_n826));
  INV_X1    g0626(.A(new_n636), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n352), .A2(new_n827), .ZN(new_n828));
  AND4_X1   g0628(.A1(new_n825), .A2(new_n826), .A3(new_n828), .A4(new_n597), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n344), .B1(new_n346), .B2(new_n348), .ZN(new_n830));
  AOI21_X1  g0630(.A(KEYINPUT16), .B1(new_n830), .B2(KEYINPUT98), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT98), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n832), .B(new_n344), .C1(new_n346), .C2(new_n348), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n351), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n827), .B1(new_n834), .B2(new_n295), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n831), .A2(new_n833), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n295), .B1(new_n836), .B2(new_n315), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n835), .B(new_n597), .C1(new_n339), .C2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n829), .B1(KEYINPUT37), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n606), .A2(new_n607), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n835), .B1(new_n840), .B2(new_n600), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n824), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n597), .B1(new_n837), .B2(new_n636), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n837), .A2(new_n339), .ZN(new_n844));
  OAI21_X1  g0644(.A(KEYINPUT37), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n826), .A2(new_n828), .A3(new_n825), .A4(new_n597), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n835), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n365), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n847), .A2(new_n849), .A3(KEYINPUT38), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n823), .B1(new_n842), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n828), .B1(new_n610), .B2(new_n600), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n826), .A2(new_n828), .A3(new_n597), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT37), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n846), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n824), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n845), .A2(new_n846), .B1(new_n365), .B2(new_n848), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT39), .B1(new_n858), .B2(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT100), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n851), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n857), .A2(new_n859), .A3(KEYINPUT100), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n822), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n639), .B(new_n778), .C1(new_n628), .C2(new_n630), .ZN(new_n865));
  INV_X1    g0665(.A(new_n775), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n842), .A2(new_n850), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n414), .A2(new_n638), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n440), .A2(new_n444), .A3(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n414), .B(new_n638), .C1(new_n437), .C2(new_n439), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n867), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n611), .A2(new_n636), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n817), .B1(new_n864), .B2(new_n875), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n340), .A2(KEYINPUT82), .A3(new_n355), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT82), .B1(new_n340), .B2(new_n355), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n600), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n828), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n881), .B2(new_n855), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n850), .A2(new_n823), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n861), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n868), .A2(KEYINPUT39), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(new_n863), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n821), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n865), .A2(new_n866), .B1(new_n870), .B2(new_n871), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n888), .A2(new_n868), .B1(new_n611), .B2(new_n636), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n887), .A2(KEYINPUT101), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n876), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n654), .A2(new_n660), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n447), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n614), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n891), .B(new_n894), .Z(new_n895));
  NAND3_X1  g0695(.A1(new_n677), .A2(KEYINPUT31), .A3(new_n638), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n678), .A2(new_n679), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n661), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n380), .A2(new_n393), .B1(new_n397), .B2(new_n638), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n866), .B1(new_n899), .B2(new_n602), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n870), .B2(new_n871), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n868), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n857), .A2(new_n850), .ZN(new_n904));
  AND4_X1   g0704(.A1(KEYINPUT40), .A2(new_n872), .A3(new_n898), .A4(new_n778), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n902), .A2(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(new_n447), .A3(new_n898), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(G330), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n906), .B1(new_n447), .B2(new_n898), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n895), .A2(new_n910), .B1(new_n207), .B2(new_n751), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT102), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n895), .A2(new_n910), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n911), .A2(KEYINPUT102), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n816), .B1(new_n914), .B2(new_n915), .ZN(G367));
  NAND2_X1  g0716(.A1(new_n760), .A2(new_n236), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n768), .B1(new_n687), .B2(new_n382), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n753), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n543), .A2(new_n639), .ZN(new_n920));
  MUX2_X1   g0720(.A(new_n560), .B(new_n630), .S(new_n920), .Z(new_n921));
  OAI221_X1 g0721(.A(new_n347), .B1(new_n739), .B2(new_n713), .C1(new_n718), .C2(new_n470), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(G317), .B2(new_n730), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT46), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n709), .A2(new_n924), .A3(new_n463), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n924), .B1(new_n709), .B2(new_n463), .ZN(new_n926));
  INV_X1    g0726(.A(G294), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n926), .B1(new_n704), .B2(new_n927), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n925), .B(new_n928), .C1(G311), .C2(new_n705), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n726), .A2(new_n455), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n734), .A2(G107), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n923), .A2(new_n929), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n726), .A2(G150), .B1(new_n730), .B2(G137), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n347), .B1(new_n714), .B2(G50), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n717), .A2(G77), .B1(new_n710), .B2(G58), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n703), .A2(G159), .B1(new_n705), .B2(G143), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n933), .A2(new_n934), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n790), .A2(new_n203), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT47), .Z(new_n940));
  OAI221_X1 g0740(.A(new_n919), .B1(new_n698), .B2(new_n921), .C1(new_n940), .C2(new_n701), .ZN(new_n941));
  INV_X1    g0741(.A(new_n645), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n594), .B(new_n585), .C1(new_n592), .C2(new_n639), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n615), .A2(new_n638), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT103), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n921), .A2(KEYINPUT43), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n948), .B(new_n949), .Z(new_n950));
  NOR2_X1   g0750(.A1(new_n945), .A2(new_n650), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n952), .A2(KEYINPUT42), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n585), .B1(new_n943), .B2(new_n521), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n952), .A2(KEYINPUT42), .B1(new_n639), .B2(new_n954), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n953), .A2(new_n955), .B1(KEYINPUT43), .B2(new_n921), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n950), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n752), .A2(G1), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n892), .A2(new_n683), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n650), .A2(new_n648), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n945), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT44), .Z(new_n962));
  NOR2_X1   g0762(.A1(new_n960), .A2(new_n945), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT45), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(new_n942), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n650), .B1(new_n644), .B2(new_n649), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(new_n642), .Z(new_n968));
  OAI21_X1  g0768(.A(new_n959), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n688), .B(KEYINPUT41), .Z(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n958), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n941), .B1(new_n957), .B2(new_n972), .ZN(G387));
  OR2_X1    g0773(.A1(new_n685), .A2(new_n968), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n685), .A2(new_n968), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n974), .A2(new_n688), .A3(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n958), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n644), .A2(new_n698), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n761), .B1(new_n232), .B2(G45), .ZN(new_n979));
  INV_X1    g0779(.A(new_n690), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n979), .B1(new_n980), .B2(new_n756), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n292), .A2(new_n201), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT50), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n256), .B1(new_n203), .B2(new_n387), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n983), .A2(new_n980), .A3(new_n984), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n981), .A2(new_n985), .B1(G107), .B2(new_n211), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n753), .B1(new_n986), .B2(new_n767), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n734), .A2(new_n382), .ZN(new_n988));
  XOR2_X1   g0788(.A(KEYINPUT104), .B(G150), .Z(new_n989));
  AOI22_X1  g0789(.A1(new_n726), .A2(G50), .B1(new_n730), .B2(new_n989), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n709), .A2(new_n387), .B1(new_n713), .B2(new_n203), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n347), .B(new_n991), .C1(G97), .C2(new_n717), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n292), .A2(new_n703), .B1(G159), .B2(new_n705), .ZN(new_n993));
  AND4_X1   g0793(.A1(new_n988), .A2(new_n990), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n705), .A2(G322), .ZN(new_n995));
  INV_X1    g0795(.A(new_n455), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n995), .B1(new_n704), .B2(new_n740), .C1(new_n996), .C2(new_n713), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n726), .B2(G317), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT48), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n734), .A2(G283), .B1(G294), .B2(new_n710), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT105), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(KEYINPUT49), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n347), .B1(new_n463), .B2(new_n718), .C1(new_n731), .C2(new_n737), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n1002), .B2(KEYINPUT49), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n994), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n987), .B1(new_n1006), .B2(new_n701), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n976), .B1(new_n977), .B2(new_n968), .C1(new_n978), .C2(new_n1007), .ZN(G393));
  OAI221_X1 g0808(.A(new_n767), .B1(new_n470), .B2(new_n211), .C1(new_n761), .C2(new_n243), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n754), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n725), .A2(new_n299), .B1(new_n277), .B2(new_n706), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT51), .Z(new_n1012));
  NOR2_X1   g0812(.A1(new_n790), .A2(new_n387), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n709), .A2(new_n203), .B1(new_n713), .B2(new_n275), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n347), .B(new_n1014), .C1(G87), .C2(new_n717), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n201), .B2(new_n704), .C1(new_n794), .C2(new_n731), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n1012), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1017), .A2(KEYINPUT106), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(KEYINPUT106), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n347), .B1(new_n739), .B2(new_n709), .C1(new_n718), .C2(new_n496), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G322), .B2(new_n730), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT107), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n726), .A2(G311), .B1(G317), .B2(new_n705), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT52), .Z(new_n1024));
  OAI22_X1  g0824(.A1(new_n996), .A2(new_n704), .B1(new_n927), .B2(new_n713), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n734), .B2(G116), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1022), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1018), .A2(new_n1019), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1010), .B1(new_n1028), .B2(new_n700), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n698), .B2(new_n946), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n966), .B2(new_n977), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n688), .B1(new_n966), .B2(new_n974), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n966), .A2(new_n974), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1031), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(G390));
  AND3_X1   g0836(.A1(new_n447), .A2(G330), .A3(new_n898), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n894), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n777), .A2(new_n398), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n775), .B1(new_n659), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n682), .A2(G330), .A3(new_n778), .A4(new_n872), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n872), .A2(KEYINPUT108), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT108), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n870), .A2(new_n871), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT110), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n898), .A2(new_n778), .A3(G330), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1047), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1042), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n872), .B1(new_n683), .B2(new_n778), .ZN(new_n1053));
  AND4_X1   g0853(.A1(G330), .A2(new_n872), .A3(new_n898), .A4(new_n778), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n867), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1038), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n822), .B(new_n904), .C1(new_n1040), .C2(new_n1046), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n821), .B1(new_n867), .B2(new_n872), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1058), .B1(new_n886), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT109), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1054), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1054), .A2(KEYINPUT109), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1064), .A2(new_n683), .A3(new_n778), .A4(new_n872), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1065), .B(new_n1058), .C1(new_n886), .C2(new_n1059), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n689), .B1(new_n1057), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1057), .B2(new_n1067), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1063), .A2(new_n958), .A3(new_n1066), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n754), .B1(new_n292), .B2(new_n783), .ZN(new_n1071));
  INV_X1    g0871(.A(G128), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n704), .A2(new_n793), .B1(new_n706), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n245), .B1(new_n718), .B2(new_n201), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(KEYINPUT54), .B(G143), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1073), .B(new_n1074), .C1(new_n714), .C2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n710), .A2(new_n989), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT53), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G125), .B2(new_n730), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n726), .A2(G132), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n734), .A2(G159), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1077), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n726), .A2(G116), .B1(new_n730), .B2(G294), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n245), .B1(new_n710), .B2(G87), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n717), .A2(G68), .B1(new_n714), .B2(G97), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n703), .A2(G107), .B1(new_n705), .B2(G283), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1083), .B1(new_n1013), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1071), .B1(new_n1089), .B2(new_n700), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n886), .B2(new_n696), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT111), .Z(new_n1092));
  NAND3_X1  g0892(.A1(new_n1069), .A2(new_n1070), .A3(new_n1092), .ZN(G378));
  NAND2_X1  g0893(.A1(new_n282), .A2(new_n827), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT55), .Z(new_n1095));
  NAND2_X1  g0895(.A1(new_n291), .A2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(KEYINPUT112), .B(KEYINPUT56), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1095), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1098), .B(new_n283), .C1(new_n290), .C2(new_n289), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1097), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n906), .B2(G330), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n839), .A2(new_n841), .A3(new_n824), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT38), .B1(new_n847), .B2(new_n849), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n872), .A2(new_n898), .A3(new_n778), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n903), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n904), .A2(new_n905), .ZN(new_n1109));
  AND4_X1   g0909(.A1(G330), .A2(new_n1108), .A3(new_n1109), .A4(new_n1102), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1103), .A2(new_n1110), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n864), .A2(new_n817), .A3(new_n875), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT101), .B1(new_n887), .B2(new_n889), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1108), .A2(new_n1109), .A3(G330), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1102), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n906), .A2(G330), .A3(new_n1102), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n876), .A2(new_n1119), .A3(new_n890), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1114), .A2(KEYINPUT113), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT113), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n891), .A2(new_n1122), .A3(new_n1111), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1063), .A2(new_n1056), .A3(new_n1066), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n1038), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(KEYINPUT115), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT115), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1125), .A2(new_n1128), .A3(new_n1038), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT57), .B1(new_n1124), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n688), .B1(new_n1131), .B2(KEYINPUT117), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT57), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1125), .A2(new_n1128), .A3(new_n1038), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1128), .B1(new_n1125), .B2(new_n1038), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1137));
  OAI211_X1 g0937(.A(KEYINPUT117), .B(new_n1133), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT116), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1133), .B1(new_n1114), .B2(new_n1120), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1139), .B1(new_n1130), .B2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1140), .B(new_n1139), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1138), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1132), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1121), .A2(new_n958), .A3(new_n1123), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n726), .A2(G107), .B1(new_n730), .B2(G283), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n718), .A2(new_n202), .B1(new_n381), .B2(new_n713), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n255), .B(new_n347), .C1(new_n709), .C2(new_n387), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n704), .A2(new_n470), .B1(new_n706), .B2(new_n463), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1147), .B(new_n1151), .C1(new_n203), .C2(new_n790), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT58), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n255), .B1(new_n301), .B2(new_n303), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1152), .A2(new_n1153), .B1(new_n201), .B2(new_n1154), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n705), .A2(G125), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n709), .A2(new_n1075), .B1(new_n713), .B2(new_n793), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(G132), .C2(new_n703), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1158), .B1(new_n1072), .B2(new_n725), .C1(new_n277), .C2(new_n790), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n303), .B(new_n255), .C1(new_n718), .C2(new_n299), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G124), .B2(new_n730), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1155), .B1(new_n1153), .B2(new_n1152), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n700), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n753), .B1(new_n201), .B2(new_n782), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(new_n1102), .C2(new_n696), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1146), .A2(KEYINPUT114), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT114), .B1(new_n1146), .B2(new_n1168), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1145), .A2(new_n1171), .ZN(G375));
  OAI211_X1 g0972(.A(new_n1055), .B(new_n1052), .C1(new_n894), .C2(new_n1037), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1057), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n971), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT118), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1056), .A2(new_n958), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1177), .A2(KEYINPUT119), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1177), .A2(KEYINPUT119), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n753), .B1(new_n203), .B2(new_n782), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n726), .A2(G283), .B1(new_n730), .B2(G303), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n709), .A2(new_n470), .B1(new_n713), .B2(new_n496), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n245), .B(new_n1182), .C1(G77), .C2(new_n717), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n703), .A2(G116), .B1(new_n705), .B2(G294), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1181), .A2(new_n988), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1185), .A2(KEYINPUT120), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n709), .A2(new_n299), .B1(new_n713), .B2(new_n277), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n245), .B1(new_n718), .B2(new_n202), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(new_n703), .C2(new_n1076), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n726), .A2(G137), .B1(new_n730), .B2(G128), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n705), .A2(G132), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT121), .Z(new_n1192));
  NAND2_X1  g0992(.A1(new_n734), .A2(G50), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1185), .A2(KEYINPUT120), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1186), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1180), .B1(new_n1196), .B2(new_n701), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1046), .B2(new_n695), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1178), .A2(new_n1179), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1176), .A2(new_n1199), .ZN(G381));
  OR2_X1    g1000(.A1(G387), .A2(G390), .ZN(new_n1201));
  OR3_X1    g1001(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(G381), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT122), .Z(new_n1204));
  NOR2_X1   g1004(.A1(G375), .A2(G378), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(G407));
  NAND2_X1  g1006(.A1(new_n637), .A2(G213), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(G407), .A2(new_n1209), .A3(G213), .ZN(G409));
  XOR2_X1   g1010(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1211));
  OAI211_X1 g1011(.A(G378), .B(new_n1171), .C1(new_n1132), .C2(new_n1144), .ZN(new_n1212));
  INV_X1    g1012(.A(G378), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1136), .A2(new_n1137), .A3(new_n970), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1114), .A2(new_n1120), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1168), .B1(new_n1215), .B2(new_n977), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1213), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1212), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n1207), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1208), .A2(G2897), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT60), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n689), .B1(new_n1173), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n1174), .B2(new_n1221), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(G384), .A3(new_n1199), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G384), .B1(new_n1223), .B2(new_n1199), .ZN(new_n1226));
  OAI21_X1  g1026(.A(KEYINPUT123), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1223), .A2(new_n1199), .ZN(new_n1228));
  INV_X1    g1028(.A(G384), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT123), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(new_n1231), .A3(new_n1224), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1220), .B1(new_n1227), .B2(new_n1232), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1232), .A2(new_n1220), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1211), .B1(new_n1219), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1208), .B1(new_n1212), .B2(new_n1217), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1237), .A2(KEYINPUT62), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT62), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1236), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(G393), .B(G396), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(G387), .A2(G390), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1201), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1242), .B1(new_n1201), .B2(new_n1243), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT126), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1241), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT63), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1246), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT61), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(new_n1253), .A3(new_n1244), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1219), .B2(new_n1235), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT124), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1238), .A2(KEYINPUT63), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1218), .A2(new_n1257), .A3(new_n1207), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1251), .A2(new_n1255), .A3(new_n1256), .A4(new_n1258), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1245), .A2(KEYINPUT61), .A3(new_n1246), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1258), .B(new_n1260), .C1(new_n1261), .C2(new_n1237), .ZN(new_n1262));
  OAI21_X1  g1062(.A(KEYINPUT124), .B1(new_n1262), .B2(new_n1250), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1249), .A2(new_n1259), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT127), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT127), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1249), .A2(new_n1263), .A3(new_n1266), .A4(new_n1259), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(G405));
  AOI21_X1  g1068(.A(G378), .B1(new_n1145), .B2(new_n1171), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1212), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1271), .B(new_n1238), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(new_n1248), .ZN(G402));
endmodule


