//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT67), .Z(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G221), .A4(G218), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT68), .Z(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(G137), .A3(new_n461), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(new_n470), .ZN(G160));
  OAI21_X1  g046(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G112), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n472), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT69), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n477), .A2(new_n461), .ZN(new_n481));
  AOI211_X1 g056(.A(new_n474), .B(new_n480), .C1(G124), .C2(new_n481), .ZN(G162));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(new_n461), .A3(G138), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n477), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(G126), .B(G2105), .C1(new_n475), .C2(new_n476), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR3_X1   g063(.A1(new_n488), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n462), .A2(KEYINPUT4), .A3(new_n489), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n486), .A2(new_n487), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n487), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n497), .A2(KEYINPUT71), .A3(new_n486), .A4(new_n490), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT72), .B1(new_n501), .B2(G651), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n507), .B1(new_n504), .B2(KEYINPUT6), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n501), .A2(KEYINPUT73), .A3(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n506), .A2(new_n510), .A3(G50), .A4(G543), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n506), .A2(new_n510), .A3(G88), .A4(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G62), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n516), .B1(new_n512), .B2(new_n513), .ZN(new_n517));
  AND2_X1   g092(.A1(G75), .A2(G543), .ZN(new_n518));
  OAI21_X1  g093(.A(G651), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n511), .A2(new_n515), .A3(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT74), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n524), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n523), .A2(new_n528), .A3(new_n525), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n506), .A2(new_n510), .A3(G89), .A4(new_n514), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n506), .A2(new_n510), .A3(G51), .A4(G543), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g110(.A(KEYINPUT75), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NOR3_X1   g112(.A1(new_n532), .A2(KEYINPUT75), .A3(new_n535), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(G168));
  NAND2_X1  g115(.A1(new_n506), .A2(new_n510), .ZN(new_n541));
  INV_X1    g116(.A(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G52), .ZN(new_n544));
  INV_X1    g119(.A(new_n514), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G90), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n504), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n544), .A2(new_n547), .A3(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  NAND2_X1  g126(.A1(new_n543), .A2(G43), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n546), .A2(G81), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(new_n504), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  AND2_X1   g137(.A1(new_n506), .A2(new_n510), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT9), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n543), .A2(new_n567), .A3(G53), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n545), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n546), .A2(G91), .B1(new_n572), .B2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(new_n535), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n575), .A2(new_n576), .A3(new_n530), .A4(new_n531), .ZN(new_n577));
  AND3_X1   g152(.A1(new_n577), .A2(new_n536), .A3(KEYINPUT76), .ZN(new_n578));
  AOI21_X1  g153(.A(KEYINPUT76), .B1(new_n577), .B2(new_n536), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G286));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n520), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n511), .A2(new_n515), .A3(new_n519), .A4(KEYINPUT77), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(G303));
  OAI21_X1  g160(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT78), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n543), .A2(G49), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n546), .A2(G87), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G288));
  NAND4_X1  g165(.A1(new_n506), .A2(new_n510), .A3(G48), .A4(G543), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n506), .A2(new_n510), .A3(G86), .A4(new_n514), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n512), .B2(new_n513), .ZN(new_n594));
  AND2_X1   g169(.A1(G73), .A2(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n591), .A2(new_n592), .A3(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n543), .A2(G47), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n563), .A2(new_n514), .ZN(new_n600));
  XOR2_X1   g175(.A(KEYINPUT79), .B(G85), .Z(new_n601));
  OAI221_X1 g176(.A(new_n598), .B1(new_n504), .B2(new_n599), .C1(new_n600), .C2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  XNOR2_X1  g179(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n605));
  OR3_X1    g180(.A1(new_n600), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n600), .B2(new_n604), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n504), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(G54), .B2(new_n543), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n606), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n603), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n603), .B1(new_n612), .B2(G868), .ZN(G321));
  NOR2_X1   g189(.A1(G299), .A2(G868), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n580), .B2(G868), .ZN(G297));
  AOI21_X1  g191(.A(new_n615), .B1(new_n580), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n612), .B1(new_n618), .B2(G860), .ZN(G148));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n556), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n611), .A2(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n620), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n478), .A2(G135), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT84), .Z(new_n626));
  NAND2_X1  g201(.A1(new_n481), .A2(G123), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n461), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT85), .B(G2096), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n462), .A2(new_n468), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT82), .B(KEYINPUT13), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(KEYINPUT83), .A2(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OR3_X1    g214(.A1(new_n639), .A2(KEYINPUT83), .A3(G2100), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(KEYINPUT83), .B2(G2100), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n632), .A2(new_n640), .A3(new_n641), .ZN(G156));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(G14), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n661), .B(KEYINPUT17), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n663), .B1(new_n665), .B2(new_n662), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT87), .Z(new_n667));
  NAND3_X1  g242(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT86), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT18), .ZN(new_n670));
  OR3_X1    g245(.A1(new_n665), .A2(new_n660), .A3(new_n662), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT88), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n682));
  OR2_X1    g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n678), .A2(new_n680), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n676), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n684), .A2(new_n681), .A3(new_n676), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n682), .B1(new_n681), .B2(new_n676), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT90), .B(KEYINPUT91), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n693), .B(new_n696), .ZN(G229));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n698), .A2(G24), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G290), .B2(G16), .ZN(new_n700));
  INV_X1    g275(.A(G1986), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G25), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n478), .A2(G131), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n481), .A2(G119), .ZN(new_n706));
  INV_X1    g281(.A(G95), .ZN(new_n707));
  AND3_X1   g282(.A1(new_n707), .A2(new_n461), .A3(KEYINPUT92), .ZN(new_n708));
  AOI21_X1  g283(.A(KEYINPUT92), .B1(new_n707), .B2(new_n461), .ZN(new_n709));
  OAI221_X1 g284(.A(G2104), .B1(G107), .B2(new_n461), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n705), .A2(new_n706), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n704), .B1(new_n712), .B2(new_n703), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT35), .B(G1991), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT93), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n713), .B(new_n715), .Z(new_n716));
  INV_X1    g291(.A(new_n700), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n716), .B1(G1986), .B2(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G6), .B(G305), .S(G16), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT32), .ZN(new_n720));
  INV_X1    g295(.A(G1981), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n698), .A2(G22), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT94), .Z(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G166), .B2(new_n698), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1971), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(KEYINPUT95), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(KEYINPUT95), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n698), .A2(G23), .ZN(new_n729));
  INV_X1    g304(.A(G288), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(new_n698), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT33), .B(G1976), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n722), .A2(new_n727), .A3(new_n728), .A4(new_n733), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n702), .B(new_n718), .C1(new_n734), .C2(KEYINPUT34), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(KEYINPUT34), .B2(new_n734), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n698), .A2(G4), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n612), .B2(new_n698), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1348), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n698), .A2(G19), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n557), .B2(new_n698), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1341), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n703), .A2(G26), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT28), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n478), .A2(G140), .ZN(new_n747));
  INV_X1    g322(.A(G128), .ZN(new_n748));
  INV_X1    g323(.A(new_n481), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(KEYINPUT96), .B1(G104), .B2(G2105), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NOR3_X1   g327(.A1(KEYINPUT96), .A2(G104), .A3(G2105), .ZN(new_n753));
  OAI221_X1 g328(.A(G2104), .B1(G116), .B2(new_n461), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n750), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n746), .B1(new_n757), .B2(new_n703), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2067), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n741), .A2(new_n744), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT97), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n698), .A2(G21), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G168), .B2(new_n698), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G1966), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT101), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n763), .A2(G1966), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n698), .A2(G20), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT23), .Z(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G299), .B2(G16), .ZN(new_n769));
  INV_X1    g344(.A(G1956), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G127), .ZN(new_n772));
  INV_X1    g347(.A(G115), .ZN(new_n773));
  OAI22_X1  g348(.A1(new_n477), .A2(new_n772), .B1(new_n773), .B2(new_n467), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT98), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n461), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n775), .B2(new_n774), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT25), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G139), .B2(new_n478), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT99), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  MUX2_X1   g358(.A(G33), .B(new_n783), .S(G29), .Z(new_n784));
  AOI211_X1 g359(.A(new_n766), .B(new_n771), .C1(G2072), .C2(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n761), .A2(new_n765), .A3(new_n785), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n478), .A2(G141), .B1(G105), .B2(new_n468), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT26), .Z(new_n790));
  INV_X1    g365(.A(G129), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n749), .B2(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(new_n703), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n703), .B2(G32), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT27), .B(G1996), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT24), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n703), .B1(new_n798), .B2(G34), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n798), .B2(G34), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G160), .B2(G29), .ZN(new_n801));
  OAI22_X1  g376(.A1(new_n796), .A2(new_n797), .B1(new_n801), .B2(G2084), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n698), .A2(G5), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G171), .B2(new_n698), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n804), .A2(G1961), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT103), .ZN(new_n807));
  NOR2_X1   g382(.A1(G29), .A2(G35), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G162), .B2(G29), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT29), .ZN(new_n810));
  INV_X1    g385(.A(G2090), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(G164), .A2(G29), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G27), .B2(G29), .ZN(new_n814));
  INV_X1    g389(.A(G2078), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n801), .A2(G2084), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT31), .B(G11), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT30), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n819), .A2(KEYINPUT102), .A3(G28), .ZN(new_n820));
  AOI21_X1  g395(.A(KEYINPUT102), .B1(new_n819), .B2(G28), .ZN(new_n821));
  OAI221_X1 g396(.A(new_n703), .B1(new_n819), .B2(G28), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n818), .B(new_n822), .C1(new_n630), .C2(new_n703), .ZN(new_n823));
  AOI211_X1 g398(.A(new_n817), .B(new_n823), .C1(new_n796), .C2(new_n797), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n814), .A2(new_n815), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n804), .A2(G1961), .ZN(new_n826));
  AND4_X1   g401(.A1(new_n816), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n807), .A2(new_n812), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n784), .A2(G2072), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT100), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n786), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n738), .A2(new_n831), .ZN(G311));
  INV_X1    g407(.A(KEYINPUT104), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n738), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n833), .B1(new_n738), .B2(new_n831), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(G150));
  INV_X1    g411(.A(KEYINPUT105), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(new_n504), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n563), .A2(G55), .A3(G543), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n563), .A2(G93), .A3(new_n514), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n557), .A2(new_n837), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(KEYINPUT105), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n837), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(new_n556), .A3(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n612), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n852), .A2(new_n853), .A3(G860), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n842), .A2(G860), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT37), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n854), .A2(new_n856), .ZN(G145));
  XNOR2_X1  g432(.A(new_n783), .B(new_n794), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n493), .A2(KEYINPUT106), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT106), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n497), .A2(new_n860), .A3(new_n486), .A4(new_n490), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n858), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n481), .A2(G130), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n461), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(G142), .B2(new_n478), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n712), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n635), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n757), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n863), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n630), .B(G160), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G162), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G37), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n872), .A2(new_n874), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XOR2_X1   g454(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(G395));
  NAND2_X1  g456(.A1(new_n842), .A2(new_n620), .ZN(new_n882));
  XOR2_X1   g457(.A(G290), .B(G305), .Z(new_n883));
  XNOR2_X1  g458(.A(G288), .B(G166), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n883), .B(new_n884), .Z(new_n885));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n885), .B1(KEYINPUT108), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(KEYINPUT108), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(G299), .B(new_n611), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(KEYINPUT41), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n844), .A2(new_n847), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n622), .ZN(new_n894));
  MUX2_X1   g469(.A(new_n891), .B(new_n892), .S(new_n894), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n889), .B(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n882), .B1(new_n896), .B2(new_n620), .ZN(G295));
  OAI21_X1  g472(.A(new_n882), .B1(new_n896), .B2(new_n620), .ZN(G331));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n899));
  NOR3_X1   g474(.A1(G171), .A2(new_n537), .A3(new_n538), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT76), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n537), .B2(new_n538), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n577), .A2(new_n536), .A3(KEYINPUT76), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(G171), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n848), .A2(new_n901), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n578), .A2(new_n579), .A3(G301), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n893), .B1(new_n908), .B2(new_n900), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n848), .A2(new_n901), .A3(new_n905), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(KEYINPUT109), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n892), .A2(new_n907), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n885), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(new_n891), .A3(new_n910), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n876), .ZN(new_n916));
  INV_X1    g491(.A(new_n910), .ZN(new_n917));
  INV_X1    g492(.A(new_n909), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n892), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n890), .B1(new_n911), .B2(new_n907), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT110), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI211_X1 g497(.A(KEYINPUT110), .B(new_n890), .C1(new_n911), .C2(new_n907), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n885), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT111), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT111), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n926), .B(new_n885), .C1(new_n922), .C2(new_n923), .ZN(new_n927));
  AOI211_X1 g502(.A(new_n899), .B(new_n916), .C1(new_n925), .C2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n916), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n912), .A2(new_n914), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n885), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT43), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT44), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n934));
  AOI211_X1 g509(.A(KEYINPUT43), .B(new_n916), .C1(new_n925), .C2(new_n927), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n899), .B1(new_n929), .B2(new_n931), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n937), .ZN(G397));
  INV_X1    g513(.A(KEYINPUT125), .ZN(new_n939));
  NAND3_X1  g514(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n583), .A2(G8), .A3(new_n584), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT55), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G125), .ZN(new_n946));
  OR2_X1    g521(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n947));
  NAND2_X1  g522(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n464), .ZN(new_n950));
  OAI21_X1  g525(.A(G2105), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n951), .A2(G40), .A3(new_n469), .A4(new_n466), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n477), .A2(new_n483), .A3(new_n485), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT4), .B1(new_n462), .B2(new_n489), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(G1384), .B1(new_n956), .B2(new_n497), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n953), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(G1384), .B1(new_n495), .B2(new_n498), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n962), .A2(G1384), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n859), .A2(new_n861), .A3(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n953), .B(new_n964), .C1(new_n960), .C2(KEYINPUT45), .ZN(new_n965));
  INV_X1    g540(.A(G1971), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n961), .A2(new_n811), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G8), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n945), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT113), .ZN(new_n971));
  NAND2_X1  g546(.A1(G305), .A2(G1981), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n591), .A2(new_n592), .A3(new_n596), .A4(new_n721), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n971), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  AOI211_X1 g552(.A(KEYINPUT113), .B(new_n975), .C1(new_n972), .C2(new_n973), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n493), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n981), .A2(new_n952), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(new_n968), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n972), .A2(KEYINPUT49), .A3(new_n973), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n970), .B1(new_n979), .B2(new_n985), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n983), .A2(new_n984), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n987), .B(KEYINPUT114), .C1(new_n977), .C2(new_n978), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n965), .A2(new_n966), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n952), .B1(new_n957), .B2(new_n958), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(new_n960), .B2(new_n958), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(G2090), .ZN(new_n993));
  OAI211_X1 g568(.A(G8), .B(new_n944), .C1(new_n990), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n957), .A2(new_n953), .ZN(new_n995));
  INV_X1    g570(.A(G1976), .ZN(new_n996));
  OAI211_X1 g571(.A(G8), .B(new_n995), .C1(G288), .C2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT52), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n730), .B2(G1976), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n998), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n969), .A2(new_n989), .A3(new_n994), .A4(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n965), .B2(G2078), .ZN(new_n1005));
  INV_X1    g580(.A(G1961), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n992), .A2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(KEYINPUT116), .B(new_n953), .C1(new_n957), .C2(KEYINPUT45), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT45), .B1(new_n493), .B2(new_n980), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1009), .B1(new_n1010), .B2(new_n952), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT71), .B1(new_n956), .B2(new_n497), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n486), .A2(new_n490), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1013), .A2(new_n494), .A3(new_n496), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n963), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1008), .A2(new_n1011), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n815), .A2(KEYINPUT53), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1005), .B(new_n1007), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(G171), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1003), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n952), .B1(new_n981), .B2(new_n962), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1021), .A2(KEYINPUT116), .B1(new_n499), .B2(new_n963), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1966), .B1(new_n1022), .B2(new_n1011), .ZN(new_n1023));
  INV_X1    g598(.A(G2084), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n991), .B(new_n1024), .C1(new_n960), .C2(new_n958), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(G168), .A2(new_n968), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1966), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1016), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n968), .B1(new_n1032), .B2(new_n1025), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1033), .A2(KEYINPUT51), .A3(new_n1028), .ZN(new_n1034));
  OAI211_X1 g609(.A(KEYINPUT121), .B(G8), .C1(new_n1023), .C2(new_n1026), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n1029), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1033), .A2(KEYINPUT121), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT51), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1034), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1028), .B1(new_n1033), .B2(KEYINPUT121), .ZN(new_n1042));
  OAI21_X1  g617(.A(G8), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT121), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT122), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1030), .B1(new_n1040), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT62), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1020), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1030), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1034), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1046), .B2(KEYINPUT122), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(KEYINPUT62), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n939), .B1(new_n1050), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n965), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT56), .B(G2072), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n959), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n960), .A2(new_n958), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1956), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n1066));
  NAND2_X1  g641(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n569), .A2(new_n1068), .A3(new_n573), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1065), .A2(new_n1066), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1059), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n965), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1070), .B1(new_n1073), .B2(new_n1063), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT120), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1348), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n992), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  INV_X1    g654(.A(G2067), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n982), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1079), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1083), .A2(new_n611), .A3(new_n1084), .ZN(new_n1085));
  OAI22_X1  g660(.A1(new_n1076), .A2(new_n1085), .B1(new_n1070), .B2(new_n1065), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT61), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1073), .A2(new_n1063), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1071), .A2(new_n1090), .A3(new_n1075), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT60), .B(new_n611), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1074), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1073), .A2(new_n1070), .A3(new_n1063), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1087), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  XOR2_X1   g670(.A(KEYINPUT58), .B(G1341), .Z(new_n1096));
  NAND2_X1  g671(.A1(new_n995), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n965), .B2(G1996), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n557), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT59), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(new_n1101), .A3(new_n557), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1091), .A2(new_n1092), .A3(new_n1095), .A4(new_n1103), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1083), .A2(KEYINPUT60), .A3(new_n1084), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT119), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1108), .B2(new_n1082), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1105), .A2(new_n1109), .A3(new_n611), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1086), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT54), .B1(new_n1018), .B2(G171), .ZN(new_n1112));
  INV_X1    g687(.A(new_n862), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n962), .B1(new_n1113), .B2(G1384), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT123), .B(G2078), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1115), .A2(KEYINPUT53), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1114), .A2(new_n953), .A3(new_n964), .A4(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1117), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1118), .A2(KEYINPUT124), .ZN(new_n1119));
  AOI21_X1  g694(.A(G301), .B1(new_n1118), .B2(KEYINPUT124), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1112), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1117), .A2(G301), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT54), .B1(new_n1019), .B2(new_n1122), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1121), .A2(new_n1003), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1055), .A2(new_n1111), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n994), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1001), .B1(new_n986), .B2(new_n988), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT115), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI211_X1 g704(.A(KEYINPUT115), .B(new_n1001), .C1(new_n986), .C2(new_n988), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1126), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI211_X1 g706(.A(G1976), .B(G288), .C1(new_n986), .C2(new_n988), .ZN(new_n1132));
  INV_X1    g707(.A(new_n973), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n983), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(G8), .B(new_n580), .C1(new_n1023), .C2(new_n1026), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT117), .B1(new_n1033), .B2(new_n580), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT118), .B1(new_n1140), .B2(new_n1003), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n969), .A2(new_n994), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1033), .A2(KEYINPUT117), .A3(new_n580), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT118), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1143), .A2(new_n1146), .A3(new_n1147), .A4(new_n1127), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1141), .A2(new_n1142), .A3(new_n1148), .ZN(new_n1149));
  OAI22_X1  g724(.A1(new_n1058), .A2(G1971), .B1(G2090), .B2(new_n992), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n944), .B1(new_n1150), .B2(G8), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1126), .A2(new_n1151), .A3(new_n1142), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1152), .B(new_n1146), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1135), .B1(new_n1149), .B2(new_n1153), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1125), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1055), .A2(KEYINPUT62), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(KEYINPUT125), .A4(new_n1020), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1057), .A2(new_n1155), .A3(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n756), .B(new_n1080), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n793), .B(G1996), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n712), .A2(new_n715), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n712), .A2(new_n715), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(G290), .B(new_n701), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1114), .A2(new_n952), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1159), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1163), .ZN(new_n1172));
  OAI22_X1  g747(.A1(new_n1172), .A2(new_n1164), .B1(G2067), .B2(new_n756), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n1169), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1174), .B(KEYINPUT126), .Z(new_n1175));
  INV_X1    g750(.A(new_n1169), .ZN(new_n1176));
  OR3_X1    g751(.A1(new_n1176), .A2(G1986), .A3(G290), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT48), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  OAI22_X1  g754(.A1(new_n1177), .A2(new_n1178), .B1(new_n1166), .B2(new_n1176), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1175), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT46), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n794), .B1(new_n1182), .B2(G1996), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1169), .B1(new_n1161), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1182), .B1(new_n1176), .B2(G1996), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1185), .A2(KEYINPUT127), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1185), .A2(KEYINPUT127), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1184), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g763(.A(new_n1188), .B(KEYINPUT47), .Z(new_n1189));
  NOR2_X1   g764(.A1(new_n1181), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1171), .A2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g766(.A1(new_n935), .A2(new_n936), .ZN(new_n1193));
  OAI21_X1  g767(.A(G319), .B1(new_n656), .B2(new_n657), .ZN(new_n1194));
  NOR3_X1   g768(.A1(G229), .A2(G227), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g769(.A(new_n1195), .B1(new_n877), .B2(new_n878), .ZN(new_n1196));
  NOR2_X1   g770(.A1(new_n1193), .A2(new_n1196), .ZN(G308));
  OAI221_X1 g771(.A(new_n1195), .B1(new_n878), .B2(new_n877), .C1(new_n935), .C2(new_n936), .ZN(G225));
endmodule


