

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U555 ( .A(n551), .Z(n521) );
  NAND2_X2 U556 ( .A1(n729), .A2(G8), .ZN(n768) );
  AND2_X2 U557 ( .A1(n528), .A2(G2104), .ZN(n882) );
  NOR2_X1 U558 ( .A1(G651), .A2(G543), .ZN(n643) );
  AND2_X1 U559 ( .A1(n553), .A2(n552), .ZN(n522) );
  INV_X1 U560 ( .A(KEYINPUT29), .ZN(n709) );
  XNOR2_X1 U561 ( .A(n710), .B(n709), .ZN(n716) );
  INV_X1 U562 ( .A(KEYINPUT99), .ZN(n727) );
  XOR2_X1 U563 ( .A(KEYINPUT65), .B(n539), .Z(n646) );
  AND2_X1 U564 ( .A1(n533), .A2(n532), .ZN(G160) );
  XNOR2_X1 U565 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n524) );
  NOR2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XNOR2_X1 U567 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U568 ( .A(KEYINPUT66), .B(n525), .ZN(n603) );
  NAND2_X1 U569 ( .A1(n603), .A2(G137), .ZN(n533) );
  INV_X1 U570 ( .A(G2105), .ZN(n528) );
  NOR2_X1 U571 ( .A1(G2104), .A2(n528), .ZN(n551) );
  NAND2_X1 U572 ( .A1(G125), .A2(n521), .ZN(n527) );
  AND2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n879) );
  NAND2_X1 U574 ( .A1(G113), .A2(n879), .ZN(n526) );
  AND2_X1 U575 ( .A1(n527), .A2(n526), .ZN(n531) );
  NAND2_X1 U576 ( .A1(G101), .A2(n882), .ZN(n529) );
  XOR2_X1 U577 ( .A(KEYINPUT23), .B(n529), .Z(n530) );
  AND2_X1 U578 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U579 ( .A1(G90), .A2(n643), .ZN(n535) );
  XOR2_X1 U580 ( .A(G543), .B(KEYINPUT0), .Z(n639) );
  INV_X1 U581 ( .A(G651), .ZN(n537) );
  NOR2_X1 U582 ( .A1(n639), .A2(n537), .ZN(n645) );
  NAND2_X1 U583 ( .A1(G77), .A2(n645), .ZN(n534) );
  NAND2_X1 U584 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U585 ( .A(KEYINPUT9), .B(n536), .ZN(n544) );
  NOR2_X1 U586 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n538), .Z(n649) );
  NAND2_X1 U588 ( .A1(G64), .A2(n649), .ZN(n541) );
  NOR2_X1 U589 ( .A1(G651), .A2(n639), .ZN(n539) );
  NAND2_X1 U590 ( .A1(G52), .A2(n646), .ZN(n540) );
  NAND2_X1 U591 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U592 ( .A(KEYINPUT70), .B(n542), .Z(n543) );
  NAND2_X1 U593 ( .A1(n544), .A2(n543), .ZN(G301) );
  INV_X1 U594 ( .A(G301), .ZN(G171) );
  AND2_X1 U595 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U596 ( .A1(G65), .A2(n649), .ZN(n546) );
  NAND2_X1 U597 ( .A1(G53), .A2(n646), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U599 ( .A1(G91), .A2(n643), .ZN(n548) );
  NAND2_X1 U600 ( .A1(G78), .A2(n645), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U602 ( .A1(n550), .A2(n549), .ZN(n971) );
  INV_X1 U603 ( .A(n971), .ZN(G299) );
  AND2_X1 U604 ( .A1(n603), .A2(G138), .ZN(n556) );
  NAND2_X1 U605 ( .A1(G126), .A2(n521), .ZN(n553) );
  NAND2_X1 U606 ( .A1(G114), .A2(n879), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n882), .A2(G102), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n522), .A2(n554), .ZN(n555) );
  NOR2_X1 U609 ( .A1(n556), .A2(n555), .ZN(G164) );
  INV_X1 U610 ( .A(G57), .ZN(G237) );
  NAND2_X1 U611 ( .A1(G7), .A2(G661), .ZN(n557) );
  XNOR2_X1 U612 ( .A(n557), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U613 ( .A(G223), .ZN(n827) );
  NAND2_X1 U614 ( .A1(n827), .A2(G567), .ZN(n558) );
  XNOR2_X1 U615 ( .A(n558), .B(KEYINPUT71), .ZN(n559) );
  XNOR2_X1 U616 ( .A(KEYINPUT11), .B(n559), .ZN(G234) );
  NAND2_X1 U617 ( .A1(n643), .A2(G81), .ZN(n560) );
  XNOR2_X1 U618 ( .A(n560), .B(KEYINPUT12), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G68), .A2(n645), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U621 ( .A(n563), .B(KEYINPUT13), .ZN(n565) );
  NAND2_X1 U622 ( .A1(G43), .A2(n646), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n568) );
  NAND2_X1 U624 ( .A1(n649), .A2(G56), .ZN(n566) );
  XOR2_X1 U625 ( .A(KEYINPUT14), .B(n566), .Z(n567) );
  NOR2_X1 U626 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X2 U627 ( .A(KEYINPUT72), .B(n569), .ZN(n969) );
  NAND2_X1 U628 ( .A1(G860), .A2(n969), .ZN(G153) );
  NAND2_X1 U629 ( .A1(G868), .A2(G301), .ZN(n579) );
  NAND2_X1 U630 ( .A1(G54), .A2(n646), .ZN(n576) );
  NAND2_X1 U631 ( .A1(G92), .A2(n643), .ZN(n571) );
  NAND2_X1 U632 ( .A1(G66), .A2(n649), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n571), .A2(n570), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G79), .A2(n645), .ZN(n572) );
  XNOR2_X1 U635 ( .A(KEYINPUT73), .B(n572), .ZN(n573) );
  NOR2_X1 U636 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U638 ( .A(n577), .B(KEYINPUT15), .ZN(n970) );
  OR2_X1 U639 ( .A1(n970), .A2(G868), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n579), .A2(n578), .ZN(G284) );
  NAND2_X1 U641 ( .A1(n643), .A2(G89), .ZN(n580) );
  XNOR2_X1 U642 ( .A(n580), .B(KEYINPUT4), .ZN(n582) );
  NAND2_X1 U643 ( .A1(G76), .A2(n645), .ZN(n581) );
  NAND2_X1 U644 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U645 ( .A(n583), .B(KEYINPUT5), .ZN(n588) );
  NAND2_X1 U646 ( .A1(G63), .A2(n649), .ZN(n585) );
  NAND2_X1 U647 ( .A1(G51), .A2(n646), .ZN(n584) );
  NAND2_X1 U648 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U649 ( .A(KEYINPUT6), .B(n586), .Z(n587) );
  NAND2_X1 U650 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U651 ( .A(n589), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U652 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U653 ( .A1(G868), .A2(G299), .ZN(n590) );
  XNOR2_X1 U654 ( .A(n590), .B(KEYINPUT74), .ZN(n592) );
  INV_X1 U655 ( .A(G868), .ZN(n655) );
  NOR2_X1 U656 ( .A1(n655), .A2(G286), .ZN(n591) );
  NOR2_X1 U657 ( .A1(n592), .A2(n591), .ZN(G297) );
  INV_X1 U658 ( .A(G860), .ZN(n593) );
  NAND2_X1 U659 ( .A1(n593), .A2(G559), .ZN(n594) );
  NAND2_X1 U660 ( .A1(n594), .A2(n970), .ZN(n595) );
  XNOR2_X1 U661 ( .A(n595), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U662 ( .A1(n970), .A2(G868), .ZN(n596) );
  NOR2_X1 U663 ( .A1(G559), .A2(n596), .ZN(n598) );
  AND2_X1 U664 ( .A1(n969), .A2(n655), .ZN(n597) );
  NOR2_X1 U665 ( .A1(n598), .A2(n597), .ZN(G282) );
  NAND2_X1 U666 ( .A1(G99), .A2(n882), .ZN(n600) );
  NAND2_X1 U667 ( .A1(G111), .A2(n879), .ZN(n599) );
  NAND2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U669 ( .A(KEYINPUT76), .B(n601), .ZN(n608) );
  NAND2_X1 U670 ( .A1(n521), .A2(G123), .ZN(n602) );
  XNOR2_X1 U671 ( .A(n602), .B(KEYINPUT18), .ZN(n605) );
  BUF_X1 U672 ( .A(n603), .Z(n883) );
  NAND2_X1 U673 ( .A1(G135), .A2(n883), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U675 ( .A(KEYINPUT75), .B(n606), .Z(n607) );
  NOR2_X1 U676 ( .A1(n608), .A2(n607), .ZN(n922) );
  XNOR2_X1 U677 ( .A(n922), .B(G2096), .ZN(n610) );
  INV_X1 U678 ( .A(G2100), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n610), .A2(n609), .ZN(G156) );
  NAND2_X1 U680 ( .A1(G67), .A2(n649), .ZN(n612) );
  NAND2_X1 U681 ( .A1(G55), .A2(n646), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U683 ( .A1(n645), .A2(G80), .ZN(n613) );
  XOR2_X1 U684 ( .A(KEYINPUT78), .B(n613), .Z(n614) );
  NOR2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U686 ( .A1(n643), .A2(G93), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n617), .A2(n616), .ZN(n659) );
  XNOR2_X1 U688 ( .A(KEYINPUT77), .B(n969), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n970), .A2(G559), .ZN(n664) );
  XNOR2_X1 U690 ( .A(n618), .B(n664), .ZN(n619) );
  NOR2_X1 U691 ( .A1(G860), .A2(n619), .ZN(n620) );
  XOR2_X1 U692 ( .A(n659), .B(n620), .Z(G145) );
  NAND2_X1 U693 ( .A1(G88), .A2(n643), .ZN(n622) );
  NAND2_X1 U694 ( .A1(G75), .A2(n645), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n627) );
  NAND2_X1 U696 ( .A1(G62), .A2(n649), .ZN(n623) );
  XOR2_X1 U697 ( .A(KEYINPUT81), .B(n623), .Z(n625) );
  NAND2_X1 U698 ( .A1(n646), .A2(G50), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n627), .A2(n626), .ZN(G166) );
  XOR2_X1 U701 ( .A(KEYINPUT80), .B(KEYINPUT2), .Z(n629) );
  NAND2_X1 U702 ( .A1(G73), .A2(n645), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n629), .B(n628), .ZN(n633) );
  NAND2_X1 U704 ( .A1(G86), .A2(n643), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G48), .A2(n646), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n649), .A2(G61), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U710 ( .A1(G49), .A2(n646), .ZN(n637) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U713 ( .A1(n649), .A2(n638), .ZN(n642) );
  NAND2_X1 U714 ( .A1(G87), .A2(n639), .ZN(n640) );
  XOR2_X1 U715 ( .A(KEYINPUT79), .B(n640), .Z(n641) );
  NAND2_X1 U716 ( .A1(n642), .A2(n641), .ZN(G288) );
  NAND2_X1 U717 ( .A1(n643), .A2(G85), .ZN(n644) );
  XNOR2_X1 U718 ( .A(KEYINPUT68), .B(n644), .ZN(n654) );
  NAND2_X1 U719 ( .A1(G72), .A2(n645), .ZN(n648) );
  NAND2_X1 U720 ( .A1(G47), .A2(n646), .ZN(n647) );
  NAND2_X1 U721 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U722 ( .A1(G60), .A2(n649), .ZN(n650) );
  XNOR2_X1 U723 ( .A(KEYINPUT69), .B(n650), .ZN(n651) );
  NOR2_X1 U724 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U725 ( .A1(n654), .A2(n653), .ZN(G290) );
  NAND2_X1 U726 ( .A1(n655), .A2(n659), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n656), .B(KEYINPUT82), .ZN(n667) );
  XNOR2_X1 U728 ( .A(G166), .B(G305), .ZN(n657) );
  XNOR2_X1 U729 ( .A(n657), .B(n969), .ZN(n658) );
  XOR2_X1 U730 ( .A(n659), .B(n658), .Z(n661) );
  XNOR2_X1 U731 ( .A(G288), .B(KEYINPUT19), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U733 ( .A(n662), .B(G290), .ZN(n663) );
  XNOR2_X1 U734 ( .A(n663), .B(G299), .ZN(n895) );
  XNOR2_X1 U735 ( .A(n895), .B(n664), .ZN(n665) );
  NAND2_X1 U736 ( .A1(G868), .A2(n665), .ZN(n666) );
  NAND2_X1 U737 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U738 ( .A1(G2084), .A2(G2078), .ZN(n668) );
  XOR2_X1 U739 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n671), .A2(G2072), .ZN(n672) );
  XOR2_X1 U743 ( .A(KEYINPUT83), .B(n672), .Z(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U745 ( .A1(G132), .A2(G82), .ZN(n673) );
  XNOR2_X1 U746 ( .A(n673), .B(KEYINPUT22), .ZN(n674) );
  XNOR2_X1 U747 ( .A(n674), .B(KEYINPUT84), .ZN(n675) );
  NOR2_X1 U748 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U749 ( .A1(G96), .A2(n676), .ZN(n831) );
  NAND2_X1 U750 ( .A1(n831), .A2(G2106), .ZN(n680) );
  NAND2_X1 U751 ( .A1(G69), .A2(G120), .ZN(n677) );
  NOR2_X1 U752 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U753 ( .A1(G108), .A2(n678), .ZN(n832) );
  NAND2_X1 U754 ( .A1(n832), .A2(G567), .ZN(n679) );
  NAND2_X1 U755 ( .A1(n680), .A2(n679), .ZN(n833) );
  NAND2_X1 U756 ( .A1(G661), .A2(G483), .ZN(n681) );
  NOR2_X1 U757 ( .A1(n833), .A2(n681), .ZN(n830) );
  NAND2_X1 U758 ( .A1(n830), .A2(G36), .ZN(G176) );
  XNOR2_X1 U759 ( .A(KEYINPUT85), .B(G166), .ZN(G303) );
  NAND2_X1 U760 ( .A1(G160), .A2(G40), .ZN(n790) );
  INV_X1 U761 ( .A(n790), .ZN(n683) );
  NOR2_X1 U762 ( .A1(G164), .A2(G1384), .ZN(n791) );
  NAND2_X1 U763 ( .A1(n683), .A2(n791), .ZN(n684) );
  XNOR2_X2 U764 ( .A(n684), .B(KEYINPUT64), .ZN(n729) );
  INV_X1 U765 ( .A(n729), .ZN(n712) );
  NAND2_X1 U766 ( .A1(n712), .A2(G1996), .ZN(n685) );
  XNOR2_X1 U767 ( .A(n685), .B(KEYINPUT26), .ZN(n686) );
  NAND2_X1 U768 ( .A1(n686), .A2(n969), .ZN(n689) );
  NAND2_X1 U769 ( .A1(n729), .A2(G1341), .ZN(n687) );
  XOR2_X1 U770 ( .A(KEYINPUT96), .B(n687), .Z(n688) );
  NOR2_X2 U771 ( .A1(n689), .A2(n688), .ZN(n696) );
  NAND2_X1 U772 ( .A1(n696), .A2(n970), .ZN(n694) );
  NAND2_X1 U773 ( .A1(n729), .A2(G1348), .ZN(n692) );
  INV_X1 U774 ( .A(KEYINPUT94), .ZN(n690) );
  XNOR2_X1 U775 ( .A(n690), .B(n729), .ZN(n711) );
  NAND2_X1 U776 ( .A1(G2067), .A2(n711), .ZN(n691) );
  NAND2_X1 U777 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U778 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U779 ( .A(KEYINPUT97), .B(n695), .Z(n698) );
  OR2_X1 U780 ( .A1(n970), .A2(n696), .ZN(n697) );
  NAND2_X1 U781 ( .A1(n698), .A2(n697), .ZN(n703) );
  NAND2_X1 U782 ( .A1(n711), .A2(G2072), .ZN(n699) );
  XNOR2_X1 U783 ( .A(n699), .B(KEYINPUT27), .ZN(n701) );
  INV_X1 U784 ( .A(G1956), .ZN(n998) );
  NOR2_X1 U785 ( .A1(n998), .A2(n711), .ZN(n700) );
  NOR2_X1 U786 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U787 ( .A1(n971), .A2(n704), .ZN(n702) );
  NAND2_X1 U788 ( .A1(n703), .A2(n702), .ZN(n708) );
  NOR2_X1 U789 ( .A1(n971), .A2(n704), .ZN(n706) );
  XNOR2_X1 U790 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n705) );
  XNOR2_X1 U791 ( .A(n706), .B(n705), .ZN(n707) );
  NAND2_X1 U792 ( .A1(n708), .A2(n707), .ZN(n710) );
  XNOR2_X1 U793 ( .A(G2078), .B(KEYINPUT25), .ZN(n945) );
  NAND2_X1 U794 ( .A1(n711), .A2(n945), .ZN(n714) );
  OR2_X1 U795 ( .A1(n712), .A2(G1961), .ZN(n713) );
  NAND2_X1 U796 ( .A1(n714), .A2(n713), .ZN(n717) );
  NAND2_X1 U797 ( .A1(n717), .A2(G171), .ZN(n715) );
  NAND2_X1 U798 ( .A1(n716), .A2(n715), .ZN(n726) );
  NOR2_X1 U799 ( .A1(G171), .A2(n717), .ZN(n722) );
  NOR2_X1 U800 ( .A1(G1966), .A2(n768), .ZN(n740) );
  NOR2_X1 U801 ( .A1(n729), .A2(G2084), .ZN(n737) );
  NOR2_X1 U802 ( .A1(n740), .A2(n737), .ZN(n718) );
  NAND2_X1 U803 ( .A1(G8), .A2(n718), .ZN(n719) );
  XNOR2_X1 U804 ( .A(KEYINPUT30), .B(n719), .ZN(n720) );
  NOR2_X1 U805 ( .A1(G168), .A2(n720), .ZN(n721) );
  NOR2_X1 U806 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U807 ( .A(n723), .B(KEYINPUT31), .Z(n724) );
  XNOR2_X1 U808 ( .A(KEYINPUT98), .B(n724), .ZN(n725) );
  NAND2_X1 U809 ( .A1(n726), .A2(n725), .ZN(n738) );
  NAND2_X1 U810 ( .A1(G286), .A2(n738), .ZN(n728) );
  XNOR2_X1 U811 ( .A(n728), .B(n727), .ZN(n734) );
  NOR2_X1 U812 ( .A1(n729), .A2(G2090), .ZN(n731) );
  NOR2_X1 U813 ( .A1(G1971), .A2(n768), .ZN(n730) );
  NOR2_X1 U814 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U815 ( .A1(G303), .A2(n732), .ZN(n733) );
  NAND2_X1 U816 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U817 ( .A1(n735), .A2(G8), .ZN(n736) );
  XNOR2_X1 U818 ( .A(n736), .B(KEYINPUT32), .ZN(n744) );
  NAND2_X1 U819 ( .A1(G8), .A2(n737), .ZN(n742) );
  INV_X1 U820 ( .A(n738), .ZN(n739) );
  NOR2_X1 U821 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U822 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U823 ( .A1(n744), .A2(n743), .ZN(n753) );
  NOR2_X1 U824 ( .A1(G2090), .A2(G303), .ZN(n745) );
  NAND2_X1 U825 ( .A1(G8), .A2(n745), .ZN(n746) );
  NAND2_X1 U826 ( .A1(n753), .A2(n746), .ZN(n747) );
  XOR2_X1 U827 ( .A(KEYINPUT103), .B(n747), .Z(n748) );
  NAND2_X1 U828 ( .A1(n748), .A2(n768), .ZN(n749) );
  XNOR2_X1 U829 ( .A(n749), .B(KEYINPUT104), .ZN(n772) );
  NAND2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n977) );
  NOR2_X1 U831 ( .A1(G288), .A2(G1976), .ZN(n750) );
  XNOR2_X1 U832 ( .A(n750), .B(KEYINPUT100), .ZN(n976) );
  NOR2_X1 U833 ( .A1(G1971), .A2(G303), .ZN(n751) );
  XOR2_X1 U834 ( .A(n751), .B(KEYINPUT101), .Z(n752) );
  NOR2_X1 U835 ( .A1(n976), .A2(n752), .ZN(n754) );
  NAND2_X1 U836 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U837 ( .A1(n977), .A2(n755), .ZN(n756) );
  NOR2_X1 U838 ( .A1(n756), .A2(n768), .ZN(n757) );
  NOR2_X1 U839 ( .A1(n757), .A2(KEYINPUT33), .ZN(n763) );
  INV_X1 U840 ( .A(n976), .ZN(n758) );
  NOR2_X1 U841 ( .A1(n768), .A2(n758), .ZN(n759) );
  AND2_X1 U842 ( .A1(KEYINPUT33), .A2(n759), .ZN(n761) );
  XNOR2_X1 U843 ( .A(KEYINPUT102), .B(G1981), .ZN(n760) );
  XNOR2_X1 U844 ( .A(n760), .B(G305), .ZN(n966) );
  OR2_X1 U845 ( .A1(n761), .A2(n966), .ZN(n762) );
  NOR2_X1 U846 ( .A1(n763), .A2(n762), .ZN(n770) );
  XNOR2_X1 U847 ( .A(KEYINPUT24), .B(KEYINPUT93), .ZN(n764) );
  XNOR2_X1 U848 ( .A(n764), .B(KEYINPUT92), .ZN(n766) );
  NOR2_X1 U849 ( .A1(G1981), .A2(G305), .ZN(n765) );
  XNOR2_X1 U850 ( .A(n766), .B(n765), .ZN(n767) );
  NOR2_X1 U851 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U852 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U853 ( .A1(n772), .A2(n771), .ZN(n809) );
  NAND2_X1 U854 ( .A1(G129), .A2(n521), .ZN(n774) );
  NAND2_X1 U855 ( .A1(G117), .A2(n879), .ZN(n773) );
  NAND2_X1 U856 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U857 ( .A(KEYINPUT90), .B(n775), .ZN(n778) );
  NAND2_X1 U858 ( .A1(n882), .A2(G105), .ZN(n776) );
  XOR2_X1 U859 ( .A(KEYINPUT38), .B(n776), .Z(n777) );
  NOR2_X1 U860 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U861 ( .A1(G141), .A2(n883), .ZN(n779) );
  NAND2_X1 U862 ( .A1(n780), .A2(n779), .ZN(n889) );
  NAND2_X1 U863 ( .A1(n889), .A2(G1996), .ZN(n788) );
  NAND2_X1 U864 ( .A1(n521), .A2(G119), .ZN(n782) );
  NAND2_X1 U865 ( .A1(G131), .A2(n883), .ZN(n781) );
  NAND2_X1 U866 ( .A1(n782), .A2(n781), .ZN(n786) );
  NAND2_X1 U867 ( .A1(G95), .A2(n882), .ZN(n784) );
  NAND2_X1 U868 ( .A1(G107), .A2(n879), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n784), .A2(n783), .ZN(n785) );
  OR2_X1 U870 ( .A1(n786), .A2(n785), .ZN(n863) );
  NAND2_X1 U871 ( .A1(G1991), .A2(n863), .ZN(n787) );
  NAND2_X1 U872 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U873 ( .A(n789), .B(KEYINPUT91), .ZN(n920) );
  INV_X1 U874 ( .A(n920), .ZN(n792) );
  NOR2_X1 U875 ( .A1(n791), .A2(n790), .ZN(n821) );
  NAND2_X1 U876 ( .A1(n792), .A2(n821), .ZN(n810) );
  NAND2_X1 U877 ( .A1(n521), .A2(G128), .ZN(n793) );
  XOR2_X1 U878 ( .A(KEYINPUT89), .B(n793), .Z(n795) );
  NAND2_X1 U879 ( .A1(n879), .A2(G116), .ZN(n794) );
  NAND2_X1 U880 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U881 ( .A(KEYINPUT35), .B(n796), .Z(n803) );
  XOR2_X1 U882 ( .A(KEYINPUT88), .B(KEYINPUT34), .Z(n801) );
  NAND2_X1 U883 ( .A1(n882), .A2(G104), .ZN(n797) );
  XOR2_X1 U884 ( .A(KEYINPUT87), .B(n797), .Z(n799) );
  NAND2_X1 U885 ( .A1(G140), .A2(n883), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U887 ( .A(n801), .B(n800), .Z(n802) );
  NOR2_X1 U888 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U889 ( .A(KEYINPUT36), .B(n804), .ZN(n861) );
  XNOR2_X1 U890 ( .A(KEYINPUT37), .B(G2067), .ZN(n819) );
  NOR2_X1 U891 ( .A1(n861), .A2(n819), .ZN(n936) );
  NAND2_X1 U892 ( .A1(n821), .A2(n936), .ZN(n817) );
  AND2_X1 U893 ( .A1(n810), .A2(n817), .ZN(n807) );
  XNOR2_X1 U894 ( .A(G1986), .B(KEYINPUT86), .ZN(n805) );
  XNOR2_X1 U895 ( .A(n805), .B(G290), .ZN(n985) );
  NAND2_X1 U896 ( .A1(n985), .A2(n821), .ZN(n806) );
  AND2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U898 ( .A1(n809), .A2(n808), .ZN(n824) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n889), .ZN(n932) );
  INV_X1 U900 ( .A(n810), .ZN(n813) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n863), .ZN(n918) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n811) );
  NOR2_X1 U903 ( .A1(n918), .A2(n811), .ZN(n812) );
  NOR2_X1 U904 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U905 ( .A1(n932), .A2(n814), .ZN(n816) );
  XOR2_X1 U906 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n815) );
  XNOR2_X1 U907 ( .A(n816), .B(n815), .ZN(n818) );
  NAND2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n820) );
  NAND2_X1 U909 ( .A1(n861), .A2(n819), .ZN(n923) );
  NAND2_X1 U910 ( .A1(n820), .A2(n923), .ZN(n822) );
  NAND2_X1 U911 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U912 ( .A1(n824), .A2(n823), .ZN(n826) );
  XNOR2_X1 U913 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n825) );
  XNOR2_X1 U914 ( .A(n826), .B(n825), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n827), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U917 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U919 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U921 ( .A(G132), .ZN(G219) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G82), .ZN(G220) );
  INV_X1 U924 ( .A(G69), .ZN(G235) );
  NOR2_X1 U925 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  INV_X1 U927 ( .A(n833), .ZN(G319) );
  XNOR2_X1 U928 ( .A(G1981), .B(KEYINPUT41), .ZN(n843) );
  XOR2_X1 U929 ( .A(G1971), .B(G1966), .Z(n835) );
  XNOR2_X1 U930 ( .A(G1986), .B(G1976), .ZN(n834) );
  XNOR2_X1 U931 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U932 ( .A(G1956), .B(G1961), .Z(n837) );
  XNOR2_X1 U933 ( .A(G1996), .B(G1991), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U935 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U936 ( .A(G2474), .B(KEYINPUT108), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U938 ( .A(n843), .B(n842), .ZN(G229) );
  XOR2_X1 U939 ( .A(G2100), .B(G2096), .Z(n845) );
  XNOR2_X1 U940 ( .A(KEYINPUT42), .B(G2678), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U942 ( .A(KEYINPUT43), .B(G2090), .Z(n847) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U945 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U946 ( .A(G2084), .B(G2078), .ZN(n850) );
  XNOR2_X1 U947 ( .A(n851), .B(n850), .ZN(G227) );
  NAND2_X1 U948 ( .A1(G100), .A2(n882), .ZN(n853) );
  NAND2_X1 U949 ( .A1(G112), .A2(n879), .ZN(n852) );
  NAND2_X1 U950 ( .A1(n853), .A2(n852), .ZN(n859) );
  NAND2_X1 U951 ( .A1(n521), .A2(G124), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U953 ( .A1(G136), .A2(n883), .ZN(n855) );
  NAND2_X1 U954 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U955 ( .A(KEYINPUT109), .B(n857), .Z(n858) );
  NOR2_X1 U956 ( .A1(n859), .A2(n858), .ZN(G162) );
  XOR2_X1 U957 ( .A(G162), .B(n922), .Z(n860) );
  XNOR2_X1 U958 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U959 ( .A(G164), .B(G160), .Z(n862) );
  XNOR2_X1 U960 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U961 ( .A(n865), .B(n864), .Z(n870) );
  XOR2_X1 U962 ( .A(KEYINPUT110), .B(KEYINPUT112), .Z(n867) );
  XNOR2_X1 U963 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U965 ( .A(KEYINPUT46), .B(n868), .ZN(n869) );
  XNOR2_X1 U966 ( .A(n870), .B(n869), .ZN(n893) );
  NAND2_X1 U967 ( .A1(G127), .A2(n521), .ZN(n872) );
  NAND2_X1 U968 ( .A1(G115), .A2(n879), .ZN(n871) );
  NAND2_X1 U969 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U970 ( .A(n873), .B(KEYINPUT47), .ZN(n875) );
  NAND2_X1 U971 ( .A1(G103), .A2(n882), .ZN(n874) );
  NAND2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n878) );
  NAND2_X1 U973 ( .A1(G139), .A2(n883), .ZN(n876) );
  XNOR2_X1 U974 ( .A(KEYINPUT111), .B(n876), .ZN(n877) );
  NOR2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n925) );
  NAND2_X1 U976 ( .A1(G130), .A2(n521), .ZN(n881) );
  NAND2_X1 U977 ( .A1(G118), .A2(n879), .ZN(n880) );
  NAND2_X1 U978 ( .A1(n881), .A2(n880), .ZN(n888) );
  NAND2_X1 U979 ( .A1(n882), .A2(G106), .ZN(n885) );
  NAND2_X1 U980 ( .A1(G142), .A2(n883), .ZN(n884) );
  NAND2_X1 U981 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U982 ( .A(n886), .B(KEYINPUT45), .Z(n887) );
  NOR2_X1 U983 ( .A1(n888), .A2(n887), .ZN(n890) );
  XNOR2_X1 U984 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U985 ( .A(n925), .B(n891), .Z(n892) );
  XNOR2_X1 U986 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U987 ( .A1(G37), .A2(n894), .ZN(G395) );
  XOR2_X1 U988 ( .A(KEYINPUT114), .B(n895), .Z(n897) );
  XNOR2_X1 U989 ( .A(n970), .B(G286), .ZN(n896) );
  XNOR2_X1 U990 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U991 ( .A(G171), .B(n898), .ZN(n899) );
  NOR2_X1 U992 ( .A1(G37), .A2(n899), .ZN(G397) );
  XOR2_X1 U993 ( .A(G2454), .B(G2435), .Z(n901) );
  XNOR2_X1 U994 ( .A(G2438), .B(G2427), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n908) );
  XOR2_X1 U996 ( .A(KEYINPUT107), .B(G2446), .Z(n903) );
  XNOR2_X1 U997 ( .A(G2443), .B(G2430), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U999 ( .A(n904), .B(G2451), .Z(n906) );
  XNOR2_X1 U1000 ( .A(G1341), .B(G1348), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n909) );
  NAND2_X1 U1003 ( .A1(n909), .A2(G14), .ZN(n916) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n916), .ZN(n913) );
  NOR2_X1 U1005 ( .A1(G229), .A2(G227), .ZN(n910) );
  XOR2_X1 U1006 ( .A(KEYINPUT49), .B(n910), .Z(n911) );
  XNOR2_X1 U1007 ( .A(n911), .B(KEYINPUT115), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G96), .ZN(G221) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(n916), .ZN(G401) );
  XOR2_X1 U1015 ( .A(G160), .B(G2084), .Z(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n924) );
  NAND2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n930) );
  XOR2_X1 U1020 ( .A(G2072), .B(n925), .Z(n927) );
  XOR2_X1 U1021 ( .A(G164), .B(G2078), .Z(n926) );
  NOR2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1023 ( .A(KEYINPUT50), .B(n928), .Z(n929) );
  NOR2_X1 U1024 ( .A1(n930), .A2(n929), .ZN(n938) );
  XOR2_X1 U1025 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1027 ( .A(KEYINPUT51), .B(n933), .Z(n934) );
  XOR2_X1 U1028 ( .A(KEYINPUT116), .B(n934), .Z(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1030 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1031 ( .A(KEYINPUT52), .B(n939), .ZN(n940) );
  NAND2_X1 U1032 ( .A1(n940), .A2(G29), .ZN(n1023) );
  XNOR2_X1 U1033 ( .A(G2084), .B(G34), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n941), .B(KEYINPUT54), .ZN(n959) );
  XNOR2_X1 U1035 ( .A(G2090), .B(G35), .ZN(n956) );
  XNOR2_X1 U1036 ( .A(G2067), .B(G26), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(G33), .B(G2072), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n950) );
  XOR2_X1 U1039 ( .A(G1996), .B(G32), .Z(n944) );
  NAND2_X1 U1040 ( .A1(n944), .A2(G28), .ZN(n948) );
  XOR2_X1 U1041 ( .A(G27), .B(n945), .Z(n946) );
  XNOR2_X1 U1042 ( .A(KEYINPUT118), .B(n946), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n953) );
  XOR2_X1 U1045 ( .A(G25), .B(G1991), .Z(n951) );
  XNOR2_X1 U1046 ( .A(KEYINPUT117), .B(n951), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(KEYINPUT53), .B(n954), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(n957), .B(KEYINPUT119), .ZN(n958) );
  NOR2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(n960), .B(KEYINPUT120), .ZN(n961) );
  NOR2_X1 U1053 ( .A1(G29), .A2(n961), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(KEYINPUT55), .B(n962), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n963), .A2(G11), .ZN(n1021) );
  INV_X1 U1056 ( .A(G16), .ZN(n1017) );
  XNOR2_X1 U1057 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(n1017), .B(n964), .ZN(n992) );
  XOR2_X1 U1059 ( .A(G1966), .B(G168), .Z(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1061 ( .A(KEYINPUT57), .B(n967), .Z(n968) );
  XNOR2_X1 U1062 ( .A(KEYINPUT122), .B(n968), .ZN(n990) );
  XOR2_X1 U1063 ( .A(n969), .B(G1341), .Z(n988) );
  XNOR2_X1 U1064 ( .A(G171), .B(G1961), .ZN(n983) );
  XNOR2_X1 U1065 ( .A(n970), .B(G1348), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(n971), .B(KEYINPUT123), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(n972), .B(n998), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n981) );
  XNOR2_X1 U1069 ( .A(G1971), .B(G303), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(KEYINPUT124), .B(n979), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(KEYINPUT125), .B(n986), .ZN(n987) );
  NOR2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n1019) );
  XOR2_X1 U1080 ( .A(G1986), .B(G24), .Z(n994) );
  XOR2_X1 U1081 ( .A(G1971), .B(G22), .Z(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(G23), .B(G1976), .ZN(n995) );
  NOR2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1085 ( .A(KEYINPUT58), .B(n997), .Z(n1014) );
  XOR2_X1 U1086 ( .A(G1981), .B(G6), .Z(n1000) );
  XNOR2_X1 U1087 ( .A(n998), .B(G20), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1006) );
  XOR2_X1 U1089 ( .A(G1341), .B(G19), .Z(n1004) );
  XNOR2_X1 U1090 ( .A(KEYINPUT59), .B(G4), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(n1001), .B(KEYINPUT126), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(G1348), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(KEYINPUT60), .B(n1007), .ZN(n1009) );
  XOR2_X1 U1096 ( .A(G1961), .B(G5), .Z(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(G21), .B(G1966), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(KEYINPUT127), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1015), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1024), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

