//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n595,
    new_n596, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XOR2_X1   g020(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(KEYINPUT3), .A3(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n468), .A2(G137), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(new_n467), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(G101), .A3(new_n469), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n476));
  AND3_X1   g051(.A1(new_n471), .A2(new_n476), .A3(G125), .ZN(new_n477));
  AND2_X1   g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  OAI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n468), .A2(new_n471), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT71), .ZN(new_n485));
  INV_X1    g060(.A(G100), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n486), .A2(new_n469), .A3(KEYINPUT72), .ZN(new_n487));
  AOI21_X1  g062(.A(KEYINPUT72), .B1(new_n486), .B2(new_n469), .ZN(new_n488));
  OAI221_X1 g063(.A(G2104), .B1(G112), .B2(new_n469), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n482), .A2(new_n469), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  AND3_X1   g066(.A1(new_n485), .A2(new_n489), .A3(new_n491), .ZN(G162));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n468), .A2(new_n471), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT75), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT75), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n468), .A2(new_n497), .A3(new_n471), .A4(new_n494), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n471), .A2(new_n476), .ZN(new_n500));
  NOR4_X1   g075(.A1(new_n500), .A2(KEYINPUT4), .A3(new_n493), .A4(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n468), .A2(G126), .A3(G2105), .A4(new_n471), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT73), .A2(G114), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT73), .A2(G114), .ZN(new_n505));
  OAI21_X1  g080(.A(G2105), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(G102), .A2(G2105), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(G2104), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n503), .A2(new_n508), .A3(KEYINPUT74), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n499), .A2(new_n502), .B1(new_n511), .B2(new_n512), .ZN(G164));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT76), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT76), .A2(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT6), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n514), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT77), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT78), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT76), .B(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n518), .B1(new_n524), .B2(KEYINPUT6), .ZN(new_n525));
  AND2_X1   g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n523), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n517), .A2(new_n519), .ZN(new_n530));
  INV_X1    g105(.A(new_n528), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n530), .A2(KEYINPUT78), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(G88), .A3(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n531), .A2(G62), .ZN(new_n534));
  NAND2_X1  g109(.A1(G75), .A2(G543), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT79), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n524), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n522), .A2(new_n533), .A3(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  AND3_X1   g114(.A1(new_n529), .A2(G89), .A3(new_n532), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n520), .A2(G51), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n531), .A2(G63), .A3(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT80), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT7), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n544), .A2(new_n545), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n541), .B(new_n542), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n540), .A2(new_n548), .ZN(G168));
  NAND3_X1  g124(.A1(new_n529), .A2(G90), .A3(new_n532), .ZN(new_n550));
  XOR2_X1   g125(.A(KEYINPUT81), .B(G52), .Z(new_n551));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G64), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n528), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n520), .A2(new_n551), .B1(new_n554), .B2(new_n524), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT82), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT82), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n550), .A2(new_n558), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(G171));
  NAND3_X1  g135(.A1(new_n529), .A2(G81), .A3(new_n532), .ZN(new_n561));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G56), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n528), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n520), .A2(G43), .B1(new_n564), .B2(new_n524), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT83), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n561), .A2(new_n565), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT83), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n567), .A2(G860), .A3(new_n570), .ZN(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND4_X1  g149(.A1(G319), .A2(G483), .A3(G661), .A4(new_n574), .ZN(G188));
  INV_X1    g150(.A(G53), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT84), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n576), .B1(new_n577), .B2(KEYINPUT9), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n530), .A2(G543), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n577), .A2(KEYINPUT9), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n520), .B(new_n578), .C1(new_n577), .C2(KEYINPUT9), .ZN(new_n582));
  INV_X1    g157(.A(G65), .ZN(new_n583));
  OR2_X1    g158(.A1(KEYINPUT5), .A2(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(KEYINPUT5), .A2(G543), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n584), .A2(KEYINPUT85), .A3(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n587), .B1(new_n526), .B2(new_n527), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n583), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g164(.A1(G78), .A2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n581), .A2(new_n582), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n529), .A2(G91), .A3(new_n532), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G299));
  AND3_X1   g169(.A1(new_n550), .A2(new_n558), .A3(new_n555), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n558), .B1(new_n550), .B2(new_n555), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n595), .A2(new_n596), .ZN(G301));
  INV_X1    g172(.A(G168), .ZN(G286));
  NAND3_X1  g173(.A1(new_n529), .A2(G87), .A3(new_n532), .ZN(new_n599));
  INV_X1    g174(.A(G651), .ZN(new_n600));
  INV_X1    g175(.A(G74), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n600), .B1(new_n528), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(new_n520), .B2(G49), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(G288));
  NAND3_X1  g179(.A1(new_n529), .A2(G86), .A3(new_n532), .ZN(new_n605));
  NAND2_X1  g180(.A1(G73), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G61), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n528), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n520), .A2(G48), .B1(new_n608), .B2(new_n524), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(G305));
  NAND3_X1  g185(.A1(new_n529), .A2(G85), .A3(new_n532), .ZN(new_n611));
  NAND2_X1  g186(.A1(G72), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G60), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n528), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n520), .A2(G47), .B1(new_n614), .B2(new_n524), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(G290));
  AND2_X1   g191(.A1(G79), .A2(G543), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n586), .A2(new_n588), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G66), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(KEYINPUT86), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n600), .B1(new_n619), .B2(KEYINPUT86), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n620), .A2(new_n621), .B1(G54), .B2(new_n520), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n529), .A2(G92), .A3(new_n532), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT10), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g200(.A1(new_n529), .A2(KEYINPUT10), .A3(G92), .A4(new_n532), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(G868), .ZN(new_n629));
  MUX2_X1   g204(.A(G301), .B(new_n628), .S(new_n629), .Z(G284));
  MUX2_X1   g205(.A(G301), .B(new_n628), .S(new_n629), .Z(G321));
  NAND2_X1  g206(.A1(G299), .A2(new_n629), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n629), .B2(G168), .ZN(G297));
  OAI21_X1  g208(.A(new_n632), .B1(new_n629), .B2(G168), .ZN(G280));
  INV_X1    g209(.A(new_n628), .ZN(new_n635));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G860), .ZN(G148));
  NAND2_X1  g212(.A1(new_n567), .A2(new_n570), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(new_n629), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n628), .A2(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(new_n629), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g217(.A1(new_n473), .A2(new_n469), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n643), .A2(new_n500), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT12), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2100), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n483), .A2(G135), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n490), .A2(G123), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n469), .A2(G111), .ZN(new_n650));
  OAI21_X1  g225(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n648), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2096), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n647), .A2(new_n653), .ZN(G156));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT14), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2427), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2435), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n661), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n658), .B(new_n664), .Z(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  AND3_X1   g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT18), .Z(new_n675));
  INV_X1    g250(.A(new_n672), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n673), .B1(new_n676), .B2(new_n670), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT87), .B(KEYINPUT17), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n670), .B(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n677), .B1(new_n680), .B2(new_n676), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n676), .A3(new_n673), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n675), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2096), .B(G2100), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT88), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1956), .B(G2474), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1961), .B(G1966), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n687), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n688), .B2(new_n691), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT20), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n689), .A2(new_n690), .ZN(new_n695));
  INV_X1    g270(.A(new_n687), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n691), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n687), .A2(KEYINPUT89), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT91), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT90), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n703), .B(new_n707), .Z(G229));
  NAND2_X1  g283(.A1(new_n483), .A2(G131), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT92), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n469), .A2(G107), .ZN(new_n711));
  OAI21_X1  g286(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n490), .A2(G119), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G25), .B(new_n715), .S(G29), .Z(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT93), .Z(new_n717));
  XOR2_X1   g292(.A(KEYINPUT35), .B(G1991), .Z(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  MUX2_X1   g295(.A(G24), .B(G290), .S(G16), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1986), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G22), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G166), .B2(new_n724), .ZN(new_n726));
  INV_X1    g301(.A(G1971), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G6), .A2(G16), .ZN(new_n729));
  INV_X1    g304(.A(G305), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G16), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT32), .B(G1981), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n728), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G16), .A2(G23), .ZN(new_n735));
  NAND2_X1  g310(.A1(G288), .A2(KEYINPUT94), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT94), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n599), .A2(new_n737), .A3(new_n603), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n735), .B1(new_n739), .B2(G16), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT33), .B(G1976), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(KEYINPUT34), .B1(new_n734), .B2(new_n742), .ZN(new_n743));
  OR3_X1    g318(.A1(new_n734), .A2(new_n742), .A3(KEYINPUT34), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n717), .A2(new_n719), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n723), .A2(new_n743), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT36), .Z(new_n747));
  MUX2_X1   g322(.A(G19), .B(new_n638), .S(G16), .Z(new_n748));
  XOR2_X1   g323(.A(KEYINPUT95), .B(G1341), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n724), .A2(G4), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n635), .B2(new_n724), .ZN(new_n752));
  INV_X1    g327(.A(G1348), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G5), .A2(G16), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G171), .B2(G16), .ZN(new_n756));
  INV_X1    g331(.A(G1961), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n750), .A2(new_n754), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT24), .ZN(new_n760));
  INV_X1    g335(.A(G34), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n760), .B2(new_n761), .ZN(new_n763));
  INV_X1    g338(.A(G29), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(G160), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(G2084), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n483), .A2(G139), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT97), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  NAND2_X1  g345(.A1(G115), .A2(G2104), .ZN(new_n771));
  INV_X1    g346(.A(G127), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n500), .B2(new_n772), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n767), .B(new_n770), .C1(G2105), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G29), .ZN(new_n775));
  OR2_X1    g350(.A1(G29), .A2(G33), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT98), .B(G2072), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n766), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n779), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n777), .A2(new_n781), .B1(G2084), .B2(new_n765), .ZN(new_n782));
  NOR2_X1   g357(.A1(G164), .A2(new_n764), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G27), .B2(new_n764), .ZN(new_n784));
  INV_X1    g359(.A(G2078), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n780), .A2(new_n782), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n764), .A2(G32), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n483), .A2(G141), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n490), .A2(G129), .ZN(new_n791));
  INV_X1    g366(.A(new_n643), .ZN(new_n792));
  NAND3_X1  g367(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT26), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n792), .A2(G105), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n790), .A2(new_n791), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT99), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n789), .B1(new_n799), .B2(new_n764), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT27), .B(G1996), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT31), .B(G11), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT100), .B(G28), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n804), .A2(KEYINPUT30), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT101), .ZN(new_n806));
  AOI21_X1  g381(.A(G29), .B1(new_n804), .B2(KEYINPUT30), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n803), .B(new_n808), .C1(new_n652), .C2(new_n764), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT102), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n724), .A2(G21), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G168), .B2(new_n724), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1966), .ZN(new_n813));
  NOR4_X1   g388(.A1(new_n788), .A2(new_n802), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n724), .A2(G20), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT23), .Z(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G299), .B2(G16), .ZN(new_n817));
  INV_X1    g392(.A(G1956), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n764), .A2(G35), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G162), .B2(new_n764), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT29), .Z(new_n822));
  INV_X1    g397(.A(G2090), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n819), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n483), .A2(G140), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n490), .A2(G128), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n469), .A2(G116), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n826), .B(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G29), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n764), .A2(G26), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT28), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT96), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G2067), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n814), .A2(new_n824), .A3(new_n825), .A4(new_n836), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n747), .A2(new_n759), .A3(new_n837), .ZN(G311));
  INV_X1    g413(.A(G311), .ZN(G150));
  NAND3_X1  g414(.A1(new_n529), .A2(G93), .A3(new_n532), .ZN(new_n840));
  NAND2_X1  g415(.A1(G80), .A2(G543), .ZN(new_n841));
  INV_X1    g416(.A(G67), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n528), .B2(new_n842), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n520), .A2(G55), .B1(new_n843), .B2(new_n524), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n635), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n566), .A2(KEYINPUT103), .A3(new_n845), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT103), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n840), .A2(new_n844), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n851), .B1(new_n852), .B2(new_n568), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n567), .A2(new_n570), .A3(new_n845), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n849), .B(new_n856), .Z(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n859));
  INV_X1    g434(.A(G860), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n858), .B2(KEYINPUT39), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n847), .B1(new_n859), .B2(new_n861), .ZN(G145));
  XNOR2_X1  g437(.A(G162), .B(G160), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n652), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n715), .B(new_n645), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n483), .A2(G142), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n490), .A2(G130), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n469), .A2(G118), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n866), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n865), .B(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n871), .A2(new_n830), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n509), .B1(new_n499), .B2(new_n502), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n830), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n873), .B1(new_n872), .B2(new_n874), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n774), .A2(new_n798), .ZN(new_n878));
  INV_X1    g453(.A(new_n799), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n878), .B1(new_n774), .B2(new_n879), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n880), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n871), .B(new_n830), .ZN(new_n883));
  INV_X1    g458(.A(new_n873), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n882), .B1(new_n885), .B2(new_n875), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n864), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n880), .B1(new_n876), .B2(new_n877), .ZN(new_n889));
  INV_X1    g464(.A(new_n864), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n885), .A2(new_n875), .A3(new_n882), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g469(.A1(new_n845), .A2(new_n629), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n739), .A2(G290), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n739), .A2(G290), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n730), .A2(KEYINPUT105), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n730), .A2(KEYINPUT105), .ZN(new_n900));
  OAI21_X1  g475(.A(G166), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(G305), .B(KEYINPUT105), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(G303), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n896), .A2(new_n897), .B1(new_n901), .B2(new_n903), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT42), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n856), .B(new_n640), .Z(new_n909));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n581), .A2(new_n582), .A3(new_n591), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n529), .A2(G91), .A3(new_n532), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n592), .A2(KEYINPUT104), .A3(new_n593), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n635), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n628), .A2(new_n910), .A3(G299), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(KEYINPUT41), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n628), .A2(new_n910), .A3(G299), .ZN(new_n919));
  AND4_X1   g494(.A1(new_n627), .A2(new_n914), .A3(new_n622), .A4(new_n913), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n909), .A2(new_n917), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n919), .A2(new_n920), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(new_n909), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n908), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n895), .B1(new_n926), .B2(new_n629), .ZN(G295));
  OAI21_X1  g502(.A(new_n895), .B1(new_n926), .B2(new_n629), .ZN(G331));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT107), .B1(new_n595), .B2(new_n596), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n557), .A2(new_n932), .A3(new_n559), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n931), .A2(new_n933), .A3(G286), .ZN(new_n934));
  NAND3_X1  g509(.A1(G171), .A2(KEYINPUT107), .A3(G168), .ZN(new_n935));
  AND4_X1   g510(.A1(new_n855), .A2(new_n934), .A3(new_n854), .A4(new_n935), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n935), .A2(new_n934), .B1(new_n854), .B2(new_n855), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n923), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n935), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n856), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n934), .A2(new_n854), .A3(new_n855), .A4(new_n935), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n940), .A2(new_n921), .A3(new_n917), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n898), .B(new_n904), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n907), .A2(new_n938), .A3(new_n942), .ZN(new_n946));
  AND4_X1   g521(.A1(new_n930), .A2(new_n945), .A3(new_n888), .A4(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(G37), .B1(new_n943), .B2(new_n944), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n930), .B1(new_n948), .B2(new_n946), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT106), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT108), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n947), .B2(new_n949), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n929), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT44), .B1(new_n950), .B2(KEYINPUT108), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT109), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n951), .A2(new_n929), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n948), .A2(new_n946), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n948), .A2(new_n930), .A3(new_n946), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT108), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(KEYINPUT108), .B2(new_n950), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n957), .B(new_n958), .C1(new_n963), .C2(new_n929), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n956), .A2(new_n964), .ZN(G397));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n873), .B2(G1384), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n475), .A2(new_n968), .A3(G40), .A4(new_n479), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n479), .A2(G40), .A3(new_n474), .A4(new_n472), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT110), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n967), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G1996), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT46), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n830), .B(G2067), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT111), .ZN(new_n979));
  INV_X1    g554(.A(new_n798), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n974), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n977), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n983), .B(KEYINPUT126), .Z(new_n984));
  OR2_X1    g559(.A1(new_n984), .A2(KEYINPUT47), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(KEYINPUT47), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n798), .A2(G1996), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n979), .B(new_n987), .C1(G1996), .C2(new_n879), .ZN(new_n988));
  OR3_X1    g563(.A1(new_n988), .A2(new_n719), .A3(new_n715), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n830), .A2(G2067), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n982), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n715), .B(new_n719), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n982), .A2(G1986), .A3(G290), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n994), .A2(new_n974), .B1(KEYINPUT48), .B2(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n995), .A2(KEYINPUT48), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n991), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n985), .A2(new_n986), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n1000));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n501), .B1(new_n1002), .B2(new_n496), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1000), .B(new_n1001), .C1(new_n1003), .C2(new_n509), .ZN(new_n1004));
  AOI21_X1  g579(.A(G2090), .B1(new_n969), .B2(new_n971), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n511), .A2(new_n512), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n495), .A2(KEYINPUT75), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n502), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1384), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1004), .B(new_n1005), .C1(new_n1010), .C2(new_n1000), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT112), .ZN(new_n1012));
  OAI211_X1 g587(.A(KEYINPUT45), .B(new_n1001), .C1(new_n1003), .C2(new_n509), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n972), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT45), .B1(new_n1015), .B2(new_n1001), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n727), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1012), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT113), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1012), .A2(new_n1017), .A3(new_n1023), .A4(new_n1020), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1022), .A2(G8), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G303), .A2(G8), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1026), .B(KEYINPUT55), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  INV_X1    g605(.A(new_n509), .ZN(new_n1031));
  AOI21_X1  g606(.A(G1384), .B1(new_n1009), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1030), .B1(new_n1032), .B2(new_n972), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n736), .A2(G1976), .A3(new_n738), .ZN(new_n1034));
  INV_X1    g609(.A(G1976), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT52), .B1(G288), .B2(new_n1035), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1038), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1029), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT114), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G305), .A2(G1981), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(G305), .A2(KEYINPUT116), .A3(G1981), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT115), .B1(G305), .B2(G1981), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n1049));
  INV_X1    g624(.A(G1981), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n605), .A2(new_n1049), .A3(new_n1050), .A4(new_n609), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1046), .A2(new_n1047), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1033), .B1(new_n1052), .B2(KEYINPUT49), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1054), .A2(KEYINPUT49), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT117), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT49), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1052), .A2(KEYINPUT49), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1033), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1043), .B1(new_n1057), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1027), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1022), .A2(G8), .A3(new_n1065), .A4(new_n1024), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1010), .A2(KEYINPUT45), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n972), .A3(new_n967), .ZN(new_n1068));
  INV_X1    g643(.A(G1966), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G2084), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1018), .A2(new_n1071), .A3(new_n972), .A4(new_n1004), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1030), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT63), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1074), .A2(new_n1075), .A3(G286), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1028), .A2(new_n1064), .A3(new_n1066), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1010), .A2(new_n1000), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT50), .B1(new_n873), .B2(G1384), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(new_n972), .A3(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1017), .B1(G2090), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G8), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n1027), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1074), .A2(G286), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1064), .A2(new_n1066), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1075), .B1(new_n1085), .B2(KEYINPUT119), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1043), .ZN(new_n1089));
  AND4_X1   g664(.A1(new_n1066), .A2(new_n1088), .A3(new_n1083), .A4(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1087), .B1(new_n1090), .B2(new_n1084), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1077), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n599), .A2(new_n1035), .A3(new_n603), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(new_n1057), .B2(new_n1063), .ZN(new_n1095));
  XOR2_X1   g670(.A(new_n1055), .B(KEYINPUT118), .Z(new_n1096));
  OAI21_X1  g671(.A(new_n1033), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1064), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1066), .B2(new_n1098), .ZN(new_n1099));
  XOR2_X1   g674(.A(G299), .B(KEYINPUT57), .Z(new_n1100));
  NAND2_X1  g675(.A1(new_n1080), .A2(new_n818), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1013), .A2(new_n972), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1016), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT56), .B(G2072), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1100), .A2(new_n1101), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1100), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT120), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT61), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1102), .A2(new_n1103), .A3(new_n975), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1032), .A2(new_n972), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT58), .B(G1341), .Z(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n638), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1114), .A2(KEYINPUT59), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1018), .A2(new_n972), .A3(new_n1004), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n753), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1111), .A2(G2067), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n628), .A2(KEYINPUT60), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n1114), .B2(KEYINPUT59), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1115), .A2(new_n1121), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1117), .A2(new_n628), .A3(new_n1118), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n628), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT60), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  OAI211_X1 g701(.A(KEYINPUT120), .B(new_n1126), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1109), .A2(new_n1122), .A3(new_n1125), .A4(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1106), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1107), .B1(new_n1129), .B2(new_n1124), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1102), .A2(new_n1103), .A3(new_n785), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1132), .A2(new_n1133), .B1(new_n757), .B2(new_n1116), .ZN(new_n1134));
  OR3_X1    g709(.A1(new_n1068), .A2(new_n1133), .A3(G2078), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n1137));
  XNOR2_X1  g712(.A(G171), .B(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n475), .B(KEYINPUT122), .ZN(new_n1139));
  OAI211_X1 g714(.A(KEYINPUT53), .B(G40), .C1(KEYINPUT123), .C2(G2078), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(KEYINPUT123), .B2(G2078), .ZN(new_n1141));
  AND4_X1   g716(.A1(new_n479), .A2(new_n967), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1138), .B1(new_n1013), .B2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1136), .A2(new_n1138), .B1(new_n1143), .B2(new_n1134), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G168), .A2(new_n1030), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT121), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1148), .B(KEYINPUT51), .C1(new_n1073), .C2(new_n1147), .ZN(new_n1149));
  OR3_X1    g724(.A1(new_n1073), .A2(KEYINPUT51), .A3(new_n1147), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1144), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1064), .A2(new_n1066), .A3(new_n1083), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1099), .B1(new_n1131), .B2(new_n1153), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1092), .A2(new_n1093), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1093), .B1(new_n1092), .B2(new_n1154), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1150), .A2(new_n1149), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1136), .A2(G171), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1150), .A2(new_n1149), .A3(KEYINPUT125), .A4(KEYINPUT62), .ZN(new_n1163));
  AND4_X1   g738(.A1(new_n1090), .A2(new_n1160), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1155), .A2(new_n1156), .A3(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(G290), .B(G1986), .Z(new_n1166));
  AOI21_X1  g741(.A(new_n982), .B1(new_n993), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n999), .B1(new_n1165), .B2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g743(.A1(G227), .A2(new_n462), .ZN(new_n1170));
  XNOR2_X1  g744(.A(new_n1170), .B(KEYINPUT127), .ZN(new_n1171));
  OR3_X1    g745(.A1(G229), .A2(G401), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g746(.A(new_n1172), .ZN(new_n1173));
  OAI211_X1 g747(.A(new_n893), .B(new_n1173), .C1(new_n949), .C2(new_n947), .ZN(G225));
  INV_X1    g748(.A(G225), .ZN(G308));
endmodule


