//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1180, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1228, new_n1229, new_n1230, new_n1231;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT64), .Z(new_n208));
  INV_X1    g0008(.A(G58), .ZN(new_n209));
  INV_X1    g0009(.A(G232), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G50), .B2(G226), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n208), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n206), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n206), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  NOR3_X1   g0028(.A1(new_n221), .A2(new_n225), .A3(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(new_n210), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G1698), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G257), .ZN(new_n246));
  AND2_X1   g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  OAI221_X1 g0048(.A(new_n246), .B1(new_n212), .B2(new_n245), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n247), .A2(new_n248), .ZN(new_n250));
  INV_X1    g0050(.A(G303), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  OAI211_X1 g0054(.A(G1), .B(G13), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n249), .A2(new_n252), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT5), .B(G41), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G1), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G270), .A3(new_n255), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n258), .A2(G274), .A3(new_n260), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n257), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT76), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G116), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n266), .A2(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n267), .A2(new_n271), .A3(new_n224), .A4(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n272), .A2(new_n224), .B1(G20), .B2(new_n269), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G283), .ZN(new_n275));
  INV_X1    g0075(.A(G97), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n275), .B(new_n223), .C1(G33), .C2(new_n276), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n274), .A2(KEYINPUT20), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(KEYINPUT20), .B1(new_n274), .B2(new_n277), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n270), .B1(new_n269), .B2(new_n273), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT76), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n257), .A2(new_n262), .A3(new_n281), .A4(new_n263), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n265), .A2(new_n280), .A3(G169), .A4(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT77), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(KEYINPUT21), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n283), .A2(new_n285), .ZN(new_n287));
  INV_X1    g0087(.A(G179), .ZN(new_n288));
  OR2_X1    g0088(.A1(new_n264), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n280), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n286), .A2(new_n287), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n211), .A2(G20), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT23), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n223), .B(G87), .C1(new_n247), .C2(new_n248), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT22), .ZN(new_n296));
  OR2_X1    g0096(.A1(KEYINPUT3), .A2(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(KEYINPUT3), .A2(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT22), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n299), .A2(new_n300), .A3(new_n223), .A4(G87), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n294), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n223), .A2(G33), .A3(G116), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT78), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT24), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n272), .A2(new_n224), .ZN(new_n308));
  NAND2_X1  g0108(.A1(KEYINPUT78), .A2(KEYINPUT24), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n305), .A2(new_n306), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n302), .A2(new_n303), .A3(new_n309), .A4(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n307), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n266), .A2(G13), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT25), .B1(new_n313), .B2(new_n293), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n313), .A2(new_n293), .A3(KEYINPUT25), .ZN(new_n315));
  INV_X1    g0115(.A(new_n308), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT71), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(new_n271), .A4(new_n267), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n273), .A2(KEYINPUT71), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n315), .B1(new_n320), .B2(G107), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n312), .A2(new_n314), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n245), .B1(new_n297), .B2(new_n298), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT80), .B(G294), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n323), .A2(G257), .B1(new_n324), .B2(G33), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT79), .ZN(new_n326));
  OAI21_X1  g0126(.A(G250), .B1(new_n247), .B2(new_n248), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n326), .B1(new_n327), .B2(G1698), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n299), .A2(KEYINPUT79), .A3(G250), .A4(new_n245), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n325), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT81), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n325), .A2(KEYINPUT81), .A3(new_n328), .A4(new_n329), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(new_n256), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n256), .B1(new_n260), .B2(new_n258), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G264), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n263), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G169), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n334), .A2(new_n288), .A3(new_n263), .A4(new_n336), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n322), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n292), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G223), .A2(G1698), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n245), .A2(G222), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n299), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n345), .B(new_n256), .C1(G77), .C2(new_n299), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n347));
  INV_X1    g0147(.A(G274), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n255), .A2(new_n347), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G226), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n346), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G190), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n267), .A2(G50), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n316), .B1(G1), .B2(new_n223), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n202), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n203), .A2(G20), .ZN(new_n360));
  INV_X1    g0160(.A(G150), .ZN(new_n361));
  NOR2_X1   g0161(.A1(G20), .A2(G33), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(KEYINPUT65), .A2(G58), .ZN(new_n364));
  XOR2_X1   g0164(.A(new_n364), .B(KEYINPUT8), .Z(new_n365));
  NAND2_X1  g0165(.A1(new_n223), .A2(G33), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n360), .B1(new_n361), .B2(new_n363), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  AOI211_X1 g0167(.A(new_n357), .B(new_n359), .C1(new_n367), .C2(new_n308), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n356), .B1(new_n368), .B2(KEYINPUT9), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n354), .A2(G200), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n369), .B(new_n370), .C1(KEYINPUT9), .C2(new_n368), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT10), .ZN(new_n372));
  INV_X1    g0172(.A(new_n368), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n354), .A2(new_n338), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n373), .B(new_n374), .C1(G179), .C2(new_n354), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G238), .A2(G1698), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n299), .B(new_n377), .C1(new_n210), .C2(G1698), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n378), .B(new_n256), .C1(G107), .C2(new_n299), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n352), .A2(G244), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(new_n350), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n381), .A2(new_n355), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G20), .A2(G77), .ZN(new_n386));
  XNOR2_X1  g0186(.A(KEYINPUT15), .B(G87), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT8), .B(G58), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n386), .B1(new_n387), .B2(new_n366), .C1(new_n363), .C2(new_n388), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(new_n308), .B1(new_n217), .B2(new_n268), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n358), .A2(new_n217), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n384), .A2(new_n385), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT13), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n210), .A2(G1698), .ZN(new_n395));
  OAI221_X1 g0195(.A(new_n395), .B1(G226), .B2(G1698), .C1(new_n247), .C2(new_n248), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G33), .A2(G97), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n255), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n398), .A2(new_n349), .ZN(new_n399));
  INV_X1    g0199(.A(G238), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n351), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n394), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  NOR4_X1   g0203(.A1(new_n398), .A2(new_n401), .A3(KEYINPUT13), .A4(new_n349), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT66), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n399), .A2(new_n402), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(KEYINPUT66), .A3(KEYINPUT13), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(G190), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G68), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G20), .ZN(new_n411));
  OAI221_X1 g0211(.A(new_n411), .B1(new_n366), .B2(new_n217), .C1(new_n363), .C2(new_n202), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n412), .A2(KEYINPUT11), .A3(new_n308), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n410), .B2(new_n358), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n313), .A2(new_n411), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT12), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT11), .B1(new_n412), .B2(new_n308), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n406), .A2(KEYINPUT13), .ZN(new_n419));
  INV_X1    g0219(.A(new_n404), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G200), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n409), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT67), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT67), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n409), .A2(new_n425), .A3(new_n418), .A4(new_n422), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n382), .A2(new_n288), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n381), .A2(new_n338), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n428), .A3(new_n392), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n424), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  OR3_X1    g0230(.A1(new_n376), .A2(new_n393), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT66), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n419), .A2(new_n432), .A3(new_n420), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n288), .B1(new_n433), .B2(new_n407), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT14), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n421), .B2(G169), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n435), .B(G169), .C1(new_n403), .C2(new_n404), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  OR3_X1    g0238(.A1(new_n434), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n418), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n299), .B1(G226), .B2(new_n245), .ZN(new_n442));
  NOR2_X1   g0242(.A1(G223), .A2(G1698), .ZN(new_n443));
  INV_X1    g0243(.A(G87), .ZN(new_n444));
  OAI22_X1  g0244(.A1(new_n442), .A2(new_n443), .B1(new_n253), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n349), .B1(new_n445), .B2(new_n256), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n351), .A2(new_n210), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(G169), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT7), .B1(new_n250), .B2(new_n223), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT7), .ZN(new_n451));
  NOR4_X1   g0251(.A1(new_n247), .A2(new_n248), .A3(new_n451), .A4(G20), .ZN(new_n452));
  OAI21_X1  g0252(.A(G68), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n209), .A2(new_n410), .ZN(new_n454));
  OAI21_X1  g0254(.A(G20), .B1(new_n454), .B2(new_n201), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n362), .A2(G159), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT16), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n316), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT68), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n297), .A2(new_n223), .A3(new_n298), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n451), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n297), .A2(KEYINPUT7), .A3(new_n223), .A4(new_n298), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n457), .B1(new_n466), .B2(G68), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n462), .B1(new_n467), .B2(KEYINPUT16), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n410), .B1(new_n464), .B2(new_n465), .ZN(new_n469));
  NOR4_X1   g0269(.A1(new_n469), .A2(KEYINPUT68), .A3(new_n457), .A4(new_n460), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n461), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n365), .A2(new_n268), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n365), .B2(new_n358), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n449), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  AOI211_X1 g0275(.A(new_n447), .B(new_n349), .C1(new_n445), .C2(new_n256), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n288), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT18), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n475), .A2(KEYINPUT18), .A3(new_n477), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n446), .A2(new_n355), .A3(new_n448), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n476), .B2(G200), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT69), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n484), .A2(new_n471), .A3(new_n485), .A4(new_n474), .ZN(new_n486));
  XNOR2_X1  g0286(.A(new_n486), .B(KEYINPUT17), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n441), .A2(new_n482), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n431), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n334), .A2(new_n355), .A3(new_n263), .A4(new_n336), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n337), .A2(new_n383), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n322), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(G244), .B1(new_n247), .B2(new_n248), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n494), .A2(G1698), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n496), .B(G244), .C1(new_n248), .C2(new_n247), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n275), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n245), .B1(new_n327), .B2(KEYINPUT4), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT72), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n327), .A2(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G1698), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n493), .A2(new_n494), .B1(G33), .B2(G283), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT72), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .A4(new_n497), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n500), .A2(new_n505), .A3(new_n256), .ZN(new_n506));
  INV_X1    g0306(.A(new_n263), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n507), .B1(new_n335), .B2(G257), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G200), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n320), .A2(G97), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n268), .A2(new_n276), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g0313(.A1(KEYINPUT6), .A2(G97), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT6), .B1(G97), .B2(G107), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT70), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n516), .B1(new_n514), .B2(new_n515), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n211), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n514), .A2(new_n515), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT70), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(G107), .A3(new_n517), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n523), .A3(G20), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n466), .A2(G107), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n362), .A2(G77), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n513), .B1(new_n527), .B2(new_n308), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n506), .A2(G190), .A3(new_n508), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n510), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n509), .A2(new_n338), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n308), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n511), .A2(new_n512), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n506), .A2(new_n288), .A3(new_n508), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n492), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n245), .A2(G238), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G244), .A2(G1698), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n297), .A2(new_n298), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n253), .A2(new_n269), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n256), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n266), .A2(G45), .ZN(new_n544));
  AND2_X1   g0344(.A1(G33), .A2(G41), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n544), .B(G250), .C1(new_n545), .C2(new_n224), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n260), .A2(G274), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT73), .B1(new_n543), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n400), .A2(G1698), .ZN(new_n551));
  AND2_X1   g0351(.A1(G244), .A2(G1698), .ZN(new_n552));
  OAI22_X1  g0352(.A1(new_n551), .A2(new_n552), .B1(new_n247), .B2(new_n248), .ZN(new_n553));
  INV_X1    g0353(.A(new_n542), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n255), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT73), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n555), .A2(new_n556), .A3(new_n548), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n288), .B1(new_n550), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n555), .B2(new_n548), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n543), .A2(new_n549), .A3(KEYINPUT73), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n560), .A3(new_n338), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT74), .ZN(new_n562));
  XOR2_X1   g0362(.A(KEYINPUT15), .B(G87), .Z(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(new_n267), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n444), .A2(new_n276), .A3(new_n211), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n397), .A2(new_n223), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT19), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n223), .B(G68), .C1(new_n247), .C2(new_n248), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT19), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n366), .B2(new_n276), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n564), .B1(new_n571), .B2(new_n308), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n318), .A2(new_n319), .A3(new_n563), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n562), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n572), .A2(new_n562), .A3(new_n573), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n558), .B(new_n561), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(G190), .B1(new_n550), .B2(new_n557), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n318), .A2(new_n319), .A3(G87), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n559), .A2(new_n560), .A3(G200), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n577), .A2(new_n572), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT75), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n576), .A2(new_n580), .A3(KEYINPUT75), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n265), .A2(new_n282), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n280), .B1(new_n585), .B2(G190), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n383), .B2(new_n585), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n583), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  AND4_X1   g0388(.A1(new_n342), .A2(new_n489), .A3(new_n538), .A4(new_n588), .ZN(G372));
  NAND2_X1  g0389(.A1(new_n292), .A2(new_n341), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n572), .A2(new_n573), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n543), .A2(new_n549), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n338), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n558), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(G200), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n577), .A2(new_n595), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n572), .A2(KEYINPUT82), .A3(new_n578), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT82), .B1(new_n572), .B2(new_n578), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n594), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n538), .A2(new_n590), .A3(new_n601), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n531), .A2(new_n535), .A3(new_n534), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n583), .A2(new_n603), .A3(new_n584), .ZN(new_n604));
  XOR2_X1   g0404(.A(KEYINPUT83), .B(KEYINPUT26), .Z(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n536), .A2(new_n600), .ZN(new_n607));
  OAI22_X1  g0407(.A1(new_n604), .A2(new_n606), .B1(KEYINPUT26), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n602), .A2(new_n608), .A3(new_n594), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n489), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n482), .ZN(new_n611));
  INV_X1    g0411(.A(new_n429), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n439), .A2(new_n440), .B1(new_n423), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n611), .B1(new_n614), .B2(new_n487), .ZN(new_n615));
  INV_X1    g0415(.A(new_n372), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n375), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n610), .A2(new_n618), .ZN(G369));
  INV_X1    g0419(.A(G13), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n620), .A2(G20), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n266), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n622), .A2(KEYINPUT27), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(KEYINPUT27), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(G213), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(G343), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n280), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g0428(.A(new_n292), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n587), .ZN(new_n630));
  INV_X1    g0430(.A(G330), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n322), .A2(new_n627), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n341), .B1(new_n492), .B2(new_n634), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n341), .A2(new_n627), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n292), .A2(new_n627), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n635), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n641), .A2(new_n636), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n639), .A2(new_n642), .ZN(G399));
  NOR2_X1   g0443(.A1(new_n565), .A2(G116), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n226), .A2(new_n254), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(G1), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n222), .B2(new_n645), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(KEYINPUT28), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT29), .ZN(new_n649));
  INV_X1    g0449(.A(new_n627), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n609), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n536), .A2(new_n600), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n576), .A2(KEYINPUT75), .A3(new_n580), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT75), .B1(new_n576), .B2(new_n580), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n655), .A2(new_n656), .A3(new_n536), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n654), .B1(new_n657), .B2(new_n605), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT84), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(new_n594), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n653), .B1(new_n604), .B2(new_n606), .ZN(new_n661));
  INV_X1    g0461(.A(new_n594), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT84), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n660), .A2(new_n663), .A3(new_n602), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n650), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n651), .B1(new_n665), .B2(KEYINPUT29), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n538), .A2(new_n588), .A3(new_n342), .A4(new_n650), .ZN(new_n667));
  INV_X1    g0467(.A(new_n509), .ZN(new_n668));
  AOI211_X1 g0468(.A(new_n288), .B(new_n264), .C1(new_n559), .C2(new_n560), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n668), .A2(new_n669), .A3(new_n336), .A4(new_n334), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT30), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n668), .A2(new_n585), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(new_n288), .A3(new_n337), .A4(new_n592), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n627), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n667), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT31), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n676), .A2(new_n679), .A3(new_n627), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G330), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n666), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n648), .B1(new_n683), .B2(G1), .ZN(G364));
  NAND2_X1  g0484(.A1(new_n621), .A2(G45), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n645), .A2(G1), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n632), .B(KEYINPUT85), .ZN(new_n687));
  INV_X1    g0487(.A(new_n630), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n686), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n224), .B1(G20), .B2(new_n338), .ZN(new_n691));
  NAND3_X1  g0491(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G190), .ZN(new_n693));
  INV_X1    g0493(.A(G317), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT33), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT33), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n692), .A2(new_n355), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G326), .ZN(new_n699));
  INV_X1    g0499(.A(new_n324), .ZN(new_n700));
  NOR2_X1   g0500(.A1(G179), .A2(G200), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n223), .B1(new_n701), .B2(G190), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n697), .B(new_n699), .C1(new_n700), .C2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n223), .A2(new_n355), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n288), .A2(G200), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(KEYINPUT87), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n706), .A2(KEYINPUT87), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT89), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n383), .A2(G179), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n704), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n299), .B1(new_n715), .B2(G303), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n711), .A2(G322), .B1(new_n712), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n223), .A2(G190), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n705), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n718), .A2(new_n701), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI22_X1  g0522(.A1(G311), .A2(new_n720), .B1(new_n722), .B2(G329), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n717), .B(new_n723), .C1(new_n712), .C2(new_n716), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n713), .A2(new_n718), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI211_X1 g0526(.A(new_n703), .B(new_n724), .C1(G283), .C2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G159), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n721), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g0529(.A(KEYINPUT88), .B(KEYINPUT32), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n729), .B(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n250), .B1(new_n726), .B2(G107), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n731), .B(new_n732), .C1(new_n217), .C2(new_n719), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n714), .A2(new_n444), .ZN(new_n734));
  INV_X1    g0534(.A(new_n702), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n735), .A2(G97), .B1(G50), .B2(new_n698), .ZN(new_n736));
  INV_X1    g0536(.A(new_n693), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n736), .B1(new_n410), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n710), .A2(new_n209), .ZN(new_n739));
  NOR4_X1   g0539(.A1(new_n733), .A2(new_n734), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n691), .B1(new_n727), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n299), .A2(G355), .A3(new_n226), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n250), .A2(new_n226), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT86), .Z(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(G45), .B2(new_n222), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n240), .A2(new_n259), .ZN(new_n746));
  OAI221_X1 g0546(.A(new_n742), .B1(G116), .B2(new_n226), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n691), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n750), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n741), .B(new_n752), .C1(new_n688), .C2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n686), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n690), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT90), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n757), .B(new_n758), .ZN(G396));
  NAND2_X1  g0559(.A1(new_n429), .A2(KEYINPUT95), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT95), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n427), .A2(new_n428), .A3(new_n761), .A4(new_n392), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n393), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n609), .A2(new_n650), .A3(new_n763), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n609), .A2(new_n650), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n392), .A2(new_n627), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n612), .A2(new_n627), .ZN(new_n768));
  AND3_X1   g0568(.A1(new_n767), .A2(KEYINPUT96), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(KEYINPUT96), .B1(new_n767), .B2(new_n768), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n764), .B1(new_n765), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n682), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n774), .A2(KEYINPUT97), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(KEYINPUT97), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n772), .A2(new_n682), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n775), .A2(new_n686), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G132), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n299), .B1(new_n721), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT94), .Z(new_n781));
  OAI22_X1  g0581(.A1(new_n714), .A2(new_n202), .B1(new_n702), .B2(new_n209), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n693), .A2(G150), .B1(new_n698), .B2(G137), .ZN(new_n783));
  INV_X1    g0583(.A(G143), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n783), .B1(new_n728), .B2(new_n719), .C1(new_n710), .C2(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT93), .Z(new_n786));
  AOI211_X1 g0586(.A(new_n781), .B(new_n782), .C1(new_n786), .C2(KEYINPUT34), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n787), .B1(KEYINPUT34), .B2(new_n786), .C1(new_n410), .C2(new_n725), .ZN(new_n788));
  INV_X1    g0588(.A(G283), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n737), .A2(new_n789), .B1(new_n719), .B2(new_n269), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT91), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  INV_X1    g0593(.A(new_n698), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n792), .B(new_n793), .C1(new_n251), .C2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT92), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n711), .A2(G294), .B1(G97), .B2(new_n735), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n250), .B1(new_n721), .B2(new_n798), .C1(new_n211), .C2(new_n714), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(G87), .B2(new_n726), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n796), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n788), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n691), .A2(new_n748), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n802), .A2(new_n691), .B1(new_n217), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n767), .A2(new_n768), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n804), .B(new_n755), .C1(new_n749), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n778), .A2(new_n806), .ZN(G384));
  NAND2_X1  g0607(.A1(new_n471), .A2(new_n474), .ZN(new_n808));
  INV_X1    g0608(.A(new_n625), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n484), .A2(new_n471), .A3(new_n474), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n449), .ZN(new_n813));
  AND3_X1   g0613(.A1(new_n808), .A2(new_n813), .A3(new_n477), .ZN(new_n814));
  OAI21_X1  g0614(.A(KEYINPUT37), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT17), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n486), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n808), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n818), .A2(new_n485), .A3(KEYINPUT17), .A4(new_n484), .ZN(new_n819));
  AND4_X1   g0619(.A1(KEYINPUT18), .A2(new_n808), .A3(new_n813), .A4(new_n477), .ZN(new_n820));
  AOI21_X1  g0620(.A(KEYINPUT18), .B1(new_n475), .B2(new_n477), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n817), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n810), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n815), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n812), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n478), .A2(KEYINPUT99), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT37), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n478), .B2(KEYINPUT99), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(KEYINPUT38), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n478), .A2(KEYINPUT99), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n832), .A2(new_n828), .A3(new_n825), .A4(new_n826), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT38), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n810), .B1(new_n482), .B2(new_n487), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n833), .B(new_n834), .C1(new_n835), .C2(new_n815), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT100), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n831), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(KEYINPUT101), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT101), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n831), .A2(new_n836), .A3(new_n841), .A4(new_n838), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n441), .A2(new_n627), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n840), .A2(new_n844), .A3(new_n842), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n418), .A2(new_n650), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n441), .A2(new_n423), .A3(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n434), .A2(new_n436), .A3(new_n438), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n424), .A2(new_n854), .A3(new_n426), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n850), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT98), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT98), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n855), .A2(new_n858), .A3(new_n850), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n853), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n760), .A2(new_n650), .A3(new_n762), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n860), .B1(new_n764), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n831), .A2(new_n836), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n862), .A2(new_n863), .B1(new_n611), .B2(new_n625), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n849), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT102), .ZN(new_n866));
  INV_X1    g0666(.A(new_n489), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n866), .B1(new_n666), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n649), .B1(new_n664), .B2(new_n650), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n489), .B(KEYINPUT102), .C1(new_n869), .C2(new_n651), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n618), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n865), .B(new_n872), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n678), .A2(new_n680), .A3(new_n805), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n855), .A2(new_n858), .A3(new_n850), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n858), .B1(new_n855), .B2(new_n850), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n852), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n874), .A2(new_n863), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT40), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n874), .A2(new_n863), .A3(KEYINPUT40), .A4(new_n877), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n489), .A2(new_n681), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n882), .B(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n884), .A2(new_n631), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n873), .B(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n266), .B2(new_n621), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n520), .A2(new_n523), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT35), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n223), .B(new_n224), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n890), .B(G116), .C1(new_n889), .C2(new_n888), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT36), .ZN(new_n892));
  OAI21_X1  g0692(.A(G77), .B1(new_n209), .B2(new_n410), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n893), .A2(new_n222), .B1(G50), .B2(new_n410), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(G1), .A3(new_n620), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n887), .A2(new_n892), .A3(new_n895), .ZN(G367));
  NOR2_X1   g0696(.A1(new_n714), .A2(new_n269), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT46), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(G107), .B2(new_n735), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n720), .A2(G283), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n711), .A2(G303), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n250), .B1(new_n721), .B2(new_n694), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n700), .A2(new_n737), .B1(new_n794), .B2(new_n798), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n902), .B(new_n903), .C1(G97), .C2(new_n726), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n899), .A2(new_n900), .A3(new_n901), .A4(new_n904), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n735), .A2(G68), .B1(G143), .B2(new_n698), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n217), .B2(new_n725), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n720), .A2(G50), .B1(G159), .B2(new_n693), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(KEYINPUT108), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n908), .A2(KEYINPUT108), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(new_n250), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n909), .B(new_n911), .C1(new_n361), .C2(new_n710), .ZN(new_n912));
  AOI22_X1  g0712(.A1(G58), .A2(new_n715), .B1(new_n722), .B2(G137), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT109), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n905), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT110), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT47), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n686), .B1(new_n917), .B2(new_n691), .ZN(new_n918));
  INV_X1    g0718(.A(new_n744), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n751), .B1(new_n226), .B2(new_n387), .C1(new_n919), .C2(new_n236), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n599), .A2(new_n627), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n601), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n594), .B2(new_n921), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n918), .B(new_n920), .C1(new_n753), .C2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n528), .A2(new_n650), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n537), .A2(new_n926), .B1(new_n536), .B2(new_n650), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT103), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n928), .A2(new_n641), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT42), .Z(new_n930));
  OR2_X1    g0730(.A1(new_n928), .A2(new_n341), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n627), .B1(new_n931), .B2(new_n536), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n925), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n927), .B(KEYINPUT103), .Z(new_n934));
  NAND2_X1  g0734(.A1(new_n638), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n933), .A2(new_n936), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n938), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n940), .B1(new_n938), .B2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n685), .A2(G1), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT106), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n641), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n637), .B1(new_n292), .B2(new_n627), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n641), .A2(new_n946), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n687), .B2(KEYINPUT107), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT107), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n633), .B1(new_n687), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n951), .B1(new_n953), .B2(new_n950), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n683), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n934), .A2(new_n642), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT44), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n934), .A2(new_n642), .ZN(new_n959));
  XOR2_X1   g0759(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n639), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n958), .A2(new_n961), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n638), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n956), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n683), .ZN(new_n966));
  XOR2_X1   g0766(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n967));
  XNOR2_X1  g0767(.A(new_n645), .B(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n945), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n924), .B1(new_n944), .B2(new_n969), .ZN(G387));
  AND2_X1   g0770(.A1(new_n722), .A2(G326), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n693), .A2(G311), .B1(new_n698), .B2(G322), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n251), .B2(new_n719), .C1(new_n710), .C2(new_n694), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT48), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n974), .B1(new_n789), .B2(new_n702), .C1(new_n700), .C2(new_n714), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n299), .B(new_n971), .C1(new_n976), .C2(KEYINPUT49), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n977), .B1(KEYINPUT49), .B2(new_n976), .C1(new_n269), .C2(new_n725), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n721), .A2(new_n361), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n714), .A2(new_n217), .B1(new_n719), .B2(new_n410), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(new_n711), .B2(G50), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n365), .A2(new_n737), .B1(new_n794), .B2(new_n728), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n702), .A2(new_n387), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n250), .B1(new_n726), .B2(G97), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n981), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n978), .B1(new_n979), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n691), .ZN(new_n988));
  INV_X1    g0788(.A(new_n644), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n388), .A2(G50), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n989), .B1(new_n991), .B2(KEYINPUT50), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n992), .B(new_n259), .C1(KEYINPUT50), .C2(new_n991), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n410), .A2(new_n217), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n744), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT111), .Z(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G45), .B2(new_n233), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n989), .A2(new_n226), .A3(new_n299), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(G107), .B2(new_n226), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n751), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n988), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n637), .B2(new_n750), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n1002), .A2(new_n755), .B1(new_n945), .B2(new_n954), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n645), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n954), .B2(new_n683), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1003), .B1(new_n956), .B2(new_n1005), .ZN(G393));
  NAND2_X1  g0806(.A1(new_n964), .A2(new_n962), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n645), .B1(new_n1007), .B2(new_n955), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n965), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n964), .A2(new_n945), .A3(new_n962), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT113), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n751), .B1(new_n276), .B2(new_n226), .C1(new_n919), .C2(new_n243), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n710), .A2(new_n798), .B1(new_n694), .B2(new_n794), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT52), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n722), .A2(G322), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n737), .A2(new_n251), .B1(new_n725), .B2(new_n211), .ZN(new_n1016));
  INV_X1    g0816(.A(G294), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n714), .A2(new_n789), .B1(new_n719), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n250), .B1(new_n702), .B2(new_n269), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n1016), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1014), .A2(new_n1015), .A3(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n710), .A2(new_n728), .B1(new_n361), .B2(new_n794), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT51), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n737), .A2(new_n202), .B1(new_n719), .B2(new_n388), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n250), .B1(new_n726), .B2(G87), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n410), .B2(new_n714), .C1(new_n784), .C2(new_n721), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT112), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1024), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1023), .B(new_n1028), .C1(new_n1027), .C2(new_n1026), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n702), .A2(new_n217), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1021), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n686), .B1(new_n1031), .B2(new_n691), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1012), .B(new_n1032), .C1(new_n934), .C2(new_n753), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1010), .A2(new_n1011), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1011), .B1(new_n1010), .B2(new_n1033), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1009), .B1(new_n1035), .B2(new_n1036), .ZN(G390));
  NAND4_X1  g0837(.A1(new_n678), .A2(G330), .A3(new_n680), .A4(new_n805), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n860), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n862), .A2(new_n847), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n846), .B2(new_n848), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n664), .A2(new_n650), .A3(new_n763), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n861), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n877), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n847), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1044), .A2(new_n1045), .A3(new_n863), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1039), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n848), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n844), .B1(new_n840), .B2(new_n842), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1049), .A2(new_n1050), .B1(new_n847), .B2(new_n862), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n681), .A2(new_n877), .A3(G330), .A4(new_n805), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1051), .A2(new_n1052), .A3(new_n1046), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1048), .A2(new_n1053), .A3(new_n945), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n748), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n365), .A2(new_n803), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n725), .A2(new_n410), .B1(new_n721), .B2(new_n1017), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n711), .B2(G116), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n211), .A2(new_n737), .B1(new_n794), .B2(new_n789), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n1059), .A2(new_n299), .A3(new_n734), .A4(new_n1030), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(new_n276), .C2(new_n719), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT114), .Z(new_n1062));
  OR3_X1    g0862(.A1(new_n714), .A2(KEYINPUT53), .A3(new_n361), .ZN(new_n1063));
  OAI21_X1  g0863(.A(KEYINPUT53), .B1(new_n714), .B2(new_n361), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n728), .C2(new_n702), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n250), .B1(new_n722), .B2(G125), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n693), .A2(G137), .B1(new_n698), .B2(G128), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(new_n202), .C2(new_n725), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1065), .B(new_n1068), .C1(G132), .C2(new_n711), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT54), .B(G143), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1069), .B1(new_n719), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1062), .A2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT115), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n686), .B1(new_n1073), .B2(new_n691), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1055), .A2(new_n1056), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n764), .A2(new_n861), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n860), .A2(new_n1038), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1076), .B1(new_n1077), .B2(new_n1039), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n771), .A2(new_n678), .A3(G330), .A4(new_n680), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n860), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1052), .A2(new_n861), .A3(new_n1080), .A4(new_n1042), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n489), .A2(G330), .A3(new_n681), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n871), .A2(new_n1082), .A3(new_n618), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(new_n1048), .A3(new_n1053), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n1004), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1085), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1054), .B(new_n1075), .C1(new_n1087), .C2(new_n1088), .ZN(G378));
  XNOR2_X1  g0889(.A(new_n376), .B(KEYINPUT55), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n368), .A2(new_n625), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT56), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1090), .B(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n748), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n803), .A2(new_n202), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n202), .B1(new_n247), .B2(G41), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n719), .A2(new_n387), .B1(new_n721), .B2(new_n789), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G58), .B2(new_n726), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n217), .B2(new_n714), .C1(new_n211), .C2(new_n710), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n735), .A2(G68), .B1(G116), .B2(new_n698), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT116), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n254), .B(new_n250), .C1(new_n737), .C2(new_n276), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1099), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT58), .Z(new_n1104));
  AOI22_X1  g0904(.A1(G137), .A2(new_n720), .B1(new_n735), .B2(G150), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n779), .B2(new_n737), .ZN(new_n1106));
  INV_X1    g0906(.A(G128), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n710), .A2(new_n1107), .B1(new_n714), .B2(new_n1070), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT117), .Z(new_n1109));
  AOI211_X1 g0909(.A(new_n1106), .B(new_n1109), .C1(G125), .C2(new_n698), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1112), .B(new_n253), .C1(new_n728), .C2(new_n725), .ZN(new_n1113));
  AOI21_X1  g0913(.A(G41), .B1(new_n722), .B2(G124), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1096), .B(new_n1104), .C1(new_n1113), .C2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n686), .B1(new_n1116), .B2(new_n691), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1094), .A2(new_n1095), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n880), .A2(G330), .A3(new_n881), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1093), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n880), .A2(new_n1093), .A3(G330), .A4(new_n881), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1124), .A2(new_n849), .A3(new_n864), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n865), .A2(new_n1123), .A3(new_n1122), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1119), .B1(new_n1127), .B2(new_n945), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT119), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n871), .A2(new_n618), .A3(new_n1083), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1086), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n1127), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT121), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT57), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1086), .A2(new_n1131), .B1(new_n1126), .B2(new_n1125), .ZN(new_n1137));
  OAI21_X1  g0937(.A(KEYINPUT121), .B1(new_n1137), .B2(KEYINPUT57), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT120), .ZN(new_n1140));
  OR2_X1    g0940(.A1(new_n1126), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1125), .A2(new_n1126), .A3(new_n1140), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1132), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1004), .B1(new_n1143), .B2(new_n1135), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1129), .B1(new_n1139), .B2(new_n1144), .ZN(G375));
  INV_X1    g0945(.A(new_n1082), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1130), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n968), .A3(new_n1084), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n860), .A2(new_n748), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n250), .B1(new_n725), .B2(new_n217), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT123), .Z(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G283), .B2(new_n711), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n983), .B1(G303), .B2(new_n722), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n1017), .B2(new_n794), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n737), .A2(new_n269), .B1(new_n719), .B2(new_n211), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(KEYINPUT122), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1155), .A2(KEYINPUT122), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1152), .B(new_n1158), .C1(new_n276), .C2(new_n714), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n721), .A2(new_n1107), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n714), .A2(new_n728), .B1(new_n719), .B2(new_n361), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n711), .B2(G137), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n702), .A2(new_n202), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n737), .A2(new_n1070), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(G132), .C2(new_n698), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n250), .B1(new_n726), .B2(G58), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1162), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1159), .B1(new_n1160), .B2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1168), .A2(new_n691), .B1(new_n410), .B2(new_n803), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1149), .A2(new_n755), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n1082), .B2(new_n945), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1148), .A2(new_n1171), .ZN(G381));
  OR2_X1    g0972(.A1(G375), .A2(G378), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(G384), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1175), .A2(new_n1171), .A3(new_n1148), .ZN(new_n1176));
  OR2_X1    g0976(.A1(G393), .A2(G396), .ZN(new_n1177));
  NOR4_X1   g0977(.A1(G387), .A2(G390), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1174), .A2(new_n1178), .ZN(G407));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n626), .ZN(new_n1180));
  OAI21_X1  g0980(.A(G213), .B1(new_n1173), .B2(new_n1180), .ZN(G409));
  NAND2_X1  g0981(.A1(G375), .A2(G378), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1132), .A2(new_n968), .A3(new_n1127), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1141), .A2(new_n945), .A3(new_n1142), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(new_n1184), .A3(new_n1118), .ZN(new_n1185));
  INV_X1    g0985(.A(G213), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n1185), .A2(G378), .B1(new_n1186), .B2(G343), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT60), .B1(new_n1130), .B2(new_n1146), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1130), .A2(KEYINPUT60), .A3(new_n1146), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1190), .A2(new_n1004), .A3(new_n1084), .A4(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n1171), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n1175), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(G384), .A3(new_n1171), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1182), .A2(new_n1188), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT63), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1200), .A2(KEYINPUT61), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n626), .A2(G213), .A3(G2897), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1196), .B(new_n1202), .Z(new_n1203));
  AOI21_X1  g1003(.A(new_n1187), .B1(G375), .B2(G378), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1198), .B1(new_n1205), .B2(new_n1199), .ZN(new_n1206));
  AND2_X1   g1006(.A1(G387), .A2(G390), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT124), .B1(G387), .B2(G390), .ZN(new_n1208));
  XOR2_X1   g1008(.A(G393), .B(G396), .Z(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  OR3_X1    g1010(.A1(new_n1207), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1210), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1201), .A2(new_n1206), .A3(new_n1213), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1205), .A2(KEYINPUT61), .ZN(new_n1215));
  AOI211_X1 g1015(.A(KEYINPUT125), .B(KEYINPUT62), .C1(new_n1204), .C2(new_n1197), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT125), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT62), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1217), .B1(new_n1198), .B2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1182), .A2(KEYINPUT62), .A3(new_n1188), .A4(new_n1197), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT126), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1204), .A2(KEYINPUT126), .A3(KEYINPUT62), .A4(new_n1197), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1215), .B1(new_n1220), .B2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1214), .B1(new_n1226), .B2(new_n1213), .ZN(G405));
  NAND2_X1  g1027(.A1(new_n1197), .A2(KEYINPUT127), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1213), .B(new_n1228), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1197), .A2(KEYINPUT127), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1173), .A2(new_n1182), .A3(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1229), .B(new_n1231), .ZN(G402));
endmodule


