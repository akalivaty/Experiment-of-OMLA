//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1217, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI21_X1  g0005(.A(G50), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  AND2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR3_X1   g0011(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n211), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n204), .A2(G50), .A3(new_n205), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n213), .A2(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G116), .ZN(new_n221));
  INV_X1    g0021(.A(G270), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G50), .ZN(new_n225));
  INV_X1    g0025(.A(G226), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n203), .C2(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n223), .B(new_n228), .C1(G97), .C2(G257), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(G1), .B2(G20), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT1), .Z(new_n231));
  AOI211_X1 g0031(.A(new_n219), .B(new_n231), .C1(new_n214), .C2(new_n213), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT65), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n249), .A2(new_n251), .A3(KEYINPUT65), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G238), .A2(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(G232), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n256), .B(new_n257), .C1(new_n258), .C2(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  OAI211_X1 g0060(.A(G1), .B(G13), .C1(new_n248), .C2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n259), .B(new_n262), .C1(G107), .C2(new_n256), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G244), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n261), .A2(new_n264), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n263), .B(new_n267), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n270), .A2(G179), .ZN(new_n271));
  XOR2_X1   g0071(.A(KEYINPUT8), .B(G58), .Z(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n272), .A2(new_n273), .B1(G20), .B2(G77), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT67), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n248), .A2(G20), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  XOR2_X1   g0077(.A(KEYINPUT15), .B(G87), .Z(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n275), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n215), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G1), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n280), .A2(new_n282), .B1(new_n207), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n282), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n210), .A2(G20), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G77), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n270), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n271), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT13), .ZN(new_n296));
  INV_X1    g0096(.A(G1698), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n226), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n258), .A2(G1698), .ZN(new_n299));
  AND3_X1   g0099(.A1(new_n249), .A2(new_n251), .A3(KEYINPUT65), .ZN(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT65), .B1(new_n249), .B2(new_n251), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n298), .B(new_n299), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G97), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n262), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n267), .B1(new_n269), .B2(new_n227), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n296), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n261), .B1(new_n302), .B2(new_n303), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n309), .A2(KEYINPUT13), .A3(new_n306), .ZN(new_n310));
  OAI21_X1  g0110(.A(G169), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT70), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT70), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n313), .B(G169), .C1(new_n308), .C2(new_n310), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n312), .A2(KEYINPUT14), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT71), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n311), .A2(KEYINPUT14), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n308), .A2(new_n310), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n318), .B1(G179), .B2(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n312), .A2(KEYINPUT71), .A3(KEYINPUT14), .A4(new_n314), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n317), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT72), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT72), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n317), .A2(new_n320), .A3(new_n324), .A4(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n273), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n277), .A2(new_n207), .B1(new_n225), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n211), .A2(G68), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n282), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT11), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n288), .A2(G68), .A3(new_n289), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n330), .B2(new_n331), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n329), .A2(new_n284), .ZN(new_n335));
  XOR2_X1   g0135(.A(new_n335), .B(KEYINPUT12), .Z(new_n336));
  NOR3_X1   g0136(.A1(new_n332), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n295), .B1(new_n326), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT17), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n272), .A2(new_n289), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT75), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n286), .A2(new_n282), .ZN(new_n343));
  INV_X1    g0143(.A(new_n272), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n342), .A2(new_n343), .B1(new_n344), .B2(new_n286), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n249), .A2(new_n251), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n226), .A2(G1698), .ZN(new_n347));
  OR2_X1    g0147(.A1(G223), .A2(G1698), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G87), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n248), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n262), .ZN(new_n352));
  INV_X1    g0152(.A(new_n269), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G232), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n267), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G200), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n300), .A2(new_n301), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT7), .B1(new_n357), .B2(new_n211), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT74), .B1(new_n250), .B2(G33), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT74), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(new_n248), .A3(KEYINPUT3), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n361), .A3(new_n251), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n362), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n363));
  OAI21_X1  g0163(.A(G68), .B1(new_n358), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G159), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n365), .A2(G20), .A3(G33), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G58), .A2(G68), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n204), .A2(new_n205), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n366), .B1(new_n368), .B2(G20), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT16), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT7), .B1(new_n346), .B2(G20), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT7), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n252), .A2(new_n372), .A3(new_n211), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(G68), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT73), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  AOI211_X1 g0176(.A(KEYINPUT73), .B(new_n366), .C1(new_n368), .C2(G20), .ZN(new_n377));
  OAI211_X1 g0177(.A(KEYINPUT16), .B(new_n374), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n282), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n345), .B(new_n356), .C1(new_n370), .C2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G190), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n355), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n340), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n345), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n378), .A2(new_n282), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT16), .ZN(new_n386));
  INV_X1    g0186(.A(new_n363), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n254), .A2(new_n211), .A3(new_n255), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n372), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n203), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n369), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n386), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n384), .B1(new_n385), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n382), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n393), .A2(KEYINPUT17), .A3(new_n394), .A4(new_n356), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n383), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n345), .B1(new_n370), .B2(new_n379), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n355), .A2(G169), .ZN(new_n398));
  INV_X1    g0198(.A(G179), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(new_n355), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT18), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n397), .A2(KEYINPUT18), .A3(new_n400), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n396), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n291), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n270), .A2(G200), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n406), .B(new_n407), .C1(new_n381), .C2(new_n270), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G223), .A2(G1698), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n297), .A2(G222), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n256), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n357), .A2(new_n207), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n262), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n353), .A2(G226), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n267), .A3(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n415), .A2(new_n292), .ZN(new_n416));
  OR2_X1    g0216(.A1(KEYINPUT8), .A2(G58), .ZN(new_n417));
  NAND2_X1  g0217(.A1(KEYINPUT8), .A2(G58), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n276), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n206), .B2(new_n211), .ZN(new_n420));
  INV_X1    g0220(.A(G150), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n327), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n282), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n289), .A2(G50), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT66), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n343), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n286), .A2(new_n225), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n415), .B2(G179), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n416), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(KEYINPUT9), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT9), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n423), .A2(new_n426), .A3(new_n432), .A4(new_n427), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n431), .A2(KEYINPUT68), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT68), .B1(new_n431), .B2(new_n433), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n415), .A2(KEYINPUT69), .A3(G200), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT69), .B1(new_n415), .B2(G200), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT10), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n415), .A2(new_n381), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n436), .A2(new_n440), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n439), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n437), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n431), .A2(new_n433), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT10), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n430), .B1(new_n443), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n338), .B1(new_n319), .B2(G190), .ZN(new_n450));
  INV_X1    g0250(.A(G200), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(new_n319), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n405), .A2(new_n408), .A3(new_n449), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT76), .B1(new_n339), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n337), .B1(new_n323), .B2(new_n325), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT76), .ZN(new_n457));
  NOR4_X1   g0257(.A1(new_n456), .A2(new_n453), .A3(new_n457), .A4(new_n295), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n288), .B1(G20), .B2(new_n221), .ZN(new_n460));
  AOI21_X1  g0260(.A(G20), .B1(G33), .B2(G283), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT77), .B(G97), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(G33), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n460), .A2(KEYINPUT20), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n460), .A2(new_n463), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT20), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n210), .A2(G33), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n288), .A2(new_n285), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n464), .A2(new_n467), .B1(G116), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n285), .A2(G116), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  OR2_X1    g0274(.A1(new_n297), .A2(G264), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n346), .B(new_n475), .C1(G257), .C2(G1698), .ZN(new_n476));
  INV_X1    g0276(.A(G303), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n476), .B1(new_n256), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n262), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT80), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G45), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G1), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT5), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G41), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n261), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(new_n222), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n487), .A2(new_n265), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT79), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n490), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT79), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n492), .B(new_n493), .C1(new_n222), .C2(new_n488), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n478), .A2(KEYINPUT80), .A3(new_n262), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n481), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n474), .A2(new_n497), .A3(G169), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT21), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(G200), .ZN(new_n501));
  INV_X1    g0301(.A(new_n474), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n481), .A2(new_n495), .A3(G190), .A4(new_n496), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n497), .A2(new_n399), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n474), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n474), .A2(new_n497), .A3(KEYINPUT21), .A4(G169), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n500), .A2(new_n504), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n227), .A2(new_n297), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n268), .A2(G1698), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n249), .A2(new_n509), .A3(new_n251), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G116), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n261), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n210), .A2(G45), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n261), .A2(G250), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n483), .A2(G274), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n513), .A2(new_n517), .A3(G179), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n278), .A2(new_n285), .ZN(new_n519));
  INV_X1    g0319(.A(G107), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n462), .A2(new_n350), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT19), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n211), .B1(new_n303), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n346), .A2(new_n211), .A3(G68), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n522), .B1(new_n462), .B2(new_n277), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n519), .B1(new_n527), .B2(new_n282), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n470), .A2(new_n278), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n518), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n513), .A2(new_n517), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n292), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n513), .A2(new_n517), .A3(new_n381), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n532), .B2(G200), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n469), .A2(new_n350), .ZN(new_n537));
  AOI211_X1 g0337(.A(new_n519), .B(new_n537), .C1(new_n527), .C2(new_n282), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n508), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT24), .ZN(new_n542));
  NOR2_X1   g0342(.A1(KEYINPUT22), .A2(G20), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n256), .A2(G87), .A3(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n249), .A2(new_n251), .A3(new_n211), .A4(G87), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT22), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n546), .A2(KEYINPUT81), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT81), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n545), .B2(KEYINPUT22), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n544), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT82), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n544), .B(KEYINPUT82), .C1(new_n547), .C2(new_n549), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n211), .A2(G107), .ZN(new_n555));
  NOR2_X1   g0355(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n556));
  OR2_X1    g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n276), .A2(G116), .ZN(new_n558));
  AND2_X1   g0358(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n555), .B1(new_n559), .B2(new_n556), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n542), .B1(new_n554), .B2(new_n562), .ZN(new_n563));
  AOI211_X1 g0363(.A(KEYINPUT24), .B(new_n561), .C1(new_n552), .C2(new_n553), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n282), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n284), .A2(new_n555), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n566), .B(KEYINPUT25), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(G107), .B2(new_n470), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT84), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n346), .A2(new_n569), .A3(G250), .A4(new_n297), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n346), .A2(G257), .A3(G1698), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G294), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n249), .A2(new_n251), .A3(G250), .A4(new_n297), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT84), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n570), .A2(new_n571), .A3(new_n572), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n262), .ZN(new_n576));
  INV_X1    g0376(.A(new_n488), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G264), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n578), .A3(new_n492), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n451), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G190), .B2(new_n579), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n565), .A2(new_n568), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(G169), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT85), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n576), .A2(G179), .A3(new_n578), .A4(new_n492), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n584), .B1(new_n583), .B2(new_n585), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n553), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n546), .B(KEYINPUT81), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT82), .B1(new_n591), .B2(new_n544), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n562), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT24), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n554), .A2(new_n542), .A3(new_n562), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n288), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n568), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n589), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n273), .A2(G77), .ZN(new_n599));
  INV_X1    g0399(.A(new_n462), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n600), .A2(KEYINPUT6), .A3(new_n520), .ZN(new_n601));
  XOR2_X1   g0401(.A(G97), .B(G107), .Z(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(KEYINPUT6), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G20), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n363), .B1(new_n372), .B2(new_n388), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n599), .B(new_n604), .C1(new_n605), .C2(new_n520), .ZN(new_n606));
  INV_X1    g0406(.A(G97), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n606), .A2(new_n282), .B1(new_n607), .B2(new_n286), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n470), .A2(G97), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n577), .A2(G257), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n346), .A2(G244), .A3(new_n297), .ZN(new_n611));
  XOR2_X1   g0411(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n612));
  AOI22_X1  g0412(.A1(new_n611), .A2(new_n612), .B1(G33), .B2(G283), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n297), .A2(KEYINPUT4), .A3(G244), .ZN(new_n614));
  INV_X1    g0414(.A(G250), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(new_n297), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n256), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n610), .B1(new_n618), .B2(new_n262), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n492), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n608), .A2(new_n609), .B1(new_n292), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n399), .A3(new_n492), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n606), .A2(new_n282), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n286), .A2(new_n607), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n624), .A3(new_n609), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n261), .B1(new_n613), .B2(new_n617), .ZN(new_n627));
  NOR4_X1   g0427(.A1(new_n627), .A2(new_n381), .A3(new_n490), .A4(new_n610), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(G200), .B2(new_n620), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n621), .A2(new_n622), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n541), .A2(new_n582), .A3(new_n598), .A4(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n459), .A2(new_n631), .ZN(G372));
  NAND2_X1  g0432(.A1(new_n403), .A2(new_n404), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n383), .A2(new_n395), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n452), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n633), .B1(new_n339), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n443), .A2(new_n448), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n430), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n620), .A2(new_n292), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n625), .A2(new_n639), .A3(new_n622), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT26), .B1(new_n640), .B2(new_n540), .ZN(new_n641));
  INV_X1    g0441(.A(new_n513), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT86), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n515), .A2(new_n643), .A3(new_n516), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n515), .B2(new_n516), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n292), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n530), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT87), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n530), .A2(KEYINPUT87), .A3(new_n647), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n535), .B1(new_n646), .B2(G200), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n530), .A2(new_n647), .B1(new_n653), .B2(new_n538), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n625), .A2(new_n654), .A3(new_n639), .A4(new_n622), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n641), .B(new_n652), .C1(KEYINPUT26), .C2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n626), .A2(new_n629), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n640), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n583), .A2(new_n585), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n596), .B2(new_n597), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n500), .A2(new_n506), .A3(new_n507), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n658), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n582), .A2(new_n654), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n656), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n638), .B1(new_n459), .B2(new_n665), .ZN(G369));
  NOR2_X1   g0466(.A1(new_n283), .A2(G20), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n210), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n596), .B2(new_n597), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n598), .A2(new_n674), .A3(new_n582), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT88), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n673), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n598), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G330), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n502), .A2(new_n680), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n508), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n661), .A2(new_n683), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n565), .A2(new_n568), .B1(new_n583), .B2(new_n585), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n680), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n662), .A2(new_n673), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n677), .A2(new_n678), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n687), .A2(new_n689), .A3(new_n691), .ZN(G399));
  OR2_X1    g0492(.A1(new_n521), .A2(G116), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n693), .B(KEYINPUT89), .Z(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n212), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n218), .B2(new_n698), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT28), .Z(new_n701));
  INV_X1    g0501(.A(KEYINPUT90), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n665), .B2(new_n673), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n630), .B1(new_n688), .B2(new_n661), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n582), .A2(new_n654), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g0506(.A(KEYINPUT90), .B(new_n680), .C1(new_n706), .C2(new_n656), .ZN(new_n707));
  XOR2_X1   g0507(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n708));
  NAND3_X1  g0508(.A1(new_n703), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT92), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT26), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n534), .A2(new_n539), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n621), .A2(new_n711), .A3(new_n712), .A4(new_n622), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n655), .A2(KEYINPUT26), .ZN(new_n714));
  AND4_X1   g0514(.A1(new_n710), .A2(new_n713), .A3(new_n714), .A4(new_n652), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n655), .A2(KEYINPUT26), .B1(new_n651), .B2(new_n650), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n710), .B1(new_n716), .B2(new_n713), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n598), .A2(new_n662), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n630), .A2(KEYINPUT93), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n657), .A2(new_n640), .A3(KEYINPUT93), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n664), .B(new_n719), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n673), .B1(new_n718), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT29), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n709), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n579), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n505), .A2(new_n726), .A3(new_n619), .A4(new_n531), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n646), .A2(new_n399), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n620), .A2(new_n497), .A3(new_n579), .A4(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n727), .A2(new_n728), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n673), .ZN(new_n734));
  OAI211_X1 g0534(.A(KEYINPUT31), .B(new_n734), .C1(new_n631), .C2(new_n673), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n734), .A2(KEYINPUT31), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n725), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n701), .B1(new_n739), .B2(new_n210), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT94), .ZN(G364));
  XNOR2_X1  g0541(.A(new_n667), .B(KEYINPUT96), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n210), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n697), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n215), .B1(G20), .B2(new_n292), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n211), .A2(new_n381), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n399), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G322), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n211), .A2(G190), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G179), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G329), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n750), .A2(new_n751), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G283), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n451), .A2(G179), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n752), .ZN(new_n759));
  INV_X1    g0559(.A(G294), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n753), .A2(G190), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n357), .B1(new_n757), .B2(new_n759), .C1(new_n760), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n752), .A2(new_n749), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n756), .B(new_n764), .C1(G311), .C2(new_n766), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n211), .A2(new_n399), .A3(new_n451), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT97), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n381), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G326), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n748), .A2(new_n758), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G303), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n769), .A2(G190), .ZN(new_n775));
  XNOR2_X1  g0575(.A(KEYINPUT33), .B(G317), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n767), .A2(new_n771), .A3(new_n774), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT32), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n754), .A2(new_n365), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n779), .A2(new_n780), .B1(new_n763), .B2(new_n607), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n357), .B(new_n781), .C1(new_n779), .C2(new_n780), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G50), .A2(new_n770), .B1(new_n775), .B2(G68), .ZN(new_n783));
  INV_X1    g0583(.A(new_n759), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G107), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n202), .A2(new_n750), .B1(new_n772), .B2(new_n350), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(G77), .B2(new_n766), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n782), .A2(new_n783), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n747), .B1(new_n778), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n746), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n243), .A2(G45), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n696), .A2(new_n346), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n794), .B(new_n795), .C1(G45), .C2(new_n218), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n256), .A2(G355), .A3(new_n212), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n796), .B(new_n797), .C1(G116), .C2(new_n212), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n789), .B1(new_n793), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n684), .A2(new_n685), .ZN(new_n800));
  INV_X1    g0600(.A(new_n792), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n745), .B(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n686), .B(KEYINPUT95), .ZN(new_n803));
  INV_X1    g0603(.A(new_n745), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n800), .B2(G330), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n802), .B1(new_n803), .B2(new_n805), .ZN(G396));
  NOR2_X1   g0606(.A1(new_n665), .A2(new_n673), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n295), .A2(new_n680), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n408), .B1(new_n406), .B2(new_n680), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(new_n294), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n703), .A2(new_n707), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n813), .B2(new_n811), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(new_n738), .Z(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n804), .ZN(new_n816));
  INV_X1    g0616(.A(new_n750), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n775), .A2(G150), .B1(G143), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n770), .A2(G137), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(new_n365), .C2(new_n765), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT34), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n346), .B1(new_n754), .B2(new_n822), .C1(new_n225), .C2(new_n772), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G58), .B2(new_n762), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n821), .B(new_n824), .C1(new_n203), .C2(new_n759), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G283), .A2(new_n775), .B1(new_n770), .B2(G303), .ZN(new_n826));
  INV_X1    g0626(.A(G311), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n772), .A2(new_n520), .B1(new_n754), .B2(new_n827), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n763), .A2(new_n607), .B1(new_n750), .B2(new_n760), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(G116), .C2(new_n766), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n784), .A2(G87), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n826), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n825), .B1(new_n256), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n804), .B1(new_n833), .B2(new_n746), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n746), .A2(new_n790), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(G77), .B2(new_n836), .C1(new_n811), .C2(new_n791), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n816), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G384));
  NOR2_X1   g0639(.A1(new_n337), .A2(new_n680), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n452), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT98), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n326), .B2(new_n338), .ZN(new_n845));
  AOI211_X1 g0645(.A(KEYINPUT98), .B(new_n337), .C1(new_n323), .C2(new_n325), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n323), .A2(new_n325), .A3(new_n452), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n840), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n850), .A2(new_n737), .A3(new_n811), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n369), .B(new_n375), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT16), .B1(new_n852), .B2(new_n374), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n345), .B1(new_n853), .B2(new_n379), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT99), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT99), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n856), .B(new_n345), .C1(new_n853), .C2(new_n379), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n855), .A2(new_n400), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n671), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n855), .A2(new_n859), .A3(new_n857), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n393), .A2(new_n394), .A3(new_n356), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n397), .B1(new_n400), .B2(new_n859), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n861), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n634), .A2(new_n633), .ZN(new_n869));
  INV_X1    g0669(.A(new_n860), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n868), .A2(new_n871), .A3(KEYINPUT38), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n866), .B1(new_n862), .B2(KEYINPUT37), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n860), .B1(new_n634), .B2(new_n633), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n851), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT40), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n405), .A2(new_n393), .A3(new_n671), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n865), .B1(new_n861), .B2(new_n864), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n866), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n873), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n872), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n851), .A2(KEYINPUT40), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n459), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n888), .A2(new_n737), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n887), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(G330), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n809), .B1(new_n807), .B2(new_n811), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n849), .B2(new_n847), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n877), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n868), .B2(new_n871), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n874), .A2(new_n875), .A3(new_n873), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT39), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT100), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n884), .A2(new_n899), .A3(new_n872), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT100), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n877), .A2(new_n901), .A3(KEYINPUT39), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n898), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n326), .A2(new_n338), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT98), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n456), .A2(new_n844), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n680), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n894), .B(new_n909), .C1(new_n633), .C2(new_n859), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n709), .B(new_n724), .C1(new_n455), .C2(new_n458), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n638), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n910), .B(new_n912), .Z(new_n913));
  XNOR2_X1  g0713(.A(new_n891), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n210), .B2(new_n742), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n221), .B1(new_n603), .B2(KEYINPUT35), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n916), .B(new_n216), .C1(KEYINPUT35), .C2(new_n603), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT36), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n367), .A2(G77), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n218), .A2(new_n919), .B1(G50), .B2(new_n203), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(G1), .A3(new_n283), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n915), .A2(new_n918), .A3(new_n921), .ZN(G367));
  OAI22_X1  g0722(.A1(new_n720), .A2(new_n721), .B1(new_n626), .B2(new_n680), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n621), .A2(new_n622), .A3(new_n673), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT101), .Z(new_n926));
  INV_X1    g0726(.A(new_n598), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n640), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT102), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n928), .A2(KEYINPUT102), .A3(new_n640), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(new_n680), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n538), .A2(new_n680), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n654), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n652), .B2(new_n935), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n691), .A2(new_n923), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT42), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n933), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT103), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n938), .B1(new_n933), .B2(new_n940), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n926), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n946), .B1(new_n687), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n691), .A2(new_n689), .ZN(new_n949));
  INV_X1    g0749(.A(new_n925), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT45), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(new_n950), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT44), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(new_n687), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n681), .A2(new_n690), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n803), .B1(new_n959), .B2(new_n691), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n959), .A2(new_n691), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n960), .B1(new_n686), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n739), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n697), .B(KEYINPUT41), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n743), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n947), .A2(new_n687), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n942), .A2(new_n967), .A3(new_n945), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n948), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n795), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n793), .B1(new_n212), .B2(new_n279), .C1(new_n239), .C2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n745), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT104), .Z(new_n973));
  AOI21_X1  g0773(.A(new_n357), .B1(G58), .B2(new_n773), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n759), .A2(new_n207), .ZN(new_n975));
  INV_X1    g0775(.A(new_n754), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n975), .B1(G137), .B2(new_n976), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n766), .A2(G50), .B1(new_n762), .B2(G68), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n974), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(G143), .ZN(new_n980));
  INV_X1    g0780(.A(new_n770), .ZN(new_n981));
  INV_X1    g0781(.A(new_n775), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n980), .A2(new_n981), .B1(new_n982), .B2(new_n365), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n979), .B(new_n983), .C1(G150), .C2(new_n817), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n976), .A2(G317), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n760), .A2(new_n982), .B1(new_n981), .B2(new_n827), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n600), .A2(new_n784), .B1(new_n766), .B2(G283), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n477), .B2(new_n750), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n773), .A2(KEYINPUT46), .A3(G116), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n346), .B1(G107), .B2(new_n762), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT46), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n772), .B2(new_n221), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n986), .A2(new_n988), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n984), .B1(new_n985), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT47), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n973), .B1(new_n801), .B2(new_n937), .C1(new_n996), .C2(new_n747), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n969), .A2(new_n997), .ZN(G387));
  AND2_X1   g0798(.A1(new_n976), .A2(G326), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G311), .A2(new_n775), .B1(new_n770), .B2(G322), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT105), .Z(new_n1001));
  NAND2_X1  g0801(.A1(new_n817), .A2(G317), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(new_n477), .C2(new_n765), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT48), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n757), .B2(new_n763), .C1(new_n760), .C2(new_n772), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT49), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n346), .B(new_n999), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n1006), .B2(new_n1005), .C1(new_n221), .C2(new_n759), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n346), .B1(new_n759), .B2(new_n607), .C1(new_n981), .C2(new_n365), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n772), .A2(new_n207), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n765), .A2(new_n203), .B1(new_n754), .B2(new_n421), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1010), .B(new_n1011), .C1(G50), .C2(new_n817), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n279), .B2(new_n763), .C1(new_n982), .C2(new_n344), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1008), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n804), .B1(new_n1014), .B2(new_n746), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n694), .A2(new_n212), .A3(new_n256), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n795), .B1(new_n236), .B2(new_n482), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n344), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1018));
  OAI21_X1  g0818(.A(KEYINPUT50), .B1(new_n344), .B2(G50), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n482), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1018), .B(new_n1020), .C1(G68), .C2(G77), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1016), .A2(new_n1017), .B1(new_n695), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n212), .A2(G107), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n793), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1015), .B(new_n1024), .C1(new_n681), .C2(new_n801), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n962), .A2(new_n744), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n739), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n962), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n697), .B1(new_n962), .B2(new_n1027), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1025), .B(new_n1026), .C1(new_n1028), .C2(new_n1029), .ZN(G393));
  OR2_X1    g0830(.A1(new_n957), .A2(new_n1028), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n957), .A2(new_n1028), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1031), .A2(new_n697), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT106), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1031), .A2(KEYINPUT106), .A3(new_n697), .A4(new_n1032), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n957), .A2(new_n744), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n793), .B1(new_n212), .B2(new_n462), .C1(new_n246), .C2(new_n970), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n770), .A2(G317), .B1(G311), .B2(new_n817), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT52), .Z(new_n1041));
  OAI21_X1  g0841(.A(new_n357), .B1(new_n221), .B2(new_n763), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n785), .B1(new_n760), .B2(new_n765), .C1(new_n751), .C2(new_n754), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(G303), .C2(new_n775), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1041), .B(new_n1044), .C1(new_n757), .C2(new_n772), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n344), .A2(new_n765), .B1(new_n980), .B2(new_n754), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1047), .B(new_n831), .C1(new_n203), .C2(new_n772), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n982), .A2(new_n225), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n981), .A2(new_n421), .B1(new_n365), .B2(new_n750), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT51), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1048), .B(new_n1049), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n1051), .B2(new_n1050), .C1(new_n207), .C2(new_n763), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1045), .B1(new_n1053), .B2(new_n252), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n804), .B1(new_n1054), .B2(new_n746), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1039), .B(new_n1055), .C1(new_n926), .C2(new_n801), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1037), .A2(new_n1038), .A3(new_n1056), .ZN(G390));
  NAND4_X1  g0857(.A1(new_n735), .A2(new_n736), .A3(G330), .A4(new_n811), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n847), .B2(new_n849), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n812), .A2(new_n808), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n842), .B1(new_n905), .B2(new_n906), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n849), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n903), .B1(new_n1063), .B2(new_n907), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n907), .A2(new_n885), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n810), .A2(new_n294), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n809), .B1(new_n723), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1065), .B1(new_n850), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1059), .B1(new_n1064), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n899), .B1(new_n872), .B2(new_n876), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT100), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n900), .B(new_n1072), .C1(new_n893), .C2(new_n908), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n850), .A2(new_n1068), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1074), .A2(new_n907), .A3(new_n885), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1058), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1073), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1070), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n744), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n772), .A2(new_n421), .ZN(new_n1082));
  XOR2_X1   g0882(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n1083));
  XNOR2_X1  g0883(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n357), .B(new_n1084), .C1(G159), .C2(new_n762), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n976), .A2(G125), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G128), .A2(new_n770), .B1(new_n775), .B2(G137), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n750), .A2(new_n822), .B1(new_n759), .B2(new_n225), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(KEYINPUT54), .B(G143), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT111), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1088), .B1(new_n1090), .B2(new_n766), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .A4(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n750), .A2(new_n221), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G107), .A2(new_n775), .B1(new_n770), .B2(G283), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n759), .A2(new_n203), .B1(new_n754), .B2(new_n760), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT113), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n772), .A2(new_n350), .B1(new_n765), .B2(new_n462), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n256), .B(new_n1097), .C1(G77), .C2(new_n762), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1092), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n804), .B1(new_n1100), .B2(new_n746), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1101), .B1(new_n272), .B2(new_n836), .C1(new_n903), .C2(new_n791), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT108), .ZN(new_n1103));
  OAI211_X1 g0903(.A(G330), .B(new_n737), .C1(new_n455), .C2(new_n458), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n911), .A2(new_n1104), .A3(new_n638), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(KEYINPUT107), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT107), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n911), .A2(new_n1104), .A3(new_n1107), .A4(new_n638), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n847), .A2(new_n849), .A3(new_n1058), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n1110), .A2(new_n1059), .A3(new_n1068), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n847), .A2(new_n849), .A3(new_n1058), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n892), .B1(new_n1077), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1103), .B1(new_n1109), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1060), .B1(new_n1110), .B2(new_n1059), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1077), .A2(new_n1067), .A3(new_n1112), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1118), .A2(new_n1106), .A3(KEYINPUT108), .A4(new_n1108), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1115), .A2(new_n1079), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT110), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT109), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n1080), .ZN(new_n1124));
  AOI211_X1 g0924(.A(KEYINPUT109), .B(new_n1079), .C1(new_n1115), .C2(new_n1119), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1121), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n697), .B1(new_n1120), .B2(KEYINPUT110), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1081), .B(new_n1102), .C1(new_n1126), .C2(new_n1127), .ZN(G378));
  INV_X1    g0928(.A(new_n1109), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT55), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n449), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n449), .A2(new_n1131), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n428), .A2(new_n859), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1139), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n887), .B2(new_n682), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1143), .B(KEYINPUT117), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1146), .A2(new_n880), .A3(G330), .A4(new_n886), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1145), .A2(new_n1147), .A3(new_n910), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n910), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1130), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT57), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1130), .A2(KEYINPUT57), .A3(new_n1150), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n697), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n770), .A2(G125), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n775), .A2(G132), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1090), .A2(new_n773), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n817), .A2(G128), .B1(new_n762), .B2(G150), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G137), .B2(new_n766), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT59), .ZN(new_n1162));
  AOI21_X1  g0962(.A(G41), .B1(new_n976), .B2(G124), .ZN(new_n1163));
  AOI21_X1  g0963(.A(G33), .B1(new_n784), .B2(G159), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n770), .A2(G116), .B1(G68), .B2(new_n762), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT115), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n775), .A2(G97), .B1(new_n278), .B2(new_n766), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT114), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n784), .A2(G58), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n750), .A2(new_n520), .B1(new_n754), .B2(new_n757), .ZN(new_n1171));
  NOR4_X1   g0971(.A1(new_n1171), .A2(new_n1010), .A3(G41), .A4(new_n346), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1167), .A2(new_n1169), .A3(new_n1170), .A4(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT58), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n260), .B1(new_n250), .B2(new_n248), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1173), .A2(new_n1174), .B1(new_n225), .B2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1165), .B(new_n1176), .C1(new_n1174), .C2(new_n1173), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n804), .B1(new_n1177), .B2(new_n746), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(G50), .B2(new_n836), .C1(new_n1146), .C2(new_n791), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT118), .Z(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n744), .B2(new_n1150), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1155), .A2(new_n1181), .ZN(G375));
  NAND2_X1  g0982(.A1(new_n835), .A2(new_n203), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n850), .A2(new_n791), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1170), .A2(new_n346), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT120), .ZN(new_n1186));
  INV_X1    g0986(.A(G128), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n765), .A2(new_n421), .B1(new_n754), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G50), .B2(new_n762), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1186), .B(new_n1189), .C1(new_n365), .C2(new_n772), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1190), .A2(KEYINPUT121), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n817), .A2(G137), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1190), .A2(KEYINPUT121), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G132), .A2(new_n770), .B1(new_n775), .B2(new_n1090), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n357), .B1(new_n757), .B2(new_n750), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n772), .A2(new_n607), .B1(new_n765), .B2(new_n520), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G303), .B2(new_n976), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n279), .B2(new_n763), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1196), .B(new_n1199), .C1(G77), .C2(new_n784), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n221), .B2(new_n982), .C1(new_n760), .C2(new_n981), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n747), .B1(new_n1195), .B2(new_n1201), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n1184), .A2(new_n804), .A3(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1118), .A2(new_n744), .B1(new_n1183), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1109), .A2(new_n1114), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT119), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1206), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1204), .B1(new_n1207), .B2(new_n965), .ZN(G381));
  INV_X1    g1008(.A(G387), .ZN(new_n1209));
  INV_X1    g1009(.A(G390), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(G378), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1155), .A2(new_n1212), .A3(new_n1181), .ZN(new_n1213));
  OR2_X1    g1013(.A1(G393), .A2(G396), .ZN(new_n1214));
  OR2_X1    g1014(.A1(G381), .A2(G384), .ZN(new_n1215));
  OR4_X1    g1015(.A1(new_n1211), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(G407));
  NAND2_X1  g1016(.A1(new_n672), .A2(G213), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT122), .Z(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(G407), .B(G213), .C1(new_n1213), .C2(new_n1219), .ZN(G409));
  INV_X1    g1020(.A(KEYINPUT126), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1211), .A2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1223));
  XOR2_X1   g1023(.A(G393), .B(G396), .Z(new_n1224));
  OR3_X1    g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1224), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT62), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1154), .A2(new_n697), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT57), .B1(new_n1130), .B2(new_n1150), .ZN(new_n1230));
  OAI211_X1 g1030(.A(G378), .B(new_n1181), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT123), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT123), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1155), .A2(new_n1233), .A3(G378), .A4(new_n1181), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1130), .A2(new_n964), .A3(new_n1150), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G378), .B1(new_n1181), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1235), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT127), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1240), .A3(new_n1219), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1237), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1242));
  OAI21_X1  g1042(.A(KEYINPUT127), .B1(new_n1242), .B2(new_n1218), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT60), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1206), .B1(new_n1245), .B2(new_n1123), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT124), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n698), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1109), .A2(KEYINPUT60), .A3(new_n1114), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(new_n1247), .C2(new_n1246), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1204), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n838), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(G384), .A3(new_n1204), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1228), .B1(new_n1244), .B2(new_n1255), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1242), .A2(new_n1218), .A3(new_n1254), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT61), .B1(new_n1257), .B2(new_n1228), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1218), .A2(G2897), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n1259), .B(KEYINPUT125), .Z(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1254), .A2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1252), .A2(new_n1253), .A3(new_n1260), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1241), .A2(new_n1243), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1258), .A2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1227), .B1(new_n1256), .B2(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1242), .A2(new_n1218), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT63), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1257), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1227), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1244), .A2(KEYINPUT63), .A3(new_n1255), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1272), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1267), .A2(new_n1275), .ZN(G405));
  NAND2_X1  g1076(.A1(G375), .A2(new_n1212), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1235), .A2(new_n1277), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1225), .A2(new_n1226), .A3(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1278), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1280));
  OR3_X1    g1080(.A1(new_n1279), .A2(new_n1280), .A3(new_n1254), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1254), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(G402));
endmodule


