

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(n738), .A2(n737), .ZN(n740) );
  OR2_X1 U556 ( .A1(n701), .A2(n787), .ZN(n745) );
  NOR2_X1 U557 ( .A1(n652), .A2(n545), .ZN(n636) );
  NOR2_X1 U558 ( .A1(G543), .A2(G651), .ZN(n640) );
  XOR2_X1 U559 ( .A(KEYINPUT7), .B(n600), .Z(G168) );
  NAND2_X1 U560 ( .A1(n745), .A2(G8), .ZN(n782) );
  XOR2_X1 U561 ( .A(KEYINPUT0), .B(G543), .Z(n652) );
  NAND2_X1 U562 ( .A1(n754), .A2(n753), .ZN(n776) );
  NOR2_X1 U563 ( .A1(n705), .A2(n704), .ZN(n707) );
  NOR2_X2 U564 ( .A1(n701), .A2(n787), .ZN(n719) );
  AND2_X2 U565 ( .A1(n526), .A2(G2104), .ZN(n891) );
  INV_X1 U566 ( .A(n1002), .ZN(n771) );
  OR2_X1 U567 ( .A1(G1966), .A2(n782), .ZN(n698) );
  INV_X1 U568 ( .A(KEYINPUT31), .ZN(n706) );
  INV_X1 U569 ( .A(KEYINPUT100), .ZN(n760) );
  XNOR2_X1 U570 ( .A(n527), .B(KEYINPUT65), .ZN(n528) );
  AND2_X1 U571 ( .A1(n785), .A2(n784), .ZN(n786) );
  AND2_X1 U572 ( .A1(n783), .A2(n524), .ZN(n784) );
  NAND2_X1 U573 ( .A1(n890), .A2(G137), .ZN(n693) );
  OR2_X1 U574 ( .A1(G301), .A2(n732), .ZN(n521) );
  AND2_X1 U575 ( .A1(n763), .A2(n762), .ZN(n522) );
  NAND2_X1 U576 ( .A1(G8), .A2(n741), .ZN(n523) );
  OR2_X1 U577 ( .A1(n782), .A2(n781), .ZN(n524) );
  NOR2_X1 U578 ( .A1(n772), .A2(n771), .ZN(n525) );
  NOR2_X1 U579 ( .A1(n722), .A2(n721), .ZN(n725) );
  INV_X1 U580 ( .A(KEYINPUT29), .ZN(n730) );
  XNOR2_X1 U581 ( .A(n731), .B(n730), .ZN(n733) );
  INV_X1 U582 ( .A(n996), .ZN(n756) );
  AND2_X1 U583 ( .A1(n757), .A2(n756), .ZN(n758) );
  INV_X1 U584 ( .A(KEYINPUT97), .ZN(n739) );
  OR2_X1 U585 ( .A1(G1384), .A2(n688), .ZN(n689) );
  NAND2_X1 U586 ( .A1(n695), .A2(n694), .ZN(n787) );
  INV_X1 U587 ( .A(G2105), .ZN(n526) );
  XNOR2_X1 U588 ( .A(KEYINPUT5), .B(KEYINPUT75), .ZN(n596) );
  INV_X1 U589 ( .A(KEYINPUT17), .ZN(n532) );
  AND2_X1 U590 ( .A1(n534), .A2(G2105), .ZN(n887) );
  XNOR2_X1 U591 ( .A(n580), .B(KEYINPUT15), .ZN(n985) );
  XNOR2_X1 U592 ( .A(n597), .B(n596), .ZN(n598) );
  NAND2_X1 U593 ( .A1(G101), .A2(n891), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(KEYINPUT23), .ZN(n531) );
  AND2_X1 U595 ( .A1(G2104), .A2(G2105), .ZN(n886) );
  NAND2_X1 U596 ( .A1(G113), .A2(n886), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n529), .B(KEYINPUT66), .ZN(n530) );
  AND2_X1 U598 ( .A1(n531), .A2(n530), .ZN(n695) );
  NOR2_X1 U599 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  XNOR2_X2 U600 ( .A(n533), .B(n532), .ZN(n890) );
  INV_X1 U601 ( .A(G2104), .ZN(n534) );
  NAND2_X1 U602 ( .A1(G125), .A2(n887), .ZN(n691) );
  AND2_X1 U603 ( .A1(n693), .A2(n691), .ZN(n535) );
  AND2_X1 U604 ( .A1(n695), .A2(n535), .ZN(G160) );
  NAND2_X1 U605 ( .A1(G138), .A2(n890), .ZN(n540) );
  AND2_X1 U606 ( .A1(G102), .A2(n891), .ZN(n539) );
  NAND2_X1 U607 ( .A1(G114), .A2(n886), .ZN(n537) );
  NAND2_X1 U608 ( .A1(G126), .A2(n887), .ZN(n536) );
  NAND2_X1 U609 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U610 ( .A1(n539), .A2(n538), .ZN(n688) );
  AND2_X1 U611 ( .A1(n540), .A2(n688), .ZN(G164) );
  INV_X1 U612 ( .A(G651), .ZN(n545) );
  NOR2_X1 U613 ( .A1(G543), .A2(n545), .ZN(n541) );
  XOR2_X2 U614 ( .A(KEYINPUT1), .B(n541), .Z(n650) );
  NAND2_X1 U615 ( .A1(G64), .A2(n650), .ZN(n544) );
  NOR2_X1 U616 ( .A1(n652), .A2(G651), .ZN(n542) );
  XNOR2_X1 U617 ( .A(KEYINPUT64), .B(n542), .ZN(n575) );
  BUF_X1 U618 ( .A(n575), .Z(n646) );
  NAND2_X1 U619 ( .A1(G52), .A2(n646), .ZN(n543) );
  NAND2_X1 U620 ( .A1(n544), .A2(n543), .ZN(n551) );
  NAND2_X1 U621 ( .A1(G77), .A2(n636), .ZN(n547) );
  NAND2_X1 U622 ( .A1(G90), .A2(n640), .ZN(n546) );
  NAND2_X1 U623 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U624 ( .A(KEYINPUT9), .B(n548), .ZN(n549) );
  XNOR2_X1 U625 ( .A(KEYINPUT69), .B(n549), .ZN(n550) );
  NOR2_X1 U626 ( .A1(n551), .A2(n550), .ZN(G171) );
  AND2_X1 U627 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U628 ( .A(G57), .ZN(G237) );
  INV_X1 U629 ( .A(G108), .ZN(G238) );
  INV_X1 U630 ( .A(G132), .ZN(G219) );
  INV_X1 U631 ( .A(G82), .ZN(G220) );
  NAND2_X1 U632 ( .A1(n636), .A2(G75), .ZN(n552) );
  XNOR2_X1 U633 ( .A(n552), .B(KEYINPUT80), .ZN(n554) );
  NAND2_X1 U634 ( .A1(G62), .A2(n650), .ZN(n553) );
  NAND2_X1 U635 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U636 ( .A1(G88), .A2(n640), .ZN(n556) );
  NAND2_X1 U637 ( .A1(G50), .A2(n575), .ZN(n555) );
  NAND2_X1 U638 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U639 ( .A1(n558), .A2(n557), .ZN(G166) );
  NAND2_X1 U640 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U641 ( .A(n559), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U642 ( .A(G567), .ZN(n681) );
  NOR2_X1 U643 ( .A1(G223), .A2(n681), .ZN(n561) );
  XNOR2_X1 U644 ( .A(KEYINPUT11), .B(KEYINPUT72), .ZN(n560) );
  XNOR2_X1 U645 ( .A(n561), .B(n560), .ZN(G234) );
  XOR2_X1 U646 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n563) );
  NAND2_X1 U647 ( .A1(G56), .A2(n650), .ZN(n562) );
  XNOR2_X1 U648 ( .A(n563), .B(n562), .ZN(n572) );
  NAND2_X1 U649 ( .A1(n575), .A2(G43), .ZN(n564) );
  XNOR2_X1 U650 ( .A(n564), .B(KEYINPUT74), .ZN(n570) );
  NAND2_X1 U651 ( .A1(G68), .A2(n636), .ZN(n567) );
  NAND2_X1 U652 ( .A1(n640), .A2(G81), .ZN(n565) );
  XNOR2_X1 U653 ( .A(n565), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U654 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U655 ( .A(n568), .B(KEYINPUT13), .ZN(n569) );
  AND2_X1 U656 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U657 ( .A1(n572), .A2(n571), .ZN(n990) );
  INV_X1 U658 ( .A(G860), .ZN(n603) );
  OR2_X1 U659 ( .A1(n990), .A2(n603), .ZN(G153) );
  INV_X1 U660 ( .A(G171), .ZN(G301) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n582) );
  NAND2_X1 U662 ( .A1(G79), .A2(n636), .ZN(n574) );
  NAND2_X1 U663 ( .A1(G92), .A2(n640), .ZN(n573) );
  NAND2_X1 U664 ( .A1(n574), .A2(n573), .ZN(n579) );
  NAND2_X1 U665 ( .A1(G66), .A2(n650), .ZN(n577) );
  NAND2_X1 U666 ( .A1(G54), .A2(n575), .ZN(n576) );
  NAND2_X1 U667 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U668 ( .A1(n579), .A2(n578), .ZN(n580) );
  INV_X1 U669 ( .A(G868), .ZN(n664) );
  NAND2_X1 U670 ( .A1(n985), .A2(n664), .ZN(n581) );
  NAND2_X1 U671 ( .A1(n582), .A2(n581), .ZN(G284) );
  NAND2_X1 U672 ( .A1(G78), .A2(n636), .ZN(n584) );
  NAND2_X1 U673 ( .A1(G91), .A2(n640), .ZN(n583) );
  NAND2_X1 U674 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U675 ( .A1(G65), .A2(n650), .ZN(n586) );
  NAND2_X1 U676 ( .A1(G53), .A2(n575), .ZN(n585) );
  NAND2_X1 U677 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U678 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U679 ( .A(n589), .B(KEYINPUT70), .ZN(n998) );
  XNOR2_X1 U680 ( .A(KEYINPUT71), .B(n998), .ZN(G299) );
  NAND2_X1 U681 ( .A1(G63), .A2(n650), .ZN(n591) );
  NAND2_X1 U682 ( .A1(G51), .A2(n646), .ZN(n590) );
  NAND2_X1 U683 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U684 ( .A(KEYINPUT6), .B(n592), .ZN(n599) );
  NAND2_X1 U685 ( .A1(n640), .A2(G89), .ZN(n593) );
  XNOR2_X1 U686 ( .A(n593), .B(KEYINPUT4), .ZN(n595) );
  NAND2_X1 U687 ( .A1(G76), .A2(n636), .ZN(n594) );
  NAND2_X1 U688 ( .A1(n595), .A2(n594), .ZN(n597) );
  NOR2_X1 U689 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U690 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U691 ( .A1(G299), .A2(G868), .ZN(n602) );
  NOR2_X1 U692 ( .A1(G286), .A2(n664), .ZN(n601) );
  NOR2_X1 U693 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U694 ( .A1(n603), .A2(G559), .ZN(n604) );
  INV_X1 U695 ( .A(n985), .ZN(n624) );
  NAND2_X1 U696 ( .A1(n604), .A2(n624), .ZN(n605) );
  XNOR2_X1 U697 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U698 ( .A1(G868), .A2(n990), .ZN(n608) );
  NAND2_X1 U699 ( .A1(G868), .A2(n624), .ZN(n606) );
  NOR2_X1 U700 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U701 ( .A1(n608), .A2(n607), .ZN(G282) );
  XOR2_X1 U702 ( .A(G2100), .B(KEYINPUT76), .Z(n617) );
  NAND2_X1 U703 ( .A1(G135), .A2(n890), .ZN(n610) );
  NAND2_X1 U704 ( .A1(G111), .A2(n886), .ZN(n609) );
  NAND2_X1 U705 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U706 ( .A1(n887), .A2(G123), .ZN(n611) );
  XOR2_X1 U707 ( .A(KEYINPUT18), .B(n611), .Z(n612) );
  NOR2_X1 U708 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U709 ( .A1(n891), .A2(G99), .ZN(n614) );
  NAND2_X1 U710 ( .A1(n615), .A2(n614), .ZN(n948) );
  XOR2_X1 U711 ( .A(G2096), .B(n948), .Z(n616) );
  NAND2_X1 U712 ( .A1(n617), .A2(n616), .ZN(G156) );
  NAND2_X1 U713 ( .A1(G67), .A2(n650), .ZN(n619) );
  NAND2_X1 U714 ( .A1(G55), .A2(n646), .ZN(n618) );
  NAND2_X1 U715 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U716 ( .A1(G80), .A2(n636), .ZN(n621) );
  NAND2_X1 U717 ( .A1(G93), .A2(n640), .ZN(n620) );
  NAND2_X1 U718 ( .A1(n621), .A2(n620), .ZN(n622) );
  OR2_X1 U719 ( .A1(n623), .A2(n622), .ZN(n665) );
  NAND2_X1 U720 ( .A1(G559), .A2(n624), .ZN(n625) );
  XNOR2_X1 U721 ( .A(n625), .B(n990), .ZN(n662) );
  NOR2_X1 U722 ( .A1(G860), .A2(n662), .ZN(n626) );
  XOR2_X1 U723 ( .A(KEYINPUT77), .B(n626), .Z(n627) );
  XOR2_X1 U724 ( .A(n665), .B(n627), .Z(G145) );
  NAND2_X1 U725 ( .A1(G73), .A2(n636), .ZN(n628) );
  XOR2_X1 U726 ( .A(KEYINPUT2), .B(n628), .Z(n633) );
  NAND2_X1 U727 ( .A1(G86), .A2(n640), .ZN(n630) );
  NAND2_X1 U728 ( .A1(G61), .A2(n650), .ZN(n629) );
  NAND2_X1 U729 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U730 ( .A(KEYINPUT79), .B(n631), .Z(n632) );
  NOR2_X1 U731 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U732 ( .A1(G48), .A2(n575), .ZN(n634) );
  NAND2_X1 U733 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U734 ( .A1(G72), .A2(n636), .ZN(n637) );
  XNOR2_X1 U735 ( .A(n637), .B(KEYINPUT68), .ZN(n639) );
  NAND2_X1 U736 ( .A1(n650), .A2(G60), .ZN(n638) );
  NAND2_X1 U737 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U738 ( .A1(G85), .A2(n640), .ZN(n641) );
  XNOR2_X1 U739 ( .A(KEYINPUT67), .B(n641), .ZN(n642) );
  NOR2_X1 U740 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U741 ( .A1(G47), .A2(n646), .ZN(n644) );
  NAND2_X1 U742 ( .A1(n645), .A2(n644), .ZN(G290) );
  NAND2_X1 U743 ( .A1(G651), .A2(G74), .ZN(n648) );
  NAND2_X1 U744 ( .A1(G49), .A2(n646), .ZN(n647) );
  NAND2_X1 U745 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U746 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U747 ( .A(n651), .B(KEYINPUT78), .ZN(n654) );
  NAND2_X1 U748 ( .A1(G87), .A2(n652), .ZN(n653) );
  NAND2_X1 U749 ( .A1(n654), .A2(n653), .ZN(G288) );
  XNOR2_X1 U750 ( .A(KEYINPUT19), .B(KEYINPUT81), .ZN(n656) );
  XNOR2_X1 U751 ( .A(G305), .B(KEYINPUT82), .ZN(n655) );
  XNOR2_X1 U752 ( .A(n656), .B(n655), .ZN(n657) );
  XOR2_X1 U753 ( .A(n665), .B(n657), .Z(n659) );
  XNOR2_X1 U754 ( .A(G290), .B(G166), .ZN(n658) );
  XNOR2_X1 U755 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U756 ( .A(G299), .B(n660), .ZN(n661) );
  XNOR2_X1 U757 ( .A(n661), .B(G288), .ZN(n914) );
  XNOR2_X1 U758 ( .A(n662), .B(n914), .ZN(n663) );
  NAND2_X1 U759 ( .A1(n663), .A2(G868), .ZN(n667) );
  NAND2_X1 U760 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U761 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U762 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U763 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U764 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U765 ( .A(n670), .B(KEYINPUT84), .ZN(n672) );
  XOR2_X1 U766 ( .A(KEYINPUT21), .B(KEYINPUT83), .Z(n671) );
  XNOR2_X1 U767 ( .A(n672), .B(n671), .ZN(n673) );
  NAND2_X1 U768 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U769 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U770 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U771 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U772 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U773 ( .A1(G96), .A2(n676), .ZN(n846) );
  NAND2_X1 U774 ( .A1(G2106), .A2(n846), .ZN(n677) );
  XNOR2_X1 U775 ( .A(n677), .B(KEYINPUT85), .ZN(n683) );
  NAND2_X1 U776 ( .A1(G120), .A2(G69), .ZN(n678) );
  NOR2_X1 U777 ( .A1(G237), .A2(n678), .ZN(n679) );
  XOR2_X1 U778 ( .A(KEYINPUT86), .B(n679), .Z(n680) );
  NOR2_X1 U779 ( .A1(G238), .A2(n680), .ZN(n848) );
  NOR2_X1 U780 ( .A1(n681), .A2(n848), .ZN(n682) );
  NOR2_X1 U781 ( .A1(n683), .A2(n682), .ZN(G319) );
  INV_X1 U782 ( .A(G319), .ZN(n685) );
  NAND2_X1 U783 ( .A1(G661), .A2(G483), .ZN(n684) );
  NOR2_X1 U784 ( .A1(n685), .A2(n684), .ZN(n845) );
  NAND2_X1 U785 ( .A1(n845), .A2(G36), .ZN(G176) );
  INV_X1 U786 ( .A(G166), .ZN(G303) );
  INV_X1 U787 ( .A(G1384), .ZN(n686) );
  AND2_X1 U788 ( .A1(G138), .A2(n686), .ZN(n687) );
  NAND2_X1 U789 ( .A1(n890), .A2(n687), .ZN(n690) );
  NAND2_X1 U790 ( .A1(n690), .A2(n689), .ZN(n788) );
  INV_X1 U791 ( .A(n788), .ZN(n701) );
  AND2_X1 U792 ( .A1(n691), .A2(G40), .ZN(n692) );
  AND2_X1 U793 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U794 ( .A1(G2084), .A2(n745), .ZN(n741) );
  INV_X1 U795 ( .A(G8), .ZN(n696) );
  NOR2_X1 U796 ( .A1(n741), .A2(n696), .ZN(n697) );
  NAND2_X1 U797 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U798 ( .A(KEYINPUT30), .B(n699), .ZN(n700) );
  NOR2_X1 U799 ( .A1(G168), .A2(n700), .ZN(n705) );
  XOR2_X1 U800 ( .A(G2078), .B(KEYINPUT25), .Z(n967) );
  NOR2_X1 U801 ( .A1(n967), .A2(n745), .ZN(n703) );
  NOR2_X1 U802 ( .A1(n719), .A2(G1961), .ZN(n702) );
  NOR2_X1 U803 ( .A1(n703), .A2(n702), .ZN(n732) );
  AND2_X1 U804 ( .A1(G301), .A2(n732), .ZN(n704) );
  XNOR2_X1 U805 ( .A(n707), .B(n706), .ZN(n735) );
  AND2_X1 U806 ( .A1(n745), .A2(G1341), .ZN(n708) );
  NOR2_X1 U807 ( .A1(n708), .A2(n990), .ZN(n711) );
  AND2_X1 U808 ( .A1(n719), .A2(G1996), .ZN(n709) );
  XOR2_X1 U809 ( .A(n709), .B(KEYINPUT26), .Z(n710) );
  NAND2_X1 U810 ( .A1(n711), .A2(n710), .ZN(n715) );
  NAND2_X1 U811 ( .A1(G1348), .A2(n745), .ZN(n713) );
  NAND2_X1 U812 ( .A1(G2067), .A2(n719), .ZN(n712) );
  NAND2_X1 U813 ( .A1(n713), .A2(n712), .ZN(n716) );
  OR2_X1 U814 ( .A1(n985), .A2(n716), .ZN(n714) );
  NAND2_X1 U815 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U816 ( .A1(n985), .A2(n716), .ZN(n717) );
  NAND2_X1 U817 ( .A1(n718), .A2(n717), .ZN(n724) );
  NAND2_X1 U818 ( .A1(n719), .A2(G2072), .ZN(n720) );
  XNOR2_X1 U819 ( .A(n720), .B(KEYINPUT27), .ZN(n722) );
  XNOR2_X1 U820 ( .A(G1956), .B(KEYINPUT95), .ZN(n1016) );
  NOR2_X1 U821 ( .A1(n1016), .A2(n719), .ZN(n721) );
  NAND2_X1 U822 ( .A1(n725), .A2(n998), .ZN(n723) );
  NAND2_X1 U823 ( .A1(n724), .A2(n723), .ZN(n729) );
  NOR2_X1 U824 ( .A1(n725), .A2(n998), .ZN(n727) );
  INV_X1 U825 ( .A(KEYINPUT28), .ZN(n726) );
  XNOR2_X1 U826 ( .A(n727), .B(n726), .ZN(n728) );
  NAND2_X1 U827 ( .A1(n729), .A2(n728), .ZN(n731) );
  NAND2_X1 U828 ( .A1(n733), .A2(n521), .ZN(n734) );
  NAND2_X1 U829 ( .A1(n735), .A2(n734), .ZN(n744) );
  INV_X1 U830 ( .A(KEYINPUT96), .ZN(n736) );
  XNOR2_X1 U831 ( .A(n744), .B(n736), .ZN(n738) );
  NOR2_X1 U832 ( .A1(G1966), .A2(n782), .ZN(n737) );
  XNOR2_X1 U833 ( .A(n740), .B(n739), .ZN(n742) );
  NAND2_X1 U834 ( .A1(n742), .A2(n523), .ZN(n743) );
  XNOR2_X1 U835 ( .A(n743), .B(KEYINPUT98), .ZN(n754) );
  NAND2_X1 U836 ( .A1(G286), .A2(n744), .ZN(n750) );
  NOR2_X1 U837 ( .A1(G1971), .A2(n782), .ZN(n747) );
  NOR2_X1 U838 ( .A1(G2090), .A2(n745), .ZN(n746) );
  NOR2_X1 U839 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U840 ( .A1(n748), .A2(G303), .ZN(n749) );
  NAND2_X1 U841 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U842 ( .A1(G8), .A2(n751), .ZN(n752) );
  XNOR2_X1 U843 ( .A(KEYINPUT32), .B(n752), .ZN(n753) );
  NOR2_X1 U844 ( .A1(G1971), .A2(G303), .ZN(n755) );
  XNOR2_X1 U845 ( .A(n755), .B(KEYINPUT99), .ZN(n757) );
  NOR2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n996) );
  NAND2_X1 U847 ( .A1(n776), .A2(n758), .ZN(n759) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n993) );
  NAND2_X1 U849 ( .A1(n759), .A2(n993), .ZN(n761) );
  XNOR2_X1 U850 ( .A(n761), .B(n760), .ZN(n763) );
  INV_X1 U851 ( .A(n782), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n522), .A2(n767), .ZN(n765) );
  INV_X1 U853 ( .A(KEYINPUT33), .ZN(n764) );
  NAND2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n773) );
  INV_X1 U855 ( .A(KEYINPUT101), .ZN(n767) );
  NAND2_X1 U856 ( .A1(n996), .A2(KEYINPUT33), .ZN(n766) );
  NAND2_X1 U857 ( .A1(n767), .A2(n766), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n996), .A2(KEYINPUT101), .ZN(n768) );
  NAND2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U860 ( .A1(n782), .A2(n770), .ZN(n772) );
  XOR2_X1 U861 ( .A(G1981), .B(G305), .Z(n1002) );
  NAND2_X1 U862 ( .A1(n773), .A2(n525), .ZN(n774) );
  XNOR2_X1 U863 ( .A(n774), .B(KEYINPUT102), .ZN(n785) );
  NOR2_X1 U864 ( .A1(G2090), .A2(G303), .ZN(n775) );
  NAND2_X1 U865 ( .A1(G8), .A2(n775), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n778), .A2(n782), .ZN(n783) );
  NOR2_X1 U868 ( .A1(G1981), .A2(G305), .ZN(n779) );
  XOR2_X1 U869 ( .A(n779), .B(KEYINPUT24), .Z(n780) );
  XNOR2_X1 U870 ( .A(KEYINPUT94), .B(n780), .ZN(n781) );
  XNOR2_X1 U871 ( .A(n786), .B(KEYINPUT103), .ZN(n823) );
  NOR2_X1 U872 ( .A1(n788), .A2(n787), .ZN(n836) );
  NAND2_X1 U873 ( .A1(n891), .A2(G105), .ZN(n790) );
  XNOR2_X1 U874 ( .A(KEYINPUT38), .B(KEYINPUT90), .ZN(n789) );
  XNOR2_X1 U875 ( .A(n790), .B(n789), .ZN(n797) );
  NAND2_X1 U876 ( .A1(G117), .A2(n886), .ZN(n792) );
  NAND2_X1 U877 ( .A1(G129), .A2(n887), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U879 ( .A1(G141), .A2(n890), .ZN(n793) );
  XNOR2_X1 U880 ( .A(KEYINPUT91), .B(n793), .ZN(n794) );
  NOR2_X1 U881 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U882 ( .A1(n797), .A2(n796), .ZN(n910) );
  NAND2_X1 U883 ( .A1(n910), .A2(G1996), .ZN(n807) );
  NAND2_X1 U884 ( .A1(G131), .A2(n890), .ZN(n799) );
  NAND2_X1 U885 ( .A1(G119), .A2(n887), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U887 ( .A1(n886), .A2(G107), .ZN(n800) );
  XOR2_X1 U888 ( .A(KEYINPUT88), .B(n800), .Z(n801) );
  NOR2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n804) );
  NAND2_X1 U890 ( .A1(n891), .A2(G95), .ZN(n803) );
  NAND2_X1 U891 ( .A1(n804), .A2(n803), .ZN(n899) );
  NAND2_X1 U892 ( .A1(G1991), .A2(n899), .ZN(n805) );
  XOR2_X1 U893 ( .A(KEYINPUT89), .B(n805), .Z(n806) );
  NAND2_X1 U894 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U895 ( .A(n808), .B(KEYINPUT92), .ZN(n947) );
  NAND2_X1 U896 ( .A1(n836), .A2(n947), .ZN(n826) );
  NAND2_X1 U897 ( .A1(G140), .A2(n890), .ZN(n810) );
  NAND2_X1 U898 ( .A1(G104), .A2(n891), .ZN(n809) );
  NAND2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U900 ( .A(KEYINPUT34), .B(n811), .ZN(n816) );
  NAND2_X1 U901 ( .A1(G116), .A2(n886), .ZN(n813) );
  NAND2_X1 U902 ( .A1(G128), .A2(n887), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U904 ( .A(KEYINPUT35), .B(n814), .Z(n815) );
  NOR2_X1 U905 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U906 ( .A(KEYINPUT36), .B(n817), .ZN(n911) );
  XNOR2_X1 U907 ( .A(KEYINPUT37), .B(G2067), .ZN(n834) );
  NOR2_X1 U908 ( .A1(n911), .A2(n834), .ZN(n943) );
  NAND2_X1 U909 ( .A1(n836), .A2(n943), .ZN(n833) );
  NAND2_X1 U910 ( .A1(n826), .A2(n833), .ZN(n818) );
  XOR2_X1 U911 ( .A(KEYINPUT93), .B(n818), .Z(n821) );
  XNOR2_X1 U912 ( .A(G1986), .B(G290), .ZN(n987) );
  NAND2_X1 U913 ( .A1(n836), .A2(n987), .ZN(n819) );
  XNOR2_X1 U914 ( .A(KEYINPUT87), .B(n819), .ZN(n820) );
  NOR2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n839) );
  NOR2_X1 U917 ( .A1(G1996), .A2(n910), .ZN(n940) );
  NOR2_X1 U918 ( .A1(G1991), .A2(n899), .ZN(n956) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n824) );
  NOR2_X1 U920 ( .A1(n956), .A2(n824), .ZN(n825) );
  XOR2_X1 U921 ( .A(KEYINPUT104), .B(n825), .Z(n827) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U923 ( .A(KEYINPUT105), .B(n828), .ZN(n829) );
  NOR2_X1 U924 ( .A1(n940), .A2(n829), .ZN(n831) );
  XNOR2_X1 U925 ( .A(KEYINPUT39), .B(KEYINPUT106), .ZN(n830) );
  XNOR2_X1 U926 ( .A(n831), .B(n830), .ZN(n832) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n911), .A2(n834), .ZN(n949) );
  NAND2_X1 U929 ( .A1(n835), .A2(n949), .ZN(n837) );
  NAND2_X1 U930 ( .A1(n837), .A2(n836), .ZN(n838) );
  NAND2_X1 U931 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U932 ( .A(n840), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U933 ( .A(G223), .ZN(n841) );
  NAND2_X1 U934 ( .A1(n841), .A2(G2106), .ZN(n842) );
  XOR2_X1 U935 ( .A(KEYINPUT107), .B(n842), .Z(G217) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U937 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U939 ( .A1(n845), .A2(n844), .ZN(G188) );
  INV_X1 U941 ( .A(G120), .ZN(G236) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(G69), .ZN(G235) );
  INV_X1 U944 ( .A(n846), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n848), .A2(n847), .ZN(G261) );
  INV_X1 U946 ( .A(G261), .ZN(G325) );
  XOR2_X1 U947 ( .A(KEYINPUT109), .B(KEYINPUT108), .Z(n850) );
  XNOR2_X1 U948 ( .A(G2678), .B(KEYINPUT43), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U950 ( .A(KEYINPUT42), .B(G2072), .Z(n852) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2090), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U953 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U954 ( .A(G2100), .B(G2096), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n858) );
  XOR2_X1 U956 ( .A(G2078), .B(G2084), .Z(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(G227) );
  XOR2_X1 U958 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n860) );
  XNOR2_X1 U959 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U961 ( .A(n861), .B(G2474), .Z(n863) );
  XNOR2_X1 U962 ( .A(G1996), .B(G1991), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n871) );
  XOR2_X1 U964 ( .A(G1976), .B(G1966), .Z(n865) );
  XNOR2_X1 U965 ( .A(G1971), .B(G1956), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U967 ( .A(KEYINPUT112), .B(G1981), .Z(n867) );
  XNOR2_X1 U968 ( .A(G1986), .B(G1961), .ZN(n866) );
  XNOR2_X1 U969 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U970 ( .A(n869), .B(n868), .Z(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(G229) );
  NAND2_X1 U972 ( .A1(G124), .A2(n887), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n872), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U974 ( .A1(n886), .A2(G112), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G136), .A2(n890), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G100), .A2(n891), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U979 ( .A1(n878), .A2(n877), .ZN(G162) );
  NAND2_X1 U980 ( .A1(G139), .A2(n890), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G103), .A2(n891), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G115), .A2(n886), .ZN(n882) );
  NAND2_X1 U984 ( .A1(G127), .A2(n887), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U986 ( .A(KEYINPUT47), .B(n883), .Z(n884) );
  NOR2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n935) );
  XNOR2_X1 U988 ( .A(G160), .B(G162), .ZN(n898) );
  NAND2_X1 U989 ( .A1(G118), .A2(n886), .ZN(n889) );
  NAND2_X1 U990 ( .A1(G130), .A2(n887), .ZN(n888) );
  NAND2_X1 U991 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U992 ( .A1(G142), .A2(n890), .ZN(n893) );
  NAND2_X1 U993 ( .A1(G106), .A2(n891), .ZN(n892) );
  NAND2_X1 U994 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U995 ( .A(KEYINPUT45), .B(n894), .Z(n895) );
  NOR2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n902) );
  XNOR2_X1 U998 ( .A(G164), .B(n899), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n900), .B(n948), .ZN(n901) );
  XOR2_X1 U1000 ( .A(n902), .B(n901), .Z(n907) );
  XOR2_X1 U1001 ( .A(KEYINPUT116), .B(KEYINPUT114), .Z(n904) );
  XNOR2_X1 U1002 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(KEYINPUT46), .B(n905), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1006 ( .A(n935), .B(n908), .Z(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n912) );
  XOR2_X1 U1008 ( .A(n912), .B(n911), .Z(n913) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n913), .ZN(G395) );
  XNOR2_X1 U1010 ( .A(G171), .B(n985), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(n990), .B(G286), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n918), .ZN(G397) );
  XOR2_X1 U1015 ( .A(G2451), .B(G2430), .Z(n920) );
  XNOR2_X1 U1016 ( .A(G2438), .B(G2443), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(n920), .B(n919), .ZN(n926) );
  XOR2_X1 U1018 ( .A(G2435), .B(G2454), .Z(n922) );
  XNOR2_X1 U1019 ( .A(G1341), .B(G1348), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(n922), .B(n921), .ZN(n924) );
  XOR2_X1 U1021 ( .A(G2446), .B(G2427), .Z(n923) );
  XNOR2_X1 U1022 ( .A(n924), .B(n923), .ZN(n925) );
  XOR2_X1 U1023 ( .A(n926), .B(n925), .Z(n927) );
  NAND2_X1 U1024 ( .A1(G14), .A2(n927), .ZN(n934) );
  NAND2_X1 U1025 ( .A1(G319), .A2(n934), .ZN(n931) );
  NOR2_X1 U1026 ( .A1(G227), .A2(G229), .ZN(n928) );
  XOR2_X1 U1027 ( .A(KEYINPUT117), .B(n928), .Z(n929) );
  XNOR2_X1 U1028 ( .A(n929), .B(KEYINPUT49), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n933) );
  NOR2_X1 U1030 ( .A1(G395), .A2(G397), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(G225) );
  INV_X1 U1032 ( .A(G225), .ZN(G308) );
  INV_X1 U1033 ( .A(n934), .ZN(G401) );
  XNOR2_X1 U1034 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n958) );
  XOR2_X1 U1035 ( .A(G2072), .B(n935), .Z(n937) );
  XOR2_X1 U1036 ( .A(G164), .B(G2078), .Z(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(KEYINPUT50), .B(n938), .ZN(n945) );
  XOR2_X1 U1039 ( .A(G2090), .B(G162), .Z(n939) );
  NOR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1041 ( .A(n941), .B(KEYINPUT51), .ZN(n942) );
  NOR2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n954) );
  NAND2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n952) );
  XOR2_X1 U1046 ( .A(G2084), .B(G160), .Z(n950) );
  XNOR2_X1 U1047 ( .A(KEYINPUT118), .B(n950), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n958), .B(n957), .ZN(n959) );
  OR2_X1 U1052 ( .A1(KEYINPUT55), .A2(n959), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n960), .A2(G29), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(n961), .B(KEYINPUT120), .ZN(n1041) );
  XOR2_X1 U1055 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n981) );
  XNOR2_X1 U1056 ( .A(G2090), .B(G35), .ZN(n976) );
  XOR2_X1 U1057 ( .A(G2072), .B(G33), .Z(n962) );
  NAND2_X1 U1058 ( .A1(n962), .A2(G28), .ZN(n973) );
  XNOR2_X1 U1059 ( .A(G25), .B(G1991), .ZN(n963) );
  XNOR2_X1 U1060 ( .A(n963), .B(KEYINPUT121), .ZN(n971) );
  XOR2_X1 U1061 ( .A(G2067), .B(G26), .Z(n966) );
  INV_X1 U1062 ( .A(G1996), .ZN(n964) );
  XNOR2_X1 U1063 ( .A(n964), .B(G32), .ZN(n965) );
  NAND2_X1 U1064 ( .A1(n966), .A2(n965), .ZN(n969) );
  XNOR2_X1 U1065 ( .A(G27), .B(n967), .ZN(n968) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(KEYINPUT53), .B(n974), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n979) );
  XOR2_X1 U1071 ( .A(G2084), .B(G34), .Z(n977) );
  XNOR2_X1 U1072 ( .A(KEYINPUT54), .B(n977), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(n981), .B(n980), .ZN(n983) );
  INV_X1 U1075 ( .A(G29), .ZN(n982) );
  NAND2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(G11), .A2(n984), .ZN(n1039) );
  XNOR2_X1 U1078 ( .A(G16), .B(KEYINPUT56), .ZN(n1011) );
  XNOR2_X1 U1079 ( .A(G171), .B(G1961), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(G1348), .B(n985), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(G1341), .B(n990), .ZN(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n1009) );
  XNOR2_X1 U1085 ( .A(G166), .B(G1971), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1088 ( .A(KEYINPUT124), .B(n997), .Z(n1000) );
  XOR2_X1 U1089 ( .A(n998), .B(G1956), .Z(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(KEYINPUT125), .B(n1001), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(G168), .B(G1966), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(n1004), .B(KEYINPUT123), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(KEYINPUT57), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1037) );
  INV_X1 U1099 ( .A(G16), .ZN(n1035) );
  XNOR2_X1 U1100 ( .A(G1961), .B(G5), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(G1966), .B(G21), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1025) );
  XOR2_X1 U1103 ( .A(KEYINPUT126), .B(G4), .Z(n1015) );
  XNOR2_X1 U1104 ( .A(G1348), .B(KEYINPUT59), .ZN(n1014) );
  XNOR2_X1 U1105 ( .A(n1015), .B(n1014), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(G20), .B(n1016), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(G1341), .B(G19), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(G1981), .B(G6), .ZN(n1017) );
  NOR2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1112 ( .A(n1023), .B(KEYINPUT60), .ZN(n1024) );
  NAND2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1032) );
  XNOR2_X1 U1114 ( .A(G1971), .B(G22), .ZN(n1027) );
  XNOR2_X1 U1115 ( .A(G23), .B(G1976), .ZN(n1026) );
  NOR2_X1 U1116 ( .A1(n1027), .A2(n1026), .ZN(n1029) );
  XOR2_X1 U1117 ( .A(G1986), .B(G24), .Z(n1028) );
  NAND2_X1 U1118 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1119 ( .A(KEYINPUT58), .B(n1030), .ZN(n1031) );
  NOR2_X1 U1120 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1121 ( .A(KEYINPUT61), .B(n1033), .ZN(n1034) );
  NAND2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1123 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NOR2_X1 U1124 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NAND2_X1 U1125 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XOR2_X1 U1126 ( .A(KEYINPUT62), .B(n1042), .Z(G311) );
  INV_X1 U1127 ( .A(G311), .ZN(G150) );
endmodule

