//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203));
  AOI21_X1  g002(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT89), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(G71gat), .A2(G78gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n208), .ZN(new_n210));
  OR2_X1    g009(.A1(G57gat), .A2(G64gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G57gat), .A2(G64gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n211), .B(new_n212), .C1(new_n206), .C2(KEYINPUT9), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n210), .B1(new_n213), .B2(KEYINPUT89), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n202), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n205), .A2(new_n208), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n210), .A2(new_n213), .A3(KEYINPUT89), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT90), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(KEYINPUT21), .ZN(new_n220));
  XOR2_X1   g019(.A(G127gat), .B(G155gat), .Z(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(G15gat), .B(G22gat), .Z(new_n224));
  INV_X1    g023(.A(G1gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(G1gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n229), .A3(KEYINPUT84), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n230), .A2(G8gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(G8gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n233), .B1(new_n219), .B2(KEYINPUT21), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(KEYINPUT91), .ZN(new_n235));
  AND2_X1   g034(.A1(G231gat), .A2(G233gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n235), .A2(new_n236), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n223), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n239), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(new_n237), .A3(new_n222), .ZN(new_n242));
  XOR2_X1   g041(.A(G183gat), .B(G211gat), .Z(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n240), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n245), .B1(new_n240), .B2(new_n242), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT95), .ZN(new_n250));
  NAND2_X1  g049(.A1(G232gat), .A2(G233gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT92), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT41), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n254), .B(KEYINPUT93), .Z(new_n255));
  INV_X1    g054(.A(KEYINPUT83), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT14), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n256), .B(new_n257), .C1(G29gat), .C2(G36gat), .ZN(new_n258));
  INV_X1    g057(.A(G29gat), .ZN(new_n259));
  INV_X1    g058(.A(G36gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(G29gat), .A2(G36gat), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n257), .B1(new_n262), .B2(KEYINPUT83), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n256), .B1(G29gat), .B2(G36gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(G43gat), .B(G50gat), .Z(new_n266));
  INV_X1    g065(.A(KEYINPUT15), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n267), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n265), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n263), .A2(new_n264), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n268), .B1(new_n272), .B2(new_n261), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT17), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n271), .A2(KEYINPUT17), .A3(new_n273), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G99gat), .A2(G106gat), .ZN(new_n279));
  INV_X1    g078(.A(G85gat), .ZN(new_n280));
  INV_X1    g079(.A(G92gat), .ZN(new_n281));
  AOI22_X1  g080(.A1(KEYINPUT8), .A2(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT7), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(new_n280), .B2(new_n281), .ZN(new_n284));
  NAND3_X1  g083(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n282), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G99gat), .B(G106gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n278), .A2(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G190gat), .B(G218gat), .Z(new_n291));
  INV_X1    g090(.A(KEYINPUT94), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI22_X1  g092(.A1(new_n252), .A2(new_n253), .B1(new_n291), .B2(new_n292), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n294), .B1(new_n274), .B2(new_n288), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n290), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n293), .B1(new_n290), .B2(new_n295), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n255), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n298), .ZN(new_n300));
  INV_X1    g099(.A(new_n255), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n301), .A3(new_n296), .ZN(new_n302));
  XNOR2_X1  g101(.A(G134gat), .B(G162gat), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n299), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n303), .B1(new_n299), .B2(new_n302), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n249), .A2(new_n250), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n306), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT95), .B1(new_n248), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G230gat), .A2(G233gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT97), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n286), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n288), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n287), .ZN(new_n317));
  OAI22_X1  g116(.A1(new_n209), .A2(new_n214), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT96), .B1(new_n219), .B2(new_n288), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT96), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n289), .A2(new_n321), .A3(new_n218), .A4(new_n215), .ZN(new_n322));
  AOI211_X1 g121(.A(KEYINPUT10), .B(new_n319), .C1(new_n320), .C2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n219), .A2(KEYINPUT10), .A3(new_n288), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n312), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n319), .B1(new_n320), .B2(new_n322), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n312), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G120gat), .B(G148gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(G176gat), .B(G204gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n326), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT98), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n334), .B1(new_n326), .B2(new_n330), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n337), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n308), .A2(new_n311), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n233), .B(new_n274), .ZN(new_n343));
  NAND2_X1  g142(.A1(G229gat), .A2(G233gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n344), .B(KEYINPUT13), .Z(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(KEYINPUT87), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n233), .A2(new_n274), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n231), .A2(new_n232), .B1(new_n271), .B2(new_n273), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n345), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT87), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT85), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n231), .A2(new_n353), .A3(new_n232), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n353), .B1(new_n231), .B2(new_n232), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n277), .B(new_n276), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT86), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n233), .A2(KEYINPUT85), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n231), .A2(new_n353), .A3(new_n232), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT86), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n278), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n348), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n357), .A2(new_n362), .A3(new_n344), .A4(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT18), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n352), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n348), .B1(new_n356), .B2(KEYINPUT86), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n367), .A2(KEYINPUT18), .A3(new_n344), .A4(new_n362), .ZN(new_n368));
  XNOR2_X1  g167(.A(G113gat), .B(G141gat), .ZN(new_n369));
  INV_X1    g168(.A(G197gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT11), .B(G169gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT12), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n366), .A2(new_n368), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n374), .B1(new_n366), .B2(new_n368), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT88), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n366), .A2(new_n368), .ZN(new_n378));
  INV_X1    g177(.A(new_n374), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT88), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n368), .A3(new_n374), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G8gat), .B(G36gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(G64gat), .B(G92gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G197gat), .B(G204gat), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT22), .ZN(new_n389));
  INV_X1    g188(.A(G211gat), .ZN(new_n390));
  INV_X1    g189(.A(G218gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G211gat), .B(G218gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n388), .A3(new_n392), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT28), .ZN(new_n400));
  INV_X1    g199(.A(G183gat), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT27), .B1(new_n401), .B2(KEYINPUT67), .ZN(new_n402));
  INV_X1    g201(.A(G190gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n401), .A2(KEYINPUT67), .A3(KEYINPUT27), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n400), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT27), .B(G183gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT28), .A3(new_n403), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT69), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT68), .B(KEYINPUT26), .ZN(new_n412));
  INV_X1    g211(.A(G169gat), .ZN(new_n413));
  INV_X1    g212(.A(G176gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n411), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(G169gat), .A2(G176gat), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT26), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n418), .A2(KEYINPUT68), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(KEYINPUT68), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT69), .B(new_n417), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G169gat), .A2(G176gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n423), .B1(KEYINPUT26), .B2(new_n415), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n416), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G183gat), .A2(G190gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT70), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n425), .A2(KEYINPUT70), .A3(new_n426), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n410), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT24), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(G183gat), .A2(G190gat), .ZN(new_n435));
  OR3_X1    g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n417), .A2(KEYINPUT23), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n437), .A2(KEYINPUT25), .A3(new_n422), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT23), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n415), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n436), .A2(KEYINPUT66), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT66), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n440), .A2(KEYINPUT25), .A3(new_n422), .A4(new_n437), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT25), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT65), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n437), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n417), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n436), .A2(new_n451), .A3(new_n422), .A4(new_n440), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n446), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n399), .B1(new_n431), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(G226gat), .A2(G233gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n455), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(new_n431), .B2(new_n453), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n398), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n425), .A2(KEYINPUT70), .A3(new_n426), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT70), .B1(new_n425), .B2(new_n426), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n409), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n452), .A2(new_n447), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(new_n445), .A3(new_n441), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT29), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n458), .B(new_n398), .C1(new_n465), .C2(new_n457), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n387), .B1(new_n459), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n398), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n465), .A2(new_n457), .ZN(new_n470));
  INV_X1    g269(.A(new_n458), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n387), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n466), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n468), .A2(KEYINPUT30), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT30), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n472), .A2(new_n476), .A3(new_n473), .A4(new_n466), .ZN(new_n477));
  XNOR2_X1  g276(.A(G141gat), .B(G148gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(G155gat), .A2(G162gat), .ZN(new_n479));
  NOR2_X1   g278(.A1(G155gat), .A2(G162gat), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n478), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT75), .B(G155gat), .ZN(new_n483));
  INV_X1    g282(.A(G162gat), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT2), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT74), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n479), .B1(new_n478), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n479), .ZN(new_n489));
  OAI221_X1 g288(.A(new_n481), .B1(new_n489), .B2(KEYINPUT74), .C1(new_n478), .C2(KEYINPUT2), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n486), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G113gat), .B(G120gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT72), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(KEYINPUT1), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G127gat), .B(G134gat), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT71), .B1(new_n497), .B2(new_n494), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n492), .A2(KEYINPUT1), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n496), .A2(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT4), .B1(new_n491), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n478), .A2(KEYINPUT2), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n481), .B1(new_n489), .B2(KEYINPUT74), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n488), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n504), .A2(new_n505), .B1(new_n485), .B2(new_n482), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n496), .A2(new_n497), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n498), .A2(new_n499), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT4), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n506), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n501), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n491), .A2(KEYINPUT3), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT3), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n486), .B(new_n514), .C1(new_n488), .C2(new_n490), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n500), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G225gat), .A2(G233gat), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n512), .A2(new_n516), .A3(KEYINPUT5), .A4(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n512), .A2(new_n517), .A3(new_n516), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n506), .A2(new_n509), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n491), .A2(new_n500), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT5), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n518), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  XOR2_X1   g324(.A(G57gat), .B(G85gat), .Z(new_n526));
  XNOR2_X1  g325(.A(G1gat), .B(G29gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT77), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT6), .B1(new_n525), .B2(new_n531), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n512), .A2(new_n517), .A3(new_n516), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(new_n523), .B2(new_n522), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT77), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n535), .A2(new_n536), .A3(new_n530), .A4(new_n518), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n535), .A2(KEYINPUT6), .A3(new_n530), .A4(new_n518), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n475), .A2(new_n477), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G78gat), .B(G106gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT31), .B(G50gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT29), .B1(new_n396), .B2(new_n397), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n491), .B1(KEYINPUT3), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT29), .B1(new_n506), .B2(new_n514), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n545), .B1(new_n546), .B2(new_n398), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT78), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(new_n546), .B2(new_n398), .ZN(new_n549));
  NAND2_X1  g348(.A1(G228gat), .A2(G233gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  OAI221_X1 g351(.A(new_n545), .B1(new_n548), .B2(new_n550), .C1(new_n546), .C2(new_n398), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G22gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n552), .A2(G22gat), .A3(new_n553), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n543), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n555), .A2(KEYINPUT79), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n552), .A2(new_n553), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT80), .B1(new_n555), .B2(KEYINPUT79), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(new_n552), .B2(new_n553), .ZN(new_n562));
  INV_X1    g361(.A(new_n543), .ZN(new_n563));
  NOR3_X1   g362(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT80), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n556), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n558), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n540), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT37), .B1(new_n459), .B2(new_n467), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT37), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n472), .A2(new_n571), .A3(new_n466), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n387), .A3(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n573), .A2(KEYINPUT38), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n525), .A2(KEYINPUT81), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT81), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n535), .A2(new_n576), .A3(new_n518), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n530), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n533), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n579), .A2(new_n539), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n573), .A2(KEYINPUT38), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n574), .A2(new_n580), .A3(new_n474), .A4(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n517), .B1(new_n512), .B2(new_n516), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT39), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT40), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n530), .B1(KEYINPUT82), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n520), .A2(new_n521), .A3(new_n517), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT39), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n583), .B2(new_n590), .ZN(new_n591));
  OAI22_X1  g390(.A1(new_n586), .A2(new_n591), .B1(KEYINPUT82), .B2(new_n587), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n583), .A2(new_n590), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n587), .A2(KEYINPUT82), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n585), .A4(new_n588), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n475), .A2(new_n596), .A3(new_n477), .A4(new_n578), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n597), .A2(new_n568), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n569), .B1(new_n582), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G15gat), .B(G43gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(G71gat), .B(G99gat), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  NAND2_X1  g401(.A1(G227gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT64), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n500), .B1(new_n431), .B2(new_n453), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n462), .A2(new_n509), .A3(new_n464), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n602), .B1(new_n608), .B2(KEYINPUT33), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT32), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT34), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n462), .A2(new_n509), .A3(new_n464), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n509), .B1(new_n462), .B2(new_n464), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n604), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT34), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(KEYINPUT32), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n606), .A2(new_n605), .A3(new_n607), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT73), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n611), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n619), .B1(new_n611), .B2(new_n616), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n609), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n619), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n608), .A2(new_n610), .A3(KEYINPUT34), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n615), .B1(new_n614), .B2(KEYINPUT32), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n609), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n616), .A3(new_n619), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n622), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT36), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT36), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n599), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n630), .A2(new_n540), .A3(new_n568), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT35), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n567), .B1(new_n622), .B2(new_n629), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n475), .A2(new_n477), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT35), .B1(new_n579), .B2(new_n539), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n384), .B1(new_n635), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n342), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n538), .A2(new_n539), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(new_n225), .ZN(G1324gat));
  INV_X1    g446(.A(new_n644), .ZN(new_n648));
  INV_X1    g447(.A(new_n639), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(G8gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT42), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT16), .B(G8gat), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  MUX2_X1   g453(.A(new_n652), .B(KEYINPUT42), .S(new_n654), .Z(G1325gat));
  INV_X1    g454(.A(G15gat), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n632), .A2(new_n634), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n644), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n648), .A2(new_n630), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n658), .B1(new_n656), .B2(new_n659), .ZN(G1326gat));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n568), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT43), .B(G22gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1327gat));
  NOR3_X1   g462(.A1(new_n249), .A2(new_n341), .A3(new_n306), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n643), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n645), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(new_n259), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT99), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT45), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n306), .A2(KEYINPUT44), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT35), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(new_n638), .B2(new_n540), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n673), .A2(new_n675), .A3(KEYINPUT101), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n677), .B1(new_n637), .B2(new_n641), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n635), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT102), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT101), .B1(new_n673), .B2(new_n675), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n637), .A2(new_n677), .A3(new_n641), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT102), .B1(new_n684), .B2(new_n635), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n672), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n635), .A2(new_n642), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n309), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT44), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n380), .A2(new_n382), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n248), .A2(new_n340), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT100), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n694), .A2(new_n666), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n670), .B(new_n671), .C1(new_n259), .C2(new_n695), .ZN(G1328gat));
  NAND3_X1  g495(.A1(new_n665), .A2(new_n260), .A3(new_n649), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT46), .Z(new_n698));
  NAND3_X1  g497(.A1(new_n690), .A2(new_n649), .A3(new_n693), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G36gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n698), .A2(new_n700), .A3(KEYINPUT103), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(G1329gat));
  INV_X1    g504(.A(new_n665), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n706), .A2(G43gat), .A3(new_n631), .ZN(new_n707));
  INV_X1    g506(.A(new_n657), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n690), .A2(new_n708), .A3(new_n693), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n707), .B1(new_n709), .B2(G43gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g510(.A1(new_n690), .A2(G50gat), .A3(new_n567), .A4(new_n693), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n665), .A2(KEYINPUT104), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n567), .B1(new_n665), .B2(KEYINPUT104), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n712), .B1(G50gat), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g516(.A1(new_n679), .A2(new_n680), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n684), .A2(KEYINPUT102), .A3(new_n635), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR4_X1   g519(.A1(new_n308), .A2(new_n311), .A3(new_n340), .A4(new_n691), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n666), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n649), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n726));
  XOR2_X1   g525(.A(KEYINPUT49), .B(G64gat), .Z(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT105), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n726), .B(new_n730), .C1(new_n725), .C2(new_n727), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(G1333gat));
  INV_X1    g531(.A(G71gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n720), .A2(new_n721), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n734), .B2(new_n631), .ZN(new_n735));
  NOR4_X1   g534(.A1(new_n734), .A2(KEYINPUT106), .A3(new_n733), .A4(new_n657), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n657), .A2(new_n733), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n722), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n735), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g540(.A1(new_n734), .A2(new_n568), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT107), .B(G78gat), .Z(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1335gat));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n682), .A2(new_n683), .B1(new_n657), .B2(new_n599), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n249), .A2(new_n691), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n309), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n745), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n748), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n679), .A2(KEYINPUT51), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT108), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n679), .A2(new_n750), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(new_n745), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(new_n340), .ZN(new_n757));
  AOI21_X1  g556(.A(G85gat), .B1(new_n757), .B2(new_n666), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n747), .A2(new_n341), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n686), .B2(new_n689), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n645), .A2(new_n280), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(G1336gat));
  NOR2_X1   g561(.A1(new_n639), .A2(G92gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n757), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n649), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G92gat), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n764), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n749), .A2(new_n751), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n769), .A2(new_n341), .A3(new_n763), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n765), .B2(G92gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n768), .B1(new_n767), .B2(new_n771), .ZN(G1337gat));
  INV_X1    g571(.A(G99gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n773), .A3(new_n630), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n760), .A2(new_n708), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n773), .B2(new_n775), .ZN(G1338gat));
  INV_X1    g575(.A(G106gat), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n760), .B2(new_n567), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n340), .A2(G106gat), .A3(new_n568), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n752), .B2(new_n755), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n759), .ZN(new_n784));
  INV_X1    g583(.A(new_n672), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n718), .B2(new_n719), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n688), .A2(KEYINPUT44), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n567), .B(new_n784), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G106gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n769), .A2(new_n779), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n781), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT109), .B1(new_n783), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(new_n781), .A3(new_n780), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n788), .A2(G106gat), .B1(new_n769), .B2(new_n779), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n793), .B(new_n794), .C1(new_n781), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n796), .ZN(G1339gat));
  INV_X1    g596(.A(KEYINPUT10), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n327), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n329), .B1(new_n799), .B2(new_n324), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n334), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(new_n329), .A3(new_n324), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n326), .A2(KEYINPUT54), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT110), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n802), .A2(new_n804), .A3(KEYINPUT55), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(new_n335), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n805), .A2(KEYINPUT110), .A3(new_n806), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n809), .A2(new_n811), .A3(new_n691), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n344), .B1(new_n367), .B2(new_n362), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n343), .A2(new_n345), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n373), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n338), .A2(new_n339), .A3(new_n382), .A4(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n309), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n809), .A2(new_n811), .A3(new_n812), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n382), .B(new_n816), .C1(new_n304), .C2(new_n305), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n248), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n691), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n307), .A2(new_n310), .A3(new_n340), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n649), .A2(new_n645), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(new_n638), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(KEYINPUT111), .Z(new_n829));
  INV_X1    g628(.A(G113gat), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n830), .A3(new_n691), .ZN(new_n831));
  INV_X1    g630(.A(new_n828), .ZN(new_n832));
  OAI21_X1  g631(.A(G113gat), .B1(new_n832), .B2(new_n384), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1340gat));
  INV_X1    g633(.A(G120gat), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n829), .A2(new_n835), .A3(new_n341), .ZN(new_n836));
  OAI21_X1  g635(.A(G120gat), .B1(new_n832), .B2(new_n340), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1341gat));
  NAND2_X1  g637(.A1(new_n828), .A2(new_n249), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(G127gat), .ZN(G1342gat));
  INV_X1    g639(.A(KEYINPUT56), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n832), .A2(G134gat), .A3(new_n306), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT112), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n842), .A2(new_n843), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n841), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n846), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(KEYINPUT56), .A3(new_n844), .ZN(new_n849));
  OAI21_X1  g648(.A(G134gat), .B1(new_n832), .B2(new_n306), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(G1343gat));
  INV_X1    g650(.A(new_n384), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n657), .A2(new_n826), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n567), .A2(KEYINPUT57), .ZN(new_n854));
  INV_X1    g653(.A(new_n821), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n805), .A2(KEYINPUT113), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT113), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n802), .A2(new_n804), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n806), .A3(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n859), .A2(new_n377), .A3(new_n383), .A4(new_n811), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n309), .B1(new_n860), .B2(new_n817), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n855), .B1(new_n861), .B2(KEYINPUT114), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n863));
  AOI211_X1 g662(.A(new_n863), .B(new_n309), .C1(new_n860), .C2(new_n817), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n248), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n854), .B1(new_n865), .B2(new_n824), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT57), .B1(new_n825), .B2(new_n567), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n852), .B(new_n853), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(G141gat), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n384), .A2(G141gat), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n825), .A2(new_n567), .A3(new_n853), .A4(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT116), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876));
  AOI211_X1 g675(.A(new_n876), .B(new_n873), .C1(new_n868), .C2(G141gat), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n691), .B(new_n853), .C1(new_n866), .C2(new_n867), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n879), .A2(KEYINPUT115), .A3(G141gat), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT115), .B1(new_n879), .B2(G141gat), .ZN(new_n881));
  INV_X1    g680(.A(new_n871), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n878), .B1(new_n883), .B2(new_n872), .ZN(G1344gat));
  AND3_X1   g683(.A1(new_n825), .A2(new_n567), .A3(new_n853), .ZN(new_n885));
  INV_X1    g684(.A(G148gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n886), .A3(new_n341), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n853), .B1(new_n866), .B2(new_n867), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n888), .A2(new_n340), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n889), .A2(new_n890), .A3(G148gat), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n307), .A2(new_n310), .A3(new_n340), .A4(new_n384), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT118), .B1(new_n861), .B2(new_n821), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n248), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n861), .A2(KEYINPUT118), .A3(new_n821), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n568), .A2(KEYINPUT57), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n825), .A2(new_n567), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT57), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n853), .B(KEYINPUT117), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n341), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n890), .B1(new_n904), .B2(G148gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n887), .B1(new_n891), .B2(new_n905), .ZN(G1345gat));
  OR3_X1    g705(.A1(new_n888), .A2(new_n483), .A3(new_n248), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n885), .A2(new_n249), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n483), .B2(new_n909), .ZN(G1346gat));
  OAI21_X1  g709(.A(G162gat), .B1(new_n888), .B2(new_n306), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n885), .A2(new_n484), .A3(new_n309), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1347gat));
  AOI21_X1  g712(.A(new_n666), .B1(new_n822), .B2(new_n824), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n638), .A2(new_n649), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n413), .B1(new_n916), .B2(new_n823), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n852), .A2(G169gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT119), .ZN(G1348gat));
  NOR2_X1   g719(.A1(new_n916), .A2(new_n340), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(new_n414), .ZN(G1349gat));
  INV_X1    g721(.A(new_n916), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n249), .A3(new_n407), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n925));
  OAI21_X1  g724(.A(G183gat), .B1(new_n916), .B2(new_n248), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT120), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT120), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n924), .A2(new_n931), .A3(new_n926), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n930), .B1(new_n933), .B2(new_n929), .ZN(G1350gat));
  NAND2_X1  g733(.A1(new_n923), .A2(new_n309), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n935), .A2(G190gat), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n936), .A2(KEYINPUT122), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(KEYINPUT122), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(G190gat), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n939), .A2(KEYINPUT61), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n939), .A2(KEYINPUT61), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n937), .A2(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1351gat));
  NAND3_X1  g741(.A1(new_n657), .A2(new_n649), .A3(new_n567), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT123), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n944), .A2(new_n914), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n370), .A3(new_n691), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n657), .A2(new_n645), .A3(new_n649), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT124), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n902), .A2(new_n852), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n946), .B1(new_n949), .B2(new_n370), .ZN(G1352gat));
  INV_X1    g749(.A(G204gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n945), .A2(new_n951), .A3(new_n341), .ZN(new_n952));
  XOR2_X1   g751(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n953));
  XNOR2_X1  g752(.A(new_n952), .B(new_n953), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n902), .A2(new_n341), .A3(new_n948), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n951), .B2(new_n955), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n945), .A2(new_n390), .A3(new_n249), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n899), .A2(new_n249), .A3(new_n901), .A4(new_n948), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G211gat), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT63), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(KEYINPUT126), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT126), .B1(new_n959), .B2(new_n960), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n957), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  NAND3_X1  g764(.A1(new_n902), .A2(KEYINPUT127), .A3(new_n948), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(new_n309), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT127), .B1(new_n902), .B2(new_n948), .ZN(new_n968));
  OAI21_X1  g767(.A(G218gat), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n945), .A2(new_n391), .A3(new_n309), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1355gat));
endmodule


