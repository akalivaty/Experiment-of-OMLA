

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X4 U558 ( .A(n673), .Z(n523) );
  XNOR2_X1 U559 ( .A(n543), .B(n542), .ZN(n673) );
  NOR2_X1 U560 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U561 ( .A1(G651), .A2(G543), .ZN(n796) );
  OR2_X1 U562 ( .A1(n950), .A2(n619), .ZN(n618) );
  NOR2_X1 U563 ( .A1(G168), .A2(n646), .ZN(n647) );
  NAND2_X1 U564 ( .A1(n591), .A2(n685), .ZN(n664) );
  XNOR2_X1 U565 ( .A(n654), .B(KEYINPUT92), .ZN(n662) );
  XNOR2_X1 U566 ( .A(G543), .B(KEYINPUT0), .ZN(n524) );
  NOR2_X1 U567 ( .A1(G164), .A2(G1384), .ZN(n685) );
  XNOR2_X1 U568 ( .A(n524), .B(KEYINPUT67), .ZN(n585) );
  NOR2_X1 U569 ( .A1(G651), .A2(n585), .ZN(n793) );
  NOR2_X1 U570 ( .A1(G2104), .A2(n541), .ZN(n884) );
  XNOR2_X1 U571 ( .A(KEYINPUT75), .B(n601), .ZN(n950) );
  INV_X1 U572 ( .A(G651), .ZN(n531) );
  NOR2_X1 U573 ( .A1(n531), .A2(n585), .ZN(n525) );
  XNOR2_X2 U574 ( .A(KEYINPUT68), .B(n525), .ZN(n797) );
  NAND2_X1 U575 ( .A1(G76), .A2(n797), .ZN(n526) );
  XNOR2_X1 U576 ( .A(KEYINPUT76), .B(n526), .ZN(n529) );
  NAND2_X1 U577 ( .A1(n796), .A2(G89), .ZN(n527) );
  XNOR2_X1 U578 ( .A(KEYINPUT4), .B(n527), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U580 ( .A(n530), .B(KEYINPUT5), .ZN(n537) );
  NOR2_X1 U581 ( .A1(G543), .A2(n531), .ZN(n532) );
  XOR2_X1 U582 ( .A(KEYINPUT1), .B(n532), .Z(n792) );
  NAND2_X1 U583 ( .A1(G63), .A2(n792), .ZN(n534) );
  NAND2_X1 U584 ( .A1(G51), .A2(n793), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U586 ( .A(KEYINPUT6), .B(n535), .Z(n536) );
  NAND2_X1 U587 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U588 ( .A(n538), .B(KEYINPUT7), .ZN(G168) );
  INV_X1 U589 ( .A(G2105), .ZN(n541) );
  AND2_X1 U590 ( .A1(n541), .A2(G2104), .ZN(n881) );
  NAND2_X1 U591 ( .A1(G102), .A2(n881), .ZN(n540) );
  AND2_X1 U592 ( .A1(G2104), .A2(G2105), .ZN(n885) );
  NAND2_X1 U593 ( .A1(G114), .A2(n885), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n547) );
  NAND2_X1 U595 ( .A1(G126), .A2(n884), .ZN(n545) );
  XNOR2_X1 U596 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n543) );
  NOR2_X1 U597 ( .A1(G2104), .A2(G2105), .ZN(n542) );
  NAND2_X1 U598 ( .A1(G138), .A2(n523), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U600 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U601 ( .A(n548), .B(KEYINPUT84), .ZN(G164) );
  NAND2_X1 U602 ( .A1(G125), .A2(n884), .ZN(n550) );
  NAND2_X1 U603 ( .A1(G113), .A2(n885), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n557) );
  NAND2_X1 U605 ( .A1(n523), .A2(G137), .ZN(n551) );
  XNOR2_X1 U606 ( .A(n551), .B(KEYINPUT66), .ZN(n555) );
  XOR2_X1 U607 ( .A(KEYINPUT23), .B(KEYINPUT64), .Z(n553) );
  NAND2_X1 U608 ( .A1(G101), .A2(n881), .ZN(n552) );
  XNOR2_X1 U609 ( .A(n553), .B(n552), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U611 ( .A1(n557), .A2(n556), .ZN(G160) );
  NAND2_X1 U612 ( .A1(G64), .A2(n792), .ZN(n559) );
  NAND2_X1 U613 ( .A1(G52), .A2(n793), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n559), .A2(n558), .ZN(n564) );
  NAND2_X1 U615 ( .A1(G90), .A2(n796), .ZN(n561) );
  NAND2_X1 U616 ( .A1(G77), .A2(n797), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U618 ( .A(KEYINPUT9), .B(n562), .Z(n563) );
  NOR2_X1 U619 ( .A1(n564), .A2(n563), .ZN(G171) );
  INV_X1 U620 ( .A(G171), .ZN(G301) );
  XOR2_X1 U621 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U622 ( .A1(G88), .A2(n796), .ZN(n566) );
  NAND2_X1 U623 ( .A1(G75), .A2(n797), .ZN(n565) );
  NAND2_X1 U624 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U625 ( .A1(G62), .A2(n792), .ZN(n568) );
  NAND2_X1 U626 ( .A1(G50), .A2(n793), .ZN(n567) );
  NAND2_X1 U627 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U628 ( .A1(n570), .A2(n569), .ZN(G166) );
  INV_X1 U629 ( .A(G166), .ZN(G303) );
  AND2_X1 U630 ( .A1(n792), .A2(G60), .ZN(n574) );
  NAND2_X1 U631 ( .A1(G85), .A2(n796), .ZN(n572) );
  NAND2_X1 U632 ( .A1(G47), .A2(n793), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U634 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U635 ( .A1(G72), .A2(n797), .ZN(n575) );
  NAND2_X1 U636 ( .A1(n576), .A2(n575), .ZN(G290) );
  NAND2_X1 U637 ( .A1(n797), .A2(G73), .ZN(n577) );
  XNOR2_X1 U638 ( .A(n577), .B(KEYINPUT2), .ZN(n584) );
  NAND2_X1 U639 ( .A1(G86), .A2(n796), .ZN(n579) );
  NAND2_X1 U640 ( .A1(G48), .A2(n793), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U642 ( .A1(G61), .A2(n792), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT81), .B(n580), .ZN(n581) );
  NOR2_X1 U644 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n584), .A2(n583), .ZN(G305) );
  NAND2_X1 U646 ( .A1(G49), .A2(n793), .ZN(n587) );
  NAND2_X1 U647 ( .A1(G87), .A2(n585), .ZN(n586) );
  NAND2_X1 U648 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U649 ( .A1(n792), .A2(n588), .ZN(n590) );
  NAND2_X1 U650 ( .A1(G651), .A2(G74), .ZN(n589) );
  NAND2_X1 U651 ( .A1(n590), .A2(n589), .ZN(G288) );
  NAND2_X1 U652 ( .A1(G160), .A2(G40), .ZN(n684) );
  INV_X1 U653 ( .A(n684), .ZN(n591) );
  NAND2_X1 U654 ( .A1(G8), .A2(n664), .ZN(n721) );
  NOR2_X1 U655 ( .A1(G1966), .A2(n721), .ZN(n655) );
  NAND2_X1 U656 ( .A1(G79), .A2(n797), .ZN(n592) );
  XOR2_X1 U657 ( .A(n592), .B(KEYINPUT73), .Z(n594) );
  NAND2_X1 U658 ( .A1(n793), .A2(G54), .ZN(n593) );
  NAND2_X1 U659 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U660 ( .A(KEYINPUT74), .B(n595), .ZN(n599) );
  NAND2_X1 U661 ( .A1(G66), .A2(n792), .ZN(n597) );
  NAND2_X1 U662 ( .A1(G92), .A2(n796), .ZN(n596) );
  NAND2_X1 U663 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U664 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U665 ( .A(n600), .B(KEYINPUT15), .Z(n601) );
  NAND2_X1 U666 ( .A1(G1348), .A2(n664), .ZN(n603) );
  INV_X1 U667 ( .A(n664), .ZN(n639) );
  NAND2_X1 U668 ( .A1(G2067), .A2(n639), .ZN(n602) );
  NAND2_X1 U669 ( .A1(n603), .A2(n602), .ZN(n619) );
  NAND2_X1 U670 ( .A1(G56), .A2(n792), .ZN(n604) );
  XOR2_X1 U671 ( .A(KEYINPUT14), .B(n604), .Z(n610) );
  NAND2_X1 U672 ( .A1(n796), .A2(G81), .ZN(n605) );
  XNOR2_X1 U673 ( .A(n605), .B(KEYINPUT12), .ZN(n607) );
  NAND2_X1 U674 ( .A1(G68), .A2(n797), .ZN(n606) );
  NAND2_X1 U675 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U676 ( .A(KEYINPUT13), .B(n608), .Z(n609) );
  NOR2_X1 U677 ( .A1(n610), .A2(n609), .ZN(n612) );
  NAND2_X1 U678 ( .A1(n793), .A2(G43), .ZN(n611) );
  NAND2_X1 U679 ( .A1(n612), .A2(n611), .ZN(n955) );
  AND2_X1 U680 ( .A1(n639), .A2(G1996), .ZN(n613) );
  XOR2_X1 U681 ( .A(n613), .B(KEYINPUT26), .Z(n615) );
  NAND2_X1 U682 ( .A1(n664), .A2(G1341), .ZN(n614) );
  NAND2_X1 U683 ( .A1(n615), .A2(n614), .ZN(n616) );
  OR2_X1 U684 ( .A1(n955), .A2(n616), .ZN(n617) );
  NAND2_X1 U685 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U686 ( .A1(n950), .A2(n619), .ZN(n620) );
  NAND2_X1 U687 ( .A1(n621), .A2(n620), .ZN(n633) );
  NAND2_X1 U688 ( .A1(G65), .A2(n792), .ZN(n623) );
  NAND2_X1 U689 ( .A1(G53), .A2(n793), .ZN(n622) );
  NAND2_X1 U690 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U691 ( .A1(G91), .A2(n796), .ZN(n625) );
  NAND2_X1 U692 ( .A1(G78), .A2(n797), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U694 ( .A1(n627), .A2(n626), .ZN(n961) );
  NAND2_X1 U695 ( .A1(n639), .A2(G2072), .ZN(n628) );
  XNOR2_X1 U696 ( .A(n628), .B(KEYINPUT27), .ZN(n630) );
  XNOR2_X1 U697 ( .A(G1956), .B(KEYINPUT89), .ZN(n928) );
  NOR2_X1 U698 ( .A1(n928), .A2(n639), .ZN(n629) );
  NOR2_X1 U699 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U700 ( .A(KEYINPUT90), .B(n631), .ZN(n634) );
  NAND2_X1 U701 ( .A1(n961), .A2(n634), .ZN(n632) );
  NAND2_X1 U702 ( .A1(n633), .A2(n632), .ZN(n637) );
  NOR2_X1 U703 ( .A1(n961), .A2(n634), .ZN(n635) );
  XOR2_X1 U704 ( .A(n635), .B(KEYINPUT28), .Z(n636) );
  NAND2_X1 U705 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U706 ( .A(n638), .B(KEYINPUT29), .ZN(n643) );
  XOR2_X1 U707 ( .A(KEYINPUT25), .B(G2078), .Z(n976) );
  NOR2_X1 U708 ( .A1(n976), .A2(n664), .ZN(n641) );
  NOR2_X1 U709 ( .A1(n639), .A2(G1961), .ZN(n640) );
  NOR2_X1 U710 ( .A1(n641), .A2(n640), .ZN(n648) );
  NOR2_X1 U711 ( .A1(G301), .A2(n648), .ZN(n642) );
  NOR2_X1 U712 ( .A1(n643), .A2(n642), .ZN(n653) );
  NOR2_X1 U713 ( .A1(G2084), .A2(n664), .ZN(n657) );
  NOR2_X1 U714 ( .A1(n657), .A2(n655), .ZN(n644) );
  NAND2_X1 U715 ( .A1(G8), .A2(n644), .ZN(n645) );
  XNOR2_X1 U716 ( .A(KEYINPUT30), .B(n645), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n647), .B(KEYINPUT91), .ZN(n650) );
  NAND2_X1 U718 ( .A1(n648), .A2(G301), .ZN(n649) );
  NAND2_X1 U719 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U720 ( .A(KEYINPUT31), .B(n651), .Z(n652) );
  NOR2_X1 U721 ( .A1(n655), .A2(n662), .ZN(n656) );
  XNOR2_X1 U722 ( .A(KEYINPUT93), .B(n656), .ZN(n659) );
  AND2_X1 U723 ( .A1(G8), .A2(n657), .ZN(n658) );
  NOR2_X1 U724 ( .A1(n659), .A2(n658), .ZN(n661) );
  INV_X1 U725 ( .A(KEYINPUT94), .ZN(n660) );
  XNOR2_X1 U726 ( .A(n661), .B(n660), .ZN(n733) );
  INV_X1 U727 ( .A(n662), .ZN(n663) );
  NAND2_X1 U728 ( .A1(G286), .A2(n663), .ZN(n670) );
  NOR2_X1 U729 ( .A1(G1971), .A2(n721), .ZN(n666) );
  NOR2_X1 U730 ( .A1(G2090), .A2(n664), .ZN(n665) );
  NOR2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U732 ( .A1(n667), .A2(G303), .ZN(n668) );
  XOR2_X1 U733 ( .A(KEYINPUT95), .B(n668), .Z(n669) );
  NAND2_X1 U734 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U735 ( .A1(n671), .A2(G8), .ZN(n672) );
  XNOR2_X1 U736 ( .A(n672), .B(KEYINPUT32), .ZN(n731) );
  XNOR2_X1 U737 ( .A(G2067), .B(KEYINPUT37), .ZN(n756) );
  XNOR2_X1 U738 ( .A(KEYINPUT86), .B(KEYINPUT34), .ZN(n677) );
  NAND2_X1 U739 ( .A1(G104), .A2(n881), .ZN(n675) );
  NAND2_X1 U740 ( .A1(G140), .A2(n523), .ZN(n674) );
  NAND2_X1 U741 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U742 ( .A(n677), .B(n676), .ZN(n682) );
  NAND2_X1 U743 ( .A1(G128), .A2(n884), .ZN(n679) );
  NAND2_X1 U744 ( .A1(G116), .A2(n885), .ZN(n678) );
  NAND2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U746 ( .A(KEYINPUT35), .B(n680), .Z(n681) );
  NOR2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U748 ( .A(KEYINPUT36), .B(n683), .ZN(n898) );
  NOR2_X1 U749 ( .A1(n756), .A2(n898), .ZN(n1014) );
  NOR2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n759) );
  NAND2_X1 U751 ( .A1(n1014), .A2(n759), .ZN(n686) );
  XNOR2_X1 U752 ( .A(n686), .B(KEYINPUT87), .ZN(n753) );
  XNOR2_X1 U753 ( .A(G1986), .B(G290), .ZN(n957) );
  NAND2_X1 U754 ( .A1(n759), .A2(n957), .ZN(n687) );
  XNOR2_X1 U755 ( .A(KEYINPUT85), .B(n687), .ZN(n688) );
  NOR2_X1 U756 ( .A1(n753), .A2(n688), .ZN(n705) );
  NAND2_X1 U757 ( .A1(G119), .A2(n884), .ZN(n690) );
  NAND2_X1 U758 ( .A1(G131), .A2(n523), .ZN(n689) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n694) );
  NAND2_X1 U760 ( .A1(G95), .A2(n881), .ZN(n692) );
  NAND2_X1 U761 ( .A1(G107), .A2(n885), .ZN(n691) );
  NAND2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n693) );
  OR2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n876) );
  NAND2_X1 U764 ( .A1(G1991), .A2(n876), .ZN(n704) );
  XOR2_X1 U765 ( .A(KEYINPUT88), .B(KEYINPUT38), .Z(n696) );
  NAND2_X1 U766 ( .A1(G105), .A2(n881), .ZN(n695) );
  XNOR2_X1 U767 ( .A(n696), .B(n695), .ZN(n700) );
  NAND2_X1 U768 ( .A1(G129), .A2(n884), .ZN(n698) );
  NAND2_X1 U769 ( .A1(G141), .A2(n523), .ZN(n697) );
  NAND2_X1 U770 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U771 ( .A1(n700), .A2(n699), .ZN(n702) );
  NAND2_X1 U772 ( .A1(n885), .A2(G117), .ZN(n701) );
  NAND2_X1 U773 ( .A1(n702), .A2(n701), .ZN(n892) );
  NAND2_X1 U774 ( .A1(G1996), .A2(n892), .ZN(n703) );
  NAND2_X1 U775 ( .A1(n704), .A2(n703), .ZN(n1008) );
  NAND2_X1 U776 ( .A1(n759), .A2(n1008), .ZN(n745) );
  NAND2_X1 U777 ( .A1(n705), .A2(n745), .ZN(n726) );
  NOR2_X1 U778 ( .A1(G1981), .A2(G305), .ZN(n706) );
  XOR2_X1 U779 ( .A(n706), .B(KEYINPUT24), .Z(n707) );
  NOR2_X1 U780 ( .A1(n721), .A2(n707), .ZN(n712) );
  NOR2_X1 U781 ( .A1(n712), .A2(n721), .ZN(n708) );
  NOR2_X1 U782 ( .A1(n726), .A2(n708), .ZN(n710) );
  AND2_X1 U783 ( .A1(n731), .A2(n710), .ZN(n709) );
  NAND2_X1 U784 ( .A1(n733), .A2(n709), .ZN(n718) );
  INV_X1 U785 ( .A(n710), .ZN(n716) );
  NOR2_X1 U786 ( .A1(G2090), .A2(G303), .ZN(n711) );
  NAND2_X1 U787 ( .A1(G8), .A2(n711), .ZN(n714) );
  INV_X1 U788 ( .A(n712), .ZN(n713) );
  AND2_X1 U789 ( .A1(n714), .A2(n713), .ZN(n715) );
  OR2_X1 U790 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U791 ( .A1(n718), .A2(n717), .ZN(n743) );
  NAND2_X1 U792 ( .A1(G1976), .A2(G288), .ZN(n959) );
  INV_X1 U793 ( .A(n959), .ZN(n719) );
  NOR2_X1 U794 ( .A1(n719), .A2(n721), .ZN(n720) );
  OR2_X1 U795 ( .A1(KEYINPUT33), .A2(n720), .ZN(n730) );
  NOR2_X1 U796 ( .A1(G1976), .A2(G288), .ZN(n958) );
  NAND2_X1 U797 ( .A1(n958), .A2(KEYINPUT33), .ZN(n722) );
  NOR2_X1 U798 ( .A1(n722), .A2(n721), .ZN(n725) );
  XOR2_X1 U799 ( .A(G1981), .B(KEYINPUT96), .Z(n723) );
  XNOR2_X1 U800 ( .A(G305), .B(n723), .ZN(n947) );
  INV_X1 U801 ( .A(n947), .ZN(n724) );
  NOR2_X1 U802 ( .A1(n725), .A2(n724), .ZN(n728) );
  INV_X1 U803 ( .A(n726), .ZN(n727) );
  AND2_X1 U804 ( .A1(n728), .A2(n727), .ZN(n729) );
  AND2_X1 U805 ( .A1(n730), .A2(n729), .ZN(n734) );
  AND2_X1 U806 ( .A1(n731), .A2(n734), .ZN(n732) );
  NAND2_X1 U807 ( .A1(n733), .A2(n732), .ZN(n741) );
  INV_X1 U808 ( .A(n734), .ZN(n739) );
  NOR2_X1 U809 ( .A1(G1971), .A2(G303), .ZN(n735) );
  NOR2_X1 U810 ( .A1(n958), .A2(n735), .ZN(n737) );
  INV_X1 U811 ( .A(KEYINPUT33), .ZN(n736) );
  AND2_X1 U812 ( .A1(n737), .A2(n736), .ZN(n738) );
  OR2_X1 U813 ( .A1(n739), .A2(n738), .ZN(n740) );
  AND2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U815 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U816 ( .A(n744), .B(KEYINPUT97), .ZN(n761) );
  NOR2_X1 U817 ( .A1(G1996), .A2(n892), .ZN(n998) );
  INV_X1 U818 ( .A(n745), .ZN(n749) );
  NOR2_X1 U819 ( .A1(G1986), .A2(G290), .ZN(n747) );
  NOR2_X1 U820 ( .A1(G1991), .A2(n876), .ZN(n746) );
  XNOR2_X1 U821 ( .A(KEYINPUT98), .B(n746), .ZN(n1011) );
  NOR2_X1 U822 ( .A1(n747), .A2(n1011), .ZN(n748) );
  NOR2_X1 U823 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U824 ( .A(KEYINPUT99), .B(n750), .Z(n751) );
  NOR2_X1 U825 ( .A1(n998), .A2(n751), .ZN(n752) );
  XNOR2_X1 U826 ( .A(KEYINPUT39), .B(n752), .ZN(n755) );
  INV_X1 U827 ( .A(n753), .ZN(n754) );
  NAND2_X1 U828 ( .A1(n755), .A2(n754), .ZN(n757) );
  NAND2_X1 U829 ( .A1(n756), .A2(n898), .ZN(n1000) );
  NAND2_X1 U830 ( .A1(n757), .A2(n1000), .ZN(n758) );
  NAND2_X1 U831 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U832 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U833 ( .A(n762), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U834 ( .A(G120), .ZN(G236) );
  INV_X1 U835 ( .A(G82), .ZN(G220) );
  NAND2_X1 U836 ( .A1(G94), .A2(G452), .ZN(n763) );
  XNOR2_X1 U837 ( .A(n763), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U838 ( .A1(G7), .A2(G661), .ZN(n764) );
  XNOR2_X1 U839 ( .A(n764), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U840 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n766) );
  XNOR2_X1 U841 ( .A(G223), .B(KEYINPUT71), .ZN(n829) );
  NAND2_X1 U842 ( .A1(G567), .A2(n829), .ZN(n765) );
  XNOR2_X1 U843 ( .A(n766), .B(n765), .ZN(G234) );
  INV_X1 U844 ( .A(n955), .ZN(n767) );
  NAND2_X1 U845 ( .A1(n767), .A2(G860), .ZN(G153) );
  NAND2_X1 U846 ( .A1(G868), .A2(G301), .ZN(n769) );
  INV_X1 U847 ( .A(G868), .ZN(n813) );
  NAND2_X1 U848 ( .A1(n950), .A2(n813), .ZN(n768) );
  NAND2_X1 U849 ( .A1(n769), .A2(n768), .ZN(G284) );
  INV_X1 U850 ( .A(n961), .ZN(G299) );
  NOR2_X1 U851 ( .A1(G286), .A2(n813), .ZN(n771) );
  NOR2_X1 U852 ( .A1(G868), .A2(G299), .ZN(n770) );
  NOR2_X1 U853 ( .A1(n771), .A2(n770), .ZN(G297) );
  INV_X1 U854 ( .A(G559), .ZN(n772) );
  NOR2_X1 U855 ( .A1(G860), .A2(n772), .ZN(n773) );
  XNOR2_X1 U856 ( .A(KEYINPUT77), .B(n773), .ZN(n774) );
  INV_X1 U857 ( .A(n950), .ZN(n790) );
  NAND2_X1 U858 ( .A1(n774), .A2(n790), .ZN(n775) );
  XNOR2_X1 U859 ( .A(n775), .B(KEYINPUT16), .ZN(n776) );
  XNOR2_X1 U860 ( .A(KEYINPUT78), .B(n776), .ZN(G148) );
  NOR2_X1 U861 ( .A1(G559), .A2(n813), .ZN(n777) );
  NAND2_X1 U862 ( .A1(n790), .A2(n777), .ZN(n778) );
  XNOR2_X1 U863 ( .A(n778), .B(KEYINPUT79), .ZN(n780) );
  NOR2_X1 U864 ( .A1(n955), .A2(G868), .ZN(n779) );
  NOR2_X1 U865 ( .A1(n780), .A2(n779), .ZN(G282) );
  NAND2_X1 U866 ( .A1(n884), .A2(G123), .ZN(n781) );
  XNOR2_X1 U867 ( .A(n781), .B(KEYINPUT18), .ZN(n783) );
  NAND2_X1 U868 ( .A1(G111), .A2(n885), .ZN(n782) );
  NAND2_X1 U869 ( .A1(n783), .A2(n782), .ZN(n787) );
  NAND2_X1 U870 ( .A1(G99), .A2(n881), .ZN(n785) );
  NAND2_X1 U871 ( .A1(G135), .A2(n523), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n1009) );
  XOR2_X1 U874 ( .A(G2096), .B(n1009), .Z(n788) );
  NOR2_X1 U875 ( .A1(G2100), .A2(n788), .ZN(n789) );
  XOR2_X1 U876 ( .A(KEYINPUT80), .B(n789), .Z(G156) );
  NAND2_X1 U877 ( .A1(n790), .A2(G559), .ZN(n810) );
  XNOR2_X1 U878 ( .A(n955), .B(n810), .ZN(n791) );
  NOR2_X1 U879 ( .A1(n791), .A2(G860), .ZN(n802) );
  NAND2_X1 U880 ( .A1(G67), .A2(n792), .ZN(n795) );
  NAND2_X1 U881 ( .A1(G55), .A2(n793), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n801) );
  NAND2_X1 U883 ( .A1(G93), .A2(n796), .ZN(n799) );
  NAND2_X1 U884 ( .A1(G80), .A2(n797), .ZN(n798) );
  NAND2_X1 U885 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U886 ( .A1(n801), .A2(n800), .ZN(n812) );
  XNOR2_X1 U887 ( .A(n802), .B(n812), .ZN(G145) );
  XNOR2_X1 U888 ( .A(KEYINPUT19), .B(G305), .ZN(n803) );
  XNOR2_X1 U889 ( .A(n803), .B(G288), .ZN(n804) );
  XOR2_X1 U890 ( .A(n804), .B(KEYINPUT82), .Z(n806) );
  XNOR2_X1 U891 ( .A(n961), .B(n812), .ZN(n805) );
  XNOR2_X1 U892 ( .A(n806), .B(n805), .ZN(n807) );
  XNOR2_X1 U893 ( .A(G166), .B(n807), .ZN(n808) );
  XNOR2_X1 U894 ( .A(n808), .B(G290), .ZN(n809) );
  XNOR2_X1 U895 ( .A(n955), .B(n809), .ZN(n901) );
  XOR2_X1 U896 ( .A(n901), .B(n810), .Z(n811) );
  NOR2_X1 U897 ( .A1(n813), .A2(n811), .ZN(n815) );
  AND2_X1 U898 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U899 ( .A1(n815), .A2(n814), .ZN(G295) );
  NAND2_X1 U900 ( .A1(G2084), .A2(G2078), .ZN(n816) );
  XNOR2_X1 U901 ( .A(n816), .B(KEYINPUT83), .ZN(n817) );
  XNOR2_X1 U902 ( .A(n817), .B(KEYINPUT20), .ZN(n818) );
  NAND2_X1 U903 ( .A1(n818), .A2(G2090), .ZN(n819) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n819), .ZN(n820) );
  NAND2_X1 U905 ( .A1(n820), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U907 ( .A(KEYINPUT70), .B(G132), .Z(G219) );
  NOR2_X1 U908 ( .A1(G219), .A2(G220), .ZN(n821) );
  XOR2_X1 U909 ( .A(KEYINPUT22), .B(n821), .Z(n822) );
  NOR2_X1 U910 ( .A1(G218), .A2(n822), .ZN(n823) );
  NAND2_X1 U911 ( .A1(G96), .A2(n823), .ZN(n835) );
  NAND2_X1 U912 ( .A1(n835), .A2(G2106), .ZN(n827) );
  NAND2_X1 U913 ( .A1(G69), .A2(G108), .ZN(n824) );
  NOR2_X1 U914 ( .A1(G236), .A2(n824), .ZN(n825) );
  NAND2_X1 U915 ( .A1(G57), .A2(n825), .ZN(n836) );
  NAND2_X1 U916 ( .A1(n836), .A2(G567), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n827), .A2(n826), .ZN(n837) );
  NAND2_X1 U918 ( .A1(G483), .A2(G661), .ZN(n828) );
  NOR2_X1 U919 ( .A1(n837), .A2(n828), .ZN(n834) );
  NAND2_X1 U920 ( .A1(n834), .A2(G36), .ZN(G176) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n829), .ZN(G217) );
  INV_X1 U922 ( .A(G661), .ZN(n831) );
  NAND2_X1 U923 ( .A1(G2), .A2(G15), .ZN(n830) );
  NOR2_X1 U924 ( .A1(n831), .A2(n830), .ZN(n832) );
  XOR2_X1 U925 ( .A(KEYINPUT100), .B(n832), .Z(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n834), .A2(n833), .ZN(G188) );
  XNOR2_X1 U928 ( .A(G69), .B(KEYINPUT101), .ZN(G235) );
  XOR2_X1 U929 ( .A(G108), .B(KEYINPUT112), .Z(G238) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  NOR2_X1 U932 ( .A1(n836), .A2(n835), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  INV_X1 U934 ( .A(n837), .ZN(G319) );
  XOR2_X1 U935 ( .A(KEYINPUT102), .B(G2678), .Z(n839) );
  XNOR2_X1 U936 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U938 ( .A(KEYINPUT103), .B(G2090), .Z(n841) );
  XNOR2_X1 U939 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U941 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U942 ( .A(G2096), .B(G2100), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n847) );
  XOR2_X1 U944 ( .A(G2084), .B(G2078), .Z(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(G227) );
  XOR2_X1 U946 ( .A(G1976), .B(G1971), .Z(n849) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1956), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U949 ( .A(n850), .B(G2474), .Z(n852) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1981), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U952 ( .A(KEYINPUT41), .B(G1961), .Z(n854) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(G229) );
  NAND2_X1 U956 ( .A1(G136), .A2(n523), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n857), .B(KEYINPUT104), .ZN(n860) );
  NAND2_X1 U958 ( .A1(G124), .A2(n884), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n858), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n865) );
  NAND2_X1 U961 ( .A1(G100), .A2(n881), .ZN(n862) );
  NAND2_X1 U962 ( .A1(G112), .A2(n885), .ZN(n861) );
  NAND2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U964 ( .A(KEYINPUT105), .B(n863), .Z(n864) );
  NOR2_X1 U965 ( .A1(n865), .A2(n864), .ZN(G162) );
  NAND2_X1 U966 ( .A1(G106), .A2(n881), .ZN(n867) );
  NAND2_X1 U967 ( .A1(G142), .A2(n523), .ZN(n866) );
  NAND2_X1 U968 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n868), .B(KEYINPUT45), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G130), .A2(n884), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G118), .A2(n885), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U973 ( .A(KEYINPUT106), .B(n871), .Z(n872) );
  NAND2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n874), .B(G164), .ZN(n897) );
  XOR2_X1 U976 ( .A(KEYINPUT109), .B(KEYINPUT46), .Z(n875) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U978 ( .A(n877), .B(KEYINPUT107), .Z(n879) );
  XNOR2_X1 U979 ( .A(G160), .B(KEYINPUT48), .ZN(n878) );
  XNOR2_X1 U980 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n1009), .B(n880), .ZN(n894) );
  NAND2_X1 U982 ( .A1(G103), .A2(n881), .ZN(n883) );
  NAND2_X1 U983 ( .A1(G139), .A2(n523), .ZN(n882) );
  NAND2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n890) );
  NAND2_X1 U985 ( .A1(G127), .A2(n884), .ZN(n887) );
  NAND2_X1 U986 ( .A1(G115), .A2(n885), .ZN(n886) );
  NAND2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U989 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U990 ( .A(KEYINPUT108), .B(n891), .Z(n1002) );
  XNOR2_X1 U991 ( .A(n892), .B(n1002), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U993 ( .A(G162), .B(n895), .Z(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n899) );
  XOR2_X1 U995 ( .A(n899), .B(n898), .Z(n900) );
  NOR2_X1 U996 ( .A1(G37), .A2(n900), .ZN(G395) );
  XNOR2_X1 U997 ( .A(G286), .B(n950), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n904) );
  XOR2_X1 U999 ( .A(G171), .B(KEYINPUT110), .Z(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n905), .ZN(G397) );
  XOR2_X1 U1002 ( .A(G2451), .B(G2430), .Z(n907) );
  XNOR2_X1 U1003 ( .A(G2438), .B(G2443), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n913) );
  XOR2_X1 U1005 ( .A(G2435), .B(G2454), .Z(n909) );
  XNOR2_X1 U1006 ( .A(G1341), .B(G1348), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n911) );
  XOR2_X1 U1008 ( .A(G2446), .B(G2427), .Z(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1010 ( .A(n913), .B(n912), .Z(n914) );
  NAND2_X1 U1011 ( .A1(G14), .A2(n914), .ZN(n921) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n921), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n915) );
  XOR2_X1 U1014 ( .A(KEYINPUT111), .B(n915), .Z(n916) );
  XNOR2_X1 U1015 ( .A(n916), .B(KEYINPUT49), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G57), .ZN(G237) );
  INV_X1 U1021 ( .A(n921), .ZN(G401) );
  XNOR2_X1 U1022 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n1031) );
  XNOR2_X1 U1023 ( .A(G1971), .B(G22), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(G1976), .B(G23), .ZN(n922) );
  NOR2_X1 U1025 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1026 ( .A(KEYINPUT124), .B(n924), .Z(n926) );
  XNOR2_X1 U1027 ( .A(G1986), .B(G24), .ZN(n925) );
  NOR2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1029 ( .A(KEYINPUT58), .B(n927), .ZN(n943) );
  XNOR2_X1 U1030 ( .A(G1961), .B(G5), .ZN(n941) );
  XNOR2_X1 U1031 ( .A(G20), .B(n928), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(G1341), .B(G19), .ZN(n930) );
  XNOR2_X1 U1033 ( .A(G1981), .B(G6), .ZN(n929) );
  NOR2_X1 U1034 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1035 ( .A1(n932), .A2(n931), .ZN(n935) );
  XOR2_X1 U1036 ( .A(KEYINPUT59), .B(G1348), .Z(n933) );
  XNOR2_X1 U1037 ( .A(G4), .B(n933), .ZN(n934) );
  NOR2_X1 U1038 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1039 ( .A(KEYINPUT60), .B(n936), .Z(n938) );
  XNOR2_X1 U1040 ( .A(G1966), .B(G21), .ZN(n937) );
  NOR2_X1 U1041 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1042 ( .A(KEYINPUT123), .B(n939), .ZN(n940) );
  NOR2_X1 U1043 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1045 ( .A(n944), .B(KEYINPUT61), .ZN(n945) );
  XOR2_X1 U1046 ( .A(KEYINPUT125), .B(n945), .Z(n946) );
  NOR2_X1 U1047 ( .A1(G16), .A2(n946), .ZN(n1029) );
  XOR2_X1 U1048 ( .A(KEYINPUT56), .B(G16), .Z(n973) );
  XNOR2_X1 U1049 ( .A(G1966), .B(G168), .ZN(n948) );
  NAND2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1051 ( .A(n949), .B(KEYINPUT57), .ZN(n954) );
  XNOR2_X1 U1052 ( .A(G301), .B(G1961), .ZN(n952) );
  XNOR2_X1 U1053 ( .A(n950), .B(G1348), .ZN(n951) );
  NOR2_X1 U1054 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1055 ( .A1(n954), .A2(n953), .ZN(n971) );
  XNOR2_X1 U1056 ( .A(G1341), .B(n955), .ZN(n956) );
  NOR2_X1 U1057 ( .A1(n957), .A2(n956), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(KEYINPUT121), .B(n958), .ZN(n960) );
  NAND2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(n961), .B(G1956), .ZN(n962) );
  XNOR2_X1 U1061 ( .A(n962), .B(KEYINPUT120), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(G166), .B(G1971), .ZN(n963) );
  XNOR2_X1 U1063 ( .A(n963), .B(KEYINPUT122), .ZN(n964) );
  NAND2_X1 U1064 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n1026) );
  XNOR2_X1 U1069 ( .A(KEYINPUT54), .B(G34), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(n974), .B(KEYINPUT117), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(G2084), .B(n975), .ZN(n992) );
  XNOR2_X1 U1072 ( .A(G2090), .B(G35), .ZN(n990) );
  XNOR2_X1 U1073 ( .A(G1996), .B(G32), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(n976), .B(G27), .ZN(n977) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1076 ( .A(KEYINPUT116), .B(n979), .ZN(n985) );
  XOR2_X1 U1077 ( .A(G2072), .B(G33), .Z(n980) );
  NAND2_X1 U1078 ( .A1(n980), .A2(G28), .ZN(n983) );
  XOR2_X1 U1079 ( .A(G25), .B(G1991), .Z(n981) );
  XNOR2_X1 U1080 ( .A(KEYINPUT115), .B(n981), .ZN(n982) );
  NOR2_X1 U1081 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1082 ( .A1(n985), .A2(n984), .ZN(n987) );
  XNOR2_X1 U1083 ( .A(G26), .B(G2067), .ZN(n986) );
  NOR2_X1 U1084 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1085 ( .A(KEYINPUT53), .B(n988), .ZN(n989) );
  NOR2_X1 U1086 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1088 ( .A(n993), .B(KEYINPUT55), .ZN(n994) );
  XNOR2_X1 U1089 ( .A(KEYINPUT118), .B(n994), .ZN(n995) );
  NOR2_X1 U1090 ( .A1(G29), .A2(n995), .ZN(n996) );
  XNOR2_X1 U1091 ( .A(n996), .B(KEYINPUT119), .ZN(n1024) );
  XOR2_X1 U1092 ( .A(G2090), .B(G162), .Z(n997) );
  NOR2_X1 U1093 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1094 ( .A(KEYINPUT51), .B(n999), .Z(n1001) );
  NAND2_X1 U1095 ( .A1(n1001), .A2(n1000), .ZN(n1007) );
  XOR2_X1 U1096 ( .A(G164), .B(G2078), .Z(n1004) );
  XNOR2_X1 U1097 ( .A(G2072), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1098 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1099 ( .A(KEYINPUT50), .B(n1005), .Z(n1006) );
  NOR2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1017) );
  NOR2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1013) );
  XOR2_X1 U1102 ( .A(G160), .B(G2084), .Z(n1010) );
  NOR2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(KEYINPUT52), .B(n1018), .ZN(n1019) );
  XOR2_X1 U1108 ( .A(KEYINPUT113), .B(n1019), .Z(n1020) );
  NOR2_X1 U1109 ( .A1(KEYINPUT55), .A2(n1020), .ZN(n1021) );
  XOR2_X1 U1110 ( .A(KEYINPUT114), .B(n1021), .Z(n1022) );
  NAND2_X1 U1111 ( .A1(G29), .A2(n1022), .ZN(n1023) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(G11), .ZN(n1028) );
  NOR2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1116 ( .A(n1031), .B(n1030), .ZN(n1032) );
  XNOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1032), .ZN(G150) );
  INV_X1 U1118 ( .A(G150), .ZN(G311) );
endmodule

