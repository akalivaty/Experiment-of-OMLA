

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579;

  XNOR2_X1 U322 ( .A(n325), .B(n324), .ZN(n567) );
  XOR2_X1 U323 ( .A(n380), .B(n379), .Z(n290) );
  XOR2_X1 U324 ( .A(G211GAT), .B(KEYINPUT21), .Z(n291) );
  XOR2_X1 U325 ( .A(G92GAT), .B(G64GAT), .Z(n292) );
  XNOR2_X1 U326 ( .A(n423), .B(n314), .ZN(n315) );
  XNOR2_X1 U327 ( .A(n388), .B(n315), .ZN(n316) );
  NOR2_X1 U328 ( .A1(n517), .A2(n537), .ZN(n522) );
  NOR2_X1 U329 ( .A1(n462), .A2(n510), .ZN(n557) );
  NOR2_X1 U330 ( .A1(n441), .A2(n571), .ZN(n442) );
  NOR2_X1 U331 ( .A1(n466), .A2(n524), .ZN(n468) );
  XNOR2_X1 U332 ( .A(n468), .B(n467), .ZN(n555) );
  XOR2_X1 U333 ( .A(KEYINPUT41), .B(n567), .Z(n552) );
  XOR2_X1 U334 ( .A(n387), .B(n311), .Z(n515) );
  XNOR2_X1 U335 ( .A(KEYINPUT38), .B(n443), .ZN(n495) );
  XNOR2_X1 U336 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U337 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U338 ( .A(n472), .B(n471), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(n447), .B(n446), .ZN(G1330GAT) );
  XNOR2_X1 U340 ( .A(KEYINPUT83), .B(KEYINPUT84), .ZN(n293) );
  XNOR2_X1 U341 ( .A(n293), .B(G183GAT), .ZN(n294) );
  XOR2_X1 U342 ( .A(n294), .B(KEYINPUT19), .Z(n296) );
  XNOR2_X1 U343 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n387) );
  XOR2_X1 U345 ( .A(KEYINPUT85), .B(G176GAT), .Z(n298) );
  XNOR2_X1 U346 ( .A(G190GAT), .B(G99GAT), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U348 ( .A(G15GAT), .B(G127GAT), .Z(n422) );
  XOR2_X1 U349 ( .A(n299), .B(n422), .Z(n301) );
  XNOR2_X1 U350 ( .A(G169GAT), .B(G43GAT), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U352 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n303) );
  NAND2_X1 U353 ( .A1(G227GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U355 ( .A(n305), .B(n304), .Z(n310) );
  XOR2_X1 U356 ( .A(KEYINPUT81), .B(G134GAT), .Z(n307) );
  XNOR2_X1 U357 ( .A(KEYINPUT80), .B(KEYINPUT0), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U359 ( .A(G113GAT), .B(n308), .Z(n393) );
  XOR2_X1 U360 ( .A(G120GAT), .B(G71GAT), .Z(n318) );
  XNOR2_X1 U361 ( .A(n393), .B(n318), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U363 ( .A(G176GAT), .B(KEYINPUT69), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n292), .B(n312), .ZN(n313) );
  XNOR2_X1 U365 ( .A(G204GAT), .B(n313), .ZN(n388) );
  XOR2_X1 U366 ( .A(KEYINPUT13), .B(G57GAT), .Z(n423) );
  XNOR2_X1 U367 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n314) );
  XOR2_X1 U368 ( .A(G99GAT), .B(G85GAT), .Z(n347) );
  XOR2_X1 U369 ( .A(n316), .B(n347), .Z(n320) );
  XNOR2_X1 U370 ( .A(G106GAT), .B(G78GAT), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n317), .B(G148GAT), .ZN(n371) );
  XNOR2_X1 U372 ( .A(n318), .B(n371), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n320), .B(n319), .ZN(n325) );
  XOR2_X1 U374 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n322) );
  NAND2_X1 U375 ( .A1(G230GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U377 ( .A(KEYINPUT33), .B(n323), .ZN(n324) );
  XOR2_X1 U378 ( .A(G15GAT), .B(G113GAT), .Z(n327) );
  XOR2_X1 U379 ( .A(G141GAT), .B(G22GAT), .Z(n374) );
  XOR2_X1 U380 ( .A(G169GAT), .B(G8GAT), .Z(n379) );
  XNOR2_X1 U381 ( .A(n374), .B(n379), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U383 ( .A(n328), .B(G50GAT), .Z(n333) );
  XOR2_X1 U384 ( .A(KEYINPUT68), .B(KEYINPUT65), .Z(n330) );
  XNOR2_X1 U385 ( .A(G197GAT), .B(G1GAT), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n331), .B(G36GAT), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U389 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n335) );
  NAND2_X1 U390 ( .A1(G229GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U392 ( .A(n337), .B(n336), .Z(n342) );
  XOR2_X1 U393 ( .A(KEYINPUT8), .B(KEYINPUT67), .Z(n339) );
  XNOR2_X1 U394 ( .A(G43GAT), .B(G29GAT), .ZN(n338) );
  XNOR2_X1 U395 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U396 ( .A(KEYINPUT7), .B(n340), .Z(n351) );
  XNOR2_X1 U397 ( .A(n351), .B(KEYINPUT66), .ZN(n341) );
  XOR2_X1 U398 ( .A(n342), .B(n341), .Z(n497) );
  OR2_X1 U399 ( .A1(n567), .A2(n497), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n343), .B(KEYINPUT72), .ZN(n478) );
  XOR2_X1 U401 ( .A(KEYINPUT74), .B(KEYINPUT10), .Z(n345) );
  XNOR2_X1 U402 ( .A(G134GAT), .B(KEYINPUT64), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n360) );
  XNOR2_X1 U404 ( .A(G36GAT), .B(G190GAT), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n346), .B(KEYINPUT75), .ZN(n383) );
  XOR2_X1 U406 ( .A(n347), .B(n383), .Z(n349) );
  NAND2_X1 U407 ( .A1(G232GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n358) );
  XOR2_X1 U410 ( .A(KEYINPUT73), .B(KEYINPUT9), .Z(n353) );
  XNOR2_X1 U411 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U413 ( .A(n354), .B(G106GAT), .Z(n356) );
  XOR2_X1 U414 ( .A(G50GAT), .B(G162GAT), .Z(n373) );
  XNOR2_X1 U415 ( .A(G218GAT), .B(n373), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U418 ( .A(n360), .B(n359), .Z(n545) );
  INV_X1 U419 ( .A(n545), .ZN(n473) );
  XOR2_X1 U420 ( .A(KEYINPUT36), .B(n473), .Z(n574) );
  XOR2_X1 U421 ( .A(G204GAT), .B(KEYINPUT86), .Z(n362) );
  XNOR2_X1 U422 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n362), .B(n361), .ZN(n378) );
  XOR2_X1 U424 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n364) );
  NAND2_X1 U425 ( .A1(G228GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U427 ( .A(n365), .B(KEYINPUT89), .Z(n370) );
  XNOR2_X1 U428 ( .A(G197GAT), .B(G218GAT), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n291), .B(n366), .ZN(n380) );
  XOR2_X1 U430 ( .A(G155GAT), .B(KEYINPUT2), .Z(n368) );
  XNOR2_X1 U431 ( .A(KEYINPUT3), .B(KEYINPUT88), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n392) );
  XNOR2_X1 U433 ( .A(n380), .B(n392), .ZN(n369) );
  XNOR2_X1 U434 ( .A(n370), .B(n369), .ZN(n372) );
  XOR2_X1 U435 ( .A(n372), .B(n371), .Z(n376) );
  XNOR2_X1 U436 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U437 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U438 ( .A(n378), .B(n377), .Z(n463) );
  XOR2_X1 U439 ( .A(n463), .B(KEYINPUT28), .Z(n517) );
  NAND2_X1 U440 ( .A1(G226GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n290), .B(n381), .ZN(n382) );
  XOR2_X1 U442 ( .A(n382), .B(KEYINPUT93), .Z(n385) );
  XNOR2_X1 U443 ( .A(n383), .B(KEYINPUT94), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n389), .B(n388), .ZN(n512) );
  XNOR2_X1 U447 ( .A(n512), .B(KEYINPUT27), .ZN(n413) );
  XOR2_X1 U448 ( .A(KEYINPUT90), .B(G57GAT), .Z(n391) );
  XNOR2_X1 U449 ( .A(G1GAT), .B(G148GAT), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n391), .B(n390), .ZN(n397) );
  XOR2_X1 U451 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n395) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n409) );
  NAND2_X1 U455 ( .A1(G225GAT), .A2(G233GAT), .ZN(n403) );
  XOR2_X1 U456 ( .A(G162GAT), .B(G127GAT), .Z(n399) );
  XNOR2_X1 U457 ( .A(G141GAT), .B(G120GAT), .ZN(n398) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n401) );
  XOR2_X1 U459 ( .A(G29GAT), .B(G85GAT), .Z(n400) );
  XNOR2_X1 U460 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U462 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n405) );
  XNOR2_X1 U463 ( .A(KEYINPUT1), .B(KEYINPUT91), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U465 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U466 ( .A(n409), .B(n408), .Z(n418) );
  INV_X1 U467 ( .A(n418), .ZN(n510) );
  NAND2_X1 U468 ( .A1(n413), .A2(n510), .ZN(n410) );
  XOR2_X1 U469 ( .A(KEYINPUT95), .B(n410), .Z(n537) );
  XNOR2_X1 U470 ( .A(KEYINPUT96), .B(n522), .ZN(n411) );
  INV_X1 U471 ( .A(n515), .ZN(n524) );
  NAND2_X1 U472 ( .A1(n411), .A2(n524), .ZN(n421) );
  NOR2_X1 U473 ( .A1(n463), .A2(n515), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n412), .B(KEYINPUT26), .ZN(n558) );
  NAND2_X1 U475 ( .A1(n558), .A2(n413), .ZN(n417) );
  NAND2_X1 U476 ( .A1(n515), .A2(n512), .ZN(n414) );
  NAND2_X1 U477 ( .A1(n463), .A2(n414), .ZN(n415) );
  XOR2_X1 U478 ( .A(KEYINPUT25), .B(n415), .Z(n416) );
  NAND2_X1 U479 ( .A1(n417), .A2(n416), .ZN(n419) );
  NAND2_X1 U480 ( .A1(n419), .A2(n418), .ZN(n420) );
  NAND2_X1 U481 ( .A1(n421), .A2(n420), .ZN(n476) );
  NAND2_X1 U482 ( .A1(n574), .A2(n476), .ZN(n441) );
  XOR2_X1 U483 ( .A(n423), .B(n422), .Z(n425) );
  XNOR2_X1 U484 ( .A(G183GAT), .B(G71GAT), .ZN(n424) );
  XNOR2_X1 U485 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U486 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n427) );
  XNOR2_X1 U487 ( .A(G1GAT), .B(KEYINPUT14), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U489 ( .A(n429), .B(n428), .Z(n431) );
  XNOR2_X1 U490 ( .A(G22GAT), .B(G211GAT), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U492 ( .A(KEYINPUT76), .B(KEYINPUT78), .Z(n433) );
  NAND2_X1 U493 ( .A1(G231GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U495 ( .A(n435), .B(n434), .Z(n440) );
  XOR2_X1 U496 ( .A(G64GAT), .B(G78GAT), .Z(n437) );
  XNOR2_X1 U497 ( .A(G8GAT), .B(G155GAT), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n438), .B(KEYINPUT77), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n571) );
  XNOR2_X1 U501 ( .A(n442), .B(KEYINPUT37), .ZN(n509) );
  NOR2_X1 U502 ( .A1(n478), .A2(n509), .ZN(n443) );
  NAND2_X1 U503 ( .A1(n515), .A2(n495), .ZN(n447) );
  XOR2_X1 U504 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n445) );
  XNOR2_X1 U505 ( .A(G43GAT), .B(KEYINPUT104), .ZN(n444) );
  INV_X1 U506 ( .A(n497), .ZN(n560) );
  NAND2_X1 U507 ( .A1(n552), .A2(n560), .ZN(n449) );
  XOR2_X1 U508 ( .A(KEYINPUT46), .B(KEYINPUT109), .Z(n448) );
  XNOR2_X1 U509 ( .A(n449), .B(n448), .ZN(n451) );
  NOR2_X1 U510 ( .A1(n571), .A2(n545), .ZN(n450) );
  AND2_X1 U511 ( .A1(n451), .A2(n450), .ZN(n452) );
  XNOR2_X1 U512 ( .A(n452), .B(KEYINPUT47), .ZN(n458) );
  NAND2_X1 U513 ( .A1(n574), .A2(n571), .ZN(n454) );
  XOR2_X1 U514 ( .A(KEYINPUT45), .B(KEYINPUT110), .Z(n453) );
  XNOR2_X1 U515 ( .A(n454), .B(n453), .ZN(n456) );
  NOR2_X1 U516 ( .A1(n560), .A2(n567), .ZN(n455) );
  NAND2_X1 U517 ( .A1(n456), .A2(n455), .ZN(n457) );
  NAND2_X1 U518 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n459), .B(KEYINPUT48), .ZN(n535) );
  NAND2_X1 U520 ( .A1(n535), .A2(n512), .ZN(n461) );
  XOR2_X1 U521 ( .A(KEYINPUT115), .B(KEYINPUT54), .Z(n460) );
  XNOR2_X1 U522 ( .A(n461), .B(n460), .ZN(n462) );
  NAND2_X1 U523 ( .A1(n557), .A2(n463), .ZN(n465) );
  XOR2_X1 U524 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n464) );
  XNOR2_X1 U525 ( .A(n465), .B(n464), .ZN(n466) );
  INV_X1 U526 ( .A(KEYINPUT117), .ZN(n467) );
  NAND2_X1 U527 ( .A1(n555), .A2(n545), .ZN(n472) );
  XOR2_X1 U528 ( .A(KEYINPUT58), .B(KEYINPUT120), .Z(n470) );
  INV_X1 U529 ( .A(G190GAT), .ZN(n469) );
  XOR2_X1 U530 ( .A(KEYINPUT98), .B(KEYINPUT34), .Z(n481) );
  NAND2_X1 U531 ( .A1(n473), .A2(n571), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n474), .B(KEYINPUT79), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n475), .B(KEYINPUT16), .ZN(n477) );
  NAND2_X1 U534 ( .A1(n477), .A2(n476), .ZN(n498) );
  NOR2_X1 U535 ( .A1(n478), .A2(n498), .ZN(n479) );
  XOR2_X1 U536 ( .A(KEYINPUT97), .B(n479), .Z(n488) );
  NAND2_X1 U537 ( .A1(n488), .A2(n510), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U539 ( .A(G1GAT), .B(n482), .Z(G1324GAT) );
  XOR2_X1 U540 ( .A(G8GAT), .B(KEYINPUT99), .Z(n484) );
  NAND2_X1 U541 ( .A1(n488), .A2(n512), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U544 ( .A1(n488), .A2(n515), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(n487), .ZN(G1326GAT) );
  NAND2_X1 U547 ( .A1(n488), .A2(n517), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n489), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U549 ( .A1(n495), .A2(n510), .ZN(n492) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  NAND2_X1 U553 ( .A1(n495), .A2(n512), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n493), .B(KEYINPUT102), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G36GAT), .B(n494), .ZN(G1329GAT) );
  NAND2_X1 U556 ( .A1(n495), .A2(n517), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n496), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT42), .B(KEYINPUT105), .Z(n500) );
  NAND2_X1 U559 ( .A1(n552), .A2(n497), .ZN(n508) );
  NOR2_X1 U560 ( .A1(n498), .A2(n508), .ZN(n505) );
  NAND2_X1 U561 ( .A1(n505), .A2(n510), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(n501), .ZN(G1332GAT) );
  NAND2_X1 U564 ( .A1(n512), .A2(n505), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(KEYINPUT106), .ZN(n503) );
  XNOR2_X1 U566 ( .A(G64GAT), .B(n503), .ZN(G1333GAT) );
  NAND2_X1 U567 ( .A1(n505), .A2(n515), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n504), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U569 ( .A(G78GAT), .B(KEYINPUT43), .Z(n507) );
  NAND2_X1 U570 ( .A1(n505), .A2(n517), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(G1335GAT) );
  NOR2_X1 U572 ( .A1(n509), .A2(n508), .ZN(n518) );
  NAND2_X1 U573 ( .A1(n510), .A2(n518), .ZN(n511) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(n511), .ZN(G1336GAT) );
  XOR2_X1 U575 ( .A(G92GAT), .B(KEYINPUT107), .Z(n514) );
  NAND2_X1 U576 ( .A1(n518), .A2(n512), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(G1337GAT) );
  NAND2_X1 U578 ( .A1(n518), .A2(n515), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n516), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n520) );
  NAND2_X1 U581 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U582 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U583 ( .A(G106GAT), .B(n521), .Z(G1339GAT) );
  NAND2_X1 U584 ( .A1(n535), .A2(n522), .ZN(n523) );
  NOR2_X1 U585 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U586 ( .A(KEYINPUT111), .B(n525), .Z(n531) );
  NAND2_X1 U587 ( .A1(n531), .A2(n560), .ZN(n526) );
  XNOR2_X1 U588 ( .A(n526), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(G120GAT), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U590 ( .A1(n531), .A2(n552), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  NAND2_X1 U592 ( .A1(n531), .A2(n571), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n529), .B(KEYINPUT50), .ZN(n530) );
  XNOR2_X1 U594 ( .A(G127GAT), .B(n530), .ZN(G1342GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT112), .B(KEYINPUT51), .Z(n533) );
  NAND2_X1 U596 ( .A1(n531), .A2(n545), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U598 ( .A(G134GAT), .B(n534), .ZN(G1343GAT) );
  XOR2_X1 U599 ( .A(G141GAT), .B(KEYINPUT113), .Z(n539) );
  NAND2_X1 U600 ( .A1(n535), .A2(n558), .ZN(n536) );
  NOR2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n546), .A2(n560), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1344GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n541) );
  NAND2_X1 U605 ( .A1(n546), .A2(n552), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(n542), .ZN(G1345GAT) );
  NAND2_X1 U608 ( .A1(n546), .A2(n571), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n543), .B(KEYINPUT114), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G155GAT), .B(n544), .ZN(G1346GAT) );
  NAND2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n547), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U613 ( .A1(n560), .A2(n555), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G169GAT), .B(n548), .ZN(G1348GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT57), .B(KEYINPUT119), .Z(n550) );
  XNOR2_X1 U616 ( .A(G176GAT), .B(KEYINPUT118), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U618 ( .A(KEYINPUT56), .B(n551), .Z(n554) );
  NAND2_X1 U619 ( .A1(n555), .A2(n552), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1349GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n571), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n562) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(KEYINPUT121), .ZN(n575) );
  NAND2_X1 U626 ( .A1(n575), .A2(n560), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(n564) );
  INV_X1 U628 ( .A(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(n566) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(G1352GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n569) );
  NAND2_X1 U633 ( .A1(n575), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G204GAT), .B(n570), .ZN(G1353GAT) );
  XOR2_X1 U636 ( .A(G211GAT), .B(KEYINPUT125), .Z(n573) );
  NAND2_X1 U637 ( .A1(n575), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1354GAT) );
  XNOR2_X1 U639 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n579) );
  XOR2_X1 U640 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n577) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(G1355GAT) );
endmodule

