//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1336, new_n1337, new_n1338, new_n1339,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n207), .B(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n205), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT66), .ZN(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  AOI211_X1 g0023(.A(new_n209), .B(new_n217), .C1(new_n221), .C2(new_n223), .ZN(G361));
  XNOR2_X1  g0024(.A(G250), .B(G257), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT67), .ZN(new_n226));
  XOR2_X1   g0026(.A(G264), .B(G270), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n228), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G87), .B(G97), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G107), .B(G116), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  XNOR2_X1  g0041(.A(KEYINPUT3), .B(G33), .ZN(new_n242));
  INV_X1    g0042(.A(G1698), .ZN(new_n243));
  NAND3_X1  g0043(.A1(new_n242), .A2(G222), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n242), .A2(G223), .A3(G1698), .ZN(new_n245));
  INV_X1    g0045(.A(G77), .ZN(new_n246));
  OAI211_X1 g0046(.A(new_n244), .B(new_n245), .C1(new_n246), .C2(new_n242), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G1), .A3(G13), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(new_n249), .A3(G274), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n249), .A2(new_n253), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT69), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT69), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n249), .A2(new_n258), .A3(new_n253), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G226), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n251), .A2(new_n255), .A3(new_n261), .ZN(new_n262));
  OR2_X1    g0062(.A1(new_n262), .A2(G179), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n202), .A2(G20), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT71), .ZN(new_n265));
  INV_X1    g0065(.A(G58), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(KEYINPUT8), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(KEYINPUT8), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT8), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(KEYINPUT71), .A3(G58), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n219), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n271), .A2(new_n273), .B1(G150), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n264), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(KEYINPUT70), .A3(new_n218), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT70), .B1(new_n277), .B2(new_n218), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n283), .A2(new_n219), .A3(G1), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n277), .A2(new_n218), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT70), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n284), .B1(new_n287), .B2(new_n278), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n219), .A2(G1), .ZN(new_n289));
  INV_X1    g0089(.A(G50), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n288), .A2(new_n291), .B1(new_n290), .B2(new_n284), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n282), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n262), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n263), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n282), .A2(KEYINPUT9), .A3(new_n292), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT75), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n262), .A2(G200), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  INV_X1    g0100(.A(new_n292), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n287), .A2(new_n278), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(new_n264), .B2(new_n275), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n300), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT76), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n251), .A2(G190), .A3(new_n261), .A4(new_n255), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n299), .A2(new_n304), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n298), .A2(new_n307), .A3(KEYINPUT10), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT10), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT75), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n297), .B(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n307), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n296), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G68), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n274), .A2(G50), .B1(G20), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(new_n246), .B2(new_n272), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n281), .A2(new_n317), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n318), .A2(KEYINPUT11), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n284), .A2(new_n315), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT12), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(KEYINPUT11), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n288), .B(G68), .C1(G1), .C2(new_n219), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT77), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT14), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT13), .ZN(new_n329));
  INV_X1    g0129(.A(new_n255), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n260), .B2(G238), .ZN(new_n331));
  INV_X1    g0131(.A(G33), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT3), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT3), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G33), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n333), .A2(new_n335), .A3(G226), .A4(new_n243), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n333), .A2(new_n335), .A3(G232), .A4(G1698), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n250), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n329), .B1(new_n331), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n259), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n258), .B1(new_n249), .B2(new_n253), .ZN(new_n343));
  OAI21_X1  g0143(.A(G238), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AND4_X1   g0144(.A1(new_n329), .A2(new_n344), .A3(new_n340), .A4(new_n255), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n328), .B(G169), .C1(new_n341), .C2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(new_n340), .A3(new_n255), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT13), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n331), .A2(new_n329), .A3(new_n340), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(G179), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n349), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n328), .B1(new_n352), .B2(G169), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n327), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT74), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n242), .A2(G232), .A3(new_n243), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n242), .A2(G238), .A3(G1698), .ZN(new_n357));
  INV_X1    g0157(.A(G107), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n356), .B(new_n357), .C1(new_n358), .C2(new_n242), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n250), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n260), .A2(G244), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n255), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G200), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n289), .A2(new_n246), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n288), .A2(new_n365), .B1(new_n246), .B2(new_n284), .ZN(new_n366));
  XOR2_X1   g0166(.A(KEYINPUT15), .B(G87), .Z(new_n367));
  NAND3_X1  g0167(.A1(new_n367), .A2(KEYINPUT72), .A3(new_n273), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n269), .A2(G58), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n268), .A2(new_n369), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(new_n274), .B1(G20), .B2(G77), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT72), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT15), .B(G87), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n372), .B1(new_n373), .B2(new_n272), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n368), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n281), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT73), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT73), .B1(new_n375), .B2(new_n281), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n366), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n355), .B1(new_n364), .B2(new_n380), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n360), .A2(new_n255), .A3(new_n361), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G190), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n376), .B(new_n377), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n384), .A2(KEYINPUT74), .A3(new_n366), .A4(new_n363), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n352), .A2(G200), .ZN(new_n387));
  INV_X1    g0187(.A(G190), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n326), .B(new_n387), .C1(new_n388), .C2(new_n352), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n362), .A2(new_n294), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n362), .A2(G179), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n380), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n354), .A2(new_n386), .A3(new_n389), .A4(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n271), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(new_n289), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(new_n288), .B1(new_n284), .B2(new_n395), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n333), .A2(new_n335), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT7), .B1(new_n399), .B2(new_n219), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  AOI211_X1 g0201(.A(new_n401), .B(G20), .C1(new_n333), .C2(new_n335), .ZN(new_n402));
  OAI21_X1  g0202(.A(G68), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n266), .A2(new_n315), .ZN(new_n404));
  NOR2_X1   g0204(.A1(G58), .A2(G68), .ZN(new_n405));
  OAI21_X1  g0205(.A(G20), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n274), .A2(G159), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT16), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n302), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n403), .A2(KEYINPUT16), .A3(new_n409), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n398), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n333), .A2(new_n335), .A3(G223), .A4(new_n243), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n333), .A2(new_n335), .A3(G226), .A4(G1698), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G87), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n250), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n249), .A2(G232), .A3(new_n253), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n255), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT78), .B1(new_n422), .B2(G179), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n255), .A2(new_n420), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n250), .B2(new_n418), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT78), .ZN(new_n426));
  INV_X1    g0226(.A(G179), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n422), .A2(new_n294), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n423), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT18), .B1(new_n414), .B2(new_n430), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n423), .A2(new_n428), .A3(new_n429), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n401), .B1(new_n242), .B2(G20), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n399), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n315), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n411), .B1(new_n436), .B2(new_n408), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n413), .A2(new_n437), .A3(new_n281), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n397), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n432), .A2(new_n433), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n419), .A2(new_n421), .A3(new_n388), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n425), .B2(G200), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n438), .A2(new_n397), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT17), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n438), .A2(new_n442), .A3(KEYINPUT17), .A4(new_n397), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n431), .A2(new_n440), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n314), .A2(new_n394), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT81), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n358), .B1(new_n434), .B2(new_n435), .ZN(new_n451));
  INV_X1    g0251(.A(G97), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(new_n358), .A3(KEYINPUT6), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT6), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G97), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n358), .A2(KEYINPUT79), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT79), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G107), .ZN(new_n458));
  AND4_X1   g0258(.A1(new_n453), .A2(new_n455), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n453), .A2(new_n455), .B1(new_n456), .B2(new_n458), .ZN(new_n460));
  OAI21_X1  g0260(.A(G20), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n274), .A2(G77), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n451), .B1(new_n463), .B2(KEYINPUT80), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT80), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n461), .A2(new_n465), .A3(new_n462), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n302), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n284), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G97), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n252), .A2(G33), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n468), .B(new_n471), .C1(new_n279), .C2(new_n280), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n470), .B1(new_n472), .B2(new_n452), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n450), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n454), .A2(G97), .A3(G107), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n452), .A2(KEYINPUT6), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n457), .A2(G107), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n358), .A2(KEYINPUT79), .ZN(new_n478));
  OAI22_X1  g0278(.A1(new_n475), .A2(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n453), .A2(new_n455), .A3(new_n456), .A4(new_n458), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n219), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n462), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT80), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n451), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n483), .A2(new_n466), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n281), .ZN(new_n486));
  INV_X1    g0286(.A(new_n473), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(KEYINPUT81), .A3(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n333), .A2(new_n335), .A3(G244), .A4(new_n243), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n242), .A2(KEYINPUT4), .A3(G244), .A4(new_n243), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G283), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n242), .A2(G250), .A3(G1698), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n250), .ZN(new_n496));
  INV_X1    g0296(.A(G41), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n252), .B(G45), .C1(new_n497), .C2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT82), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n500), .B1(new_n501), .B2(G41), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n497), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n499), .A2(new_n504), .A3(G274), .A4(new_n249), .ZN(new_n505));
  INV_X1    g0305(.A(G45), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(G1), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n497), .A2(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n501), .A2(G41), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(G257), .A3(new_n249), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n496), .A2(new_n505), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(G200), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(G190), .B2(new_n512), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n474), .A2(new_n488), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n486), .A2(new_n487), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n496), .A2(new_n427), .A3(new_n505), .A4(new_n511), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT83), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n512), .A2(new_n294), .ZN(new_n520));
  INV_X1    g0320(.A(new_n511), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n495), .B2(new_n250), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT83), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n522), .A2(new_n523), .A3(new_n427), .A4(new_n505), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n517), .A2(new_n519), .A3(new_n520), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n516), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n333), .A2(new_n335), .A3(G264), .A4(G1698), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n333), .A2(new_n335), .A3(G257), .A4(new_n243), .ZN(new_n528));
  INV_X1    g0328(.A(G303), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n527), .B(new_n528), .C1(new_n529), .C2(new_n242), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n250), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n510), .A2(G270), .A3(new_n249), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n502), .A2(new_n503), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n249), .A2(G274), .A3(new_n509), .A4(new_n507), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(G200), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G116), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n252), .A2(new_n538), .A3(G13), .A4(G20), .ZN(new_n539));
  OR2_X1    g0339(.A1(new_n539), .A2(KEYINPUT87), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(KEYINPUT87), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n277), .A2(new_n218), .B1(G20), .B2(new_n538), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n493), .B(new_n219), .C1(G33), .C2(new_n452), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n543), .A2(KEYINPUT20), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT20), .B1(new_n543), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(KEYINPUT86), .B1(new_n472), .B2(new_n538), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT86), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n288), .A2(new_n549), .A3(G116), .A4(new_n471), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n547), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n505), .A2(new_n533), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n552), .A2(G190), .A3(new_n531), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n537), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT88), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n537), .A2(new_n551), .A3(KEYINPUT88), .A4(new_n553), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT21), .ZN(new_n559));
  OAI21_X1  g0359(.A(G169), .B1(new_n532), .B2(new_n536), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n560), .B2(new_n551), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n552), .A2(G179), .A3(new_n531), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n551), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n560), .A2(new_n551), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n563), .B1(new_n564), .B2(KEYINPUT21), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n558), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n472), .A2(new_n358), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n284), .A2(new_n358), .ZN(new_n568));
  XNOR2_X1  g0368(.A(new_n568), .B(KEYINPUT25), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n333), .A2(new_n335), .A3(new_n219), .A4(G87), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT22), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT22), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n242), .A2(new_n573), .A3(new_n219), .A4(G87), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT90), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n576), .B(KEYINPUT23), .C1(new_n219), .C2(G107), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n358), .A2(G20), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n576), .B1(new_n579), .B2(KEYINPUT23), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT23), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(new_n358), .A3(G20), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n219), .A2(G33), .A3(G116), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n578), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n575), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g0386(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n575), .A2(new_n585), .A3(new_n587), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT91), .B1(new_n591), .B2(new_n281), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n575), .A2(new_n585), .A3(new_n587), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n587), .B1(new_n575), .B2(new_n585), .ZN(new_n594));
  OAI211_X1 g0394(.A(KEYINPUT91), .B(new_n281), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n570), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n535), .A2(new_n534), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n510), .A2(G264), .A3(new_n249), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT92), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT92), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n510), .A2(new_n601), .A3(G264), .A4(new_n249), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n598), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n242), .A2(G257), .A3(G1698), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n242), .A2(G250), .A3(new_n243), .ZN(new_n605));
  INV_X1    g0405(.A(G294), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n604), .B(new_n605), .C1(new_n332), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n250), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT93), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n603), .A2(new_n608), .A3(new_n609), .A4(G179), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n603), .A2(G179), .A3(new_n608), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT93), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n294), .B1(new_n603), .B2(new_n608), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n611), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n597), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n249), .B1(G250), .B2(new_n507), .ZN(new_n619));
  INV_X1    g0419(.A(G274), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n619), .B1(new_n620), .B2(new_n507), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n333), .A2(new_n335), .A3(G238), .A4(new_n243), .ZN(new_n623));
  NAND2_X1  g0423(.A1(G33), .A2(G116), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n333), .A2(new_n335), .A3(G244), .A4(G1698), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT84), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n242), .A2(KEYINPUT84), .A3(G244), .A4(G1698), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n622), .B1(new_n630), .B2(new_n249), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n294), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n622), .B(new_n427), .C1(new_n630), .C2(new_n249), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT19), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n219), .B1(new_n338), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G87), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(new_n452), .A3(new_n358), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n333), .A2(new_n335), .A3(new_n219), .A4(G68), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n634), .B1(new_n272), .B2(new_n452), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n281), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n373), .A2(new_n284), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n288), .A2(new_n367), .A3(new_n471), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n632), .A2(new_n633), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n302), .A2(G87), .A3(new_n468), .A4(new_n471), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n642), .A3(new_n643), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n631), .B2(G200), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n628), .A2(new_n629), .ZN(new_n652));
  INV_X1    g0452(.A(new_n625), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n621), .B1(new_n654), .B2(new_n250), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n651), .A2(KEYINPUT85), .B1(G190), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n631), .A2(G200), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n649), .A2(new_n642), .A3(new_n643), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT85), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n648), .B1(new_n656), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n570), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n281), .B1(new_n593), .B2(new_n594), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n663), .B1(new_n666), .B2(new_n595), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n603), .A2(new_n608), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n513), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(G190), .B2(new_n668), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n618), .A2(new_n662), .A3(new_n671), .ZN(new_n672));
  NOR4_X1   g0472(.A1(new_n449), .A2(new_n526), .A3(new_n566), .A4(new_n672), .ZN(G372));
  INV_X1    g0473(.A(new_n296), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n351), .A2(new_n353), .ZN(new_n675));
  INV_X1    g0475(.A(new_n393), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n675), .A2(new_n327), .B1(new_n676), .B2(new_n389), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n445), .A2(new_n446), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n431), .B(new_n440), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT10), .B1(new_n298), .B2(new_n307), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n311), .A2(new_n312), .A3(new_n309), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n674), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n610), .B1(new_n613), .B2(new_n615), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n565), .B(new_n561), .C1(new_n667), .C2(new_n684), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n622), .B(G190), .C1(new_n630), .C2(new_n249), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n657), .A2(new_n658), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n647), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n667), .B2(new_n670), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n685), .A2(new_n689), .A3(new_n525), .A4(new_n516), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n647), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n519), .A2(new_n520), .A3(new_n524), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n294), .A2(new_n631), .B1(new_n644), .B2(new_n645), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n693), .A2(new_n633), .B1(new_n651), .B2(new_n686), .ZN(new_n694));
  AOI21_X1  g0494(.A(KEYINPUT81), .B1(new_n486), .B2(new_n487), .ZN(new_n695));
  AOI211_X1 g0495(.A(new_n450), .B(new_n473), .C1(new_n485), .C2(new_n281), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n692), .B(new_n694), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT26), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(KEYINPUT94), .A3(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n662), .A2(KEYINPUT26), .A3(new_n517), .A4(new_n692), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT94), .B1(new_n697), .B2(new_n698), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n691), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n683), .B1(new_n449), .B2(new_n704), .ZN(G369));
  NAND2_X1  g0505(.A1(new_n565), .A2(new_n561), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n252), .A2(new_n219), .A3(G13), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT27), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(KEYINPUT27), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G213), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G343), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n551), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n706), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n566), .B2(new_n714), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G330), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n667), .A2(new_n684), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n712), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n618), .A2(new_n671), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n667), .A2(new_n713), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n721), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n706), .A2(new_n713), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n725), .A2(new_n727), .B1(new_n719), .B2(new_n713), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n724), .A2(new_n728), .ZN(G399));
  INV_X1    g0529(.A(new_n206), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G41), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n637), .A2(G116), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(G1), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n222), .B2(new_n732), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n474), .A2(new_n488), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n737), .A2(KEYINPUT26), .A3(new_n692), .A4(new_n694), .ZN(new_n738));
  OAI211_X1 g0538(.A(KEYINPUT85), .B(new_n658), .C1(new_n655), .C2(new_n513), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n686), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n651), .A2(KEYINPUT85), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n647), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n698), .B1(new_n742), .B2(new_n525), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(new_n647), .A3(new_n690), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(KEYINPUT29), .A3(new_n713), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n703), .A2(new_n700), .A3(new_n699), .ZN(new_n747));
  INV_X1    g0547(.A(new_n691), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n712), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n746), .B1(new_n749), .B2(KEYINPUT29), .ZN(new_n750));
  INV_X1    g0550(.A(G330), .ZN(new_n751));
  AND3_X1   g0551(.A1(new_n618), .A2(new_n671), .A3(new_n662), .ZN(new_n752));
  INV_X1    g0552(.A(new_n526), .ZN(new_n753));
  INV_X1    g0553(.A(new_n566), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n752), .A2(new_n753), .A3(new_n754), .A4(new_n713), .ZN(new_n755));
  XOR2_X1   g0555(.A(KEYINPUT95), .B(KEYINPUT31), .Z(new_n756));
  AOI21_X1  g0556(.A(G179), .B1(new_n552), .B2(new_n531), .ZN(new_n757));
  AND4_X1   g0557(.A1(new_n512), .A2(new_n668), .A3(new_n757), .A4(new_n631), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n536), .B1(new_n250), .B2(new_n530), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n759), .A2(new_n603), .A3(G179), .A4(new_n608), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n654), .A2(new_n250), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n522), .A2(new_n761), .A3(new_n622), .ZN(new_n762));
  OAI21_X1  g0562(.A(KEYINPUT96), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n758), .B1(new_n763), .B2(KEYINPUT30), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT30), .ZN(new_n765));
  OAI211_X1 g0565(.A(KEYINPUT96), .B(new_n765), .C1(new_n760), .C2(new_n762), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n713), .B(new_n756), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n763), .A2(KEYINPUT30), .ZN(new_n768));
  INV_X1    g0568(.A(new_n758), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n768), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(KEYINPUT31), .B1(new_n770), .B2(new_n712), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n751), .B1(new_n755), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n750), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n736), .B1(new_n776), .B2(G1), .ZN(G364));
  NOR2_X1   g0577(.A1(new_n283), .A2(G20), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n252), .B1(new_n778), .B2(G45), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n731), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n718), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(G330), .B2(new_n716), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n242), .A2(G355), .A3(new_n206), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(G116), .B2(new_n206), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n730), .A2(new_n242), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n506), .B2(new_n223), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n240), .A2(G45), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n785), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n218), .B1(G20), .B2(new_n294), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n781), .B1(new_n790), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n427), .A2(G20), .A3(G190), .A4(G200), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G87), .ZN(new_n800));
  NAND2_X1  g0600(.A1(G20), .A2(G179), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT97), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n388), .A2(new_n513), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n242), .B(new_n800), .C1(new_n804), .C2(new_n290), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n219), .A2(G190), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n806), .A2(new_n427), .A3(G200), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT100), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n358), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n388), .A2(G200), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n802), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n805), .B(new_n812), .C1(G58), .C2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(G179), .A2(G200), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT99), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n219), .B1(new_n819), .B2(G190), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n802), .A2(new_n388), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n513), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n821), .A2(G97), .B1(G68), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n819), .A2(new_n806), .ZN(new_n825));
  INV_X1    g0625(.A(G159), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT32), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n816), .A2(new_n824), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n802), .A2(new_n388), .A3(new_n513), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n831), .A2(KEYINPUT98), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n831), .A2(KEYINPUT98), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(new_n246), .ZN(new_n835));
  XNOR2_X1  g0635(.A(KEYINPUT33), .B(G317), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n823), .A2(new_n836), .B1(new_n815), .B2(G322), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT101), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n821), .A2(G294), .B1(G311), .B2(new_n831), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n399), .B1(new_n529), .B2(new_n798), .ZN(new_n840));
  INV_X1    g0640(.A(new_n811), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(new_n841), .B2(G283), .ZN(new_n842));
  INV_X1    g0642(.A(new_n825), .ZN(new_n843));
  INV_X1    g0643(.A(new_n804), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n843), .A2(G329), .B1(G326), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n839), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n829), .A2(new_n835), .B1(new_n838), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n797), .B1(new_n847), .B2(new_n794), .ZN(new_n848));
  INV_X1    g0648(.A(new_n793), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n848), .B1(new_n716), .B2(new_n849), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n783), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(G396));
  OAI21_X1  g0652(.A(new_n380), .B1(new_n392), .B2(new_n712), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n386), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n392), .A2(KEYINPUT102), .A3(new_n380), .A4(new_n712), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n382), .A2(new_n427), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n362), .A2(new_n294), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n380), .A2(new_n856), .A3(new_n857), .A4(new_n712), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT102), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n854), .A2(new_n861), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n386), .A2(new_n853), .B1(new_n855), .B2(new_n860), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n863), .A2(new_n712), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n749), .A2(new_n862), .B1(new_n704), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n781), .B1(new_n866), .B2(new_n774), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n774), .B2(new_n866), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n794), .A2(new_n791), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n781), .B1(G77), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n834), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(G116), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n811), .A2(new_n636), .B1(new_n529), .B2(new_n804), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(G294), .B2(new_n815), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n823), .A2(G283), .ZN(new_n875));
  INV_X1    g0675(.A(G311), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n399), .B1(new_n358), .B2(new_n798), .C1(new_n825), .C2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(G97), .B2(new_n821), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n872), .A2(new_n874), .A3(new_n875), .A4(new_n878), .ZN(new_n879));
  AOI22_X1  g0679(.A1(G137), .A2(new_n844), .B1(new_n815), .B2(G143), .ZN(new_n880));
  INV_X1    g0680(.A(G150), .ZN(new_n881));
  INV_X1    g0681(.A(new_n823), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n880), .B1(new_n881), .B2(new_n882), .C1(new_n834), .C2(new_n826), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT34), .Z(new_n884));
  OAI21_X1  g0684(.A(new_n242), .B1(new_n290), .B2(new_n798), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n811), .A2(new_n315), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n885), .B(new_n886), .C1(G132), .C2(new_n843), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n266), .B2(new_n820), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n879), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n870), .B1(new_n889), .B2(new_n794), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n792), .B2(new_n862), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n891), .B(KEYINPUT103), .Z(new_n892));
  NAND2_X1  g0692(.A1(new_n868), .A2(new_n892), .ZN(G384));
  NOR2_X1   g0693(.A1(new_n459), .A2(new_n460), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n896), .A2(G116), .A3(new_n221), .A4(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT36), .ZN(new_n899));
  OAI21_X1  g0699(.A(G77), .B1(new_n266), .B2(new_n315), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n900), .A2(new_n222), .B1(G50), .B2(new_n315), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(G1), .A3(new_n283), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT104), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n448), .B(new_n746), .C1(new_n749), .C2(KEYINPUT29), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n683), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT108), .Z(new_n907));
  INV_X1    g0707(.A(new_n710), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n431), .B2(new_n440), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n393), .A2(new_n712), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n699), .A2(new_n700), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n647), .B(new_n690), .C1(new_n911), .C2(new_n702), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n910), .B1(new_n912), .B2(new_n864), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n326), .A2(new_n713), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n354), .A2(new_n915), .A3(new_n389), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(new_n354), .B2(new_n389), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n439), .A2(new_n908), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n447), .A2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n430), .A2(new_n710), .B1(new_n438), .B2(new_n397), .ZN(new_n923));
  INV_X1    g0723(.A(new_n443), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT37), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n432), .A2(new_n439), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT37), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n926), .A2(new_n927), .A3(new_n443), .A4(new_n920), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n922), .A2(KEYINPUT38), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n922), .B2(new_n929), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n909), .B1(new_n919), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT39), .B1(new_n930), .B2(new_n931), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT105), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(KEYINPUT105), .B(KEYINPUT39), .C1(new_n930), .C2(new_n931), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT107), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n414), .A2(KEYINPUT106), .A3(new_n442), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT106), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n443), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n938), .B(KEYINPUT37), .C1(new_n942), .C2(new_n923), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n443), .B(KEYINPUT106), .ZN(new_n944));
  INV_X1    g0744(.A(new_n923), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n927), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n928), .A2(KEYINPUT107), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n922), .B(new_n943), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT38), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n930), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT39), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n936), .A2(new_n937), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n675), .A2(new_n327), .A3(new_n713), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n933), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n907), .B(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n930), .B1(new_n949), .B2(new_n948), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n354), .A2(new_n389), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n914), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n354), .A2(new_n915), .A3(new_n389), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n863), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR4_X1   g0764(.A1(new_n672), .A2(new_n526), .A3(new_n566), .A4(new_n712), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n770), .A2(KEYINPUT31), .A3(new_n712), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n713), .B1(new_n764), .B2(new_n766), .ZN(new_n967));
  INV_X1    g0767(.A(new_n756), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n964), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(KEYINPUT40), .B1(new_n960), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n862), .B1(new_n916), .B2(new_n917), .ZN(new_n972));
  INV_X1    g0772(.A(new_n969), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n972), .B1(new_n973), .B2(new_n755), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT40), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n974), .A2(new_n932), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n973), .A2(new_n755), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n978), .A2(new_n448), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n751), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n979), .B2(new_n977), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n959), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n252), .B2(new_n778), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n959), .A2(new_n981), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n904), .B1(new_n983), .B2(new_n984), .ZN(G367));
  NOR2_X1   g0785(.A1(new_n695), .A2(new_n696), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n516), .B(new_n525), .C1(new_n986), .C2(new_n713), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n737), .A2(new_n692), .A3(new_n712), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n721), .A2(new_n726), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT109), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n989), .A2(KEYINPUT109), .A3(new_n990), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(KEYINPUT42), .ZN(new_n996));
  INV_X1    g0796(.A(new_n989), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n525), .B1(new_n997), .B2(new_n618), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n713), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT43), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n694), .B1(new_n658), .B2(new_n713), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n648), .A2(new_n650), .A3(new_n712), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT42), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n993), .A2(new_n1006), .A3(new_n994), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1000), .A2(new_n1001), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n996), .A2(new_n1007), .A3(new_n999), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1005), .A2(new_n1001), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1004), .A2(KEYINPUT43), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n724), .A2(new_n997), .ZN(new_n1013));
  AND3_X1   g0813(.A1(new_n1008), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1013), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n731), .B(KEYINPUT41), .Z(new_n1017));
  INV_X1    g0817(.A(KEYINPUT45), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n725), .A2(new_n727), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n618), .B2(new_n712), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1018), .B1(new_n1020), .B2(new_n997), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n728), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1020), .A2(KEYINPUT44), .A3(new_n997), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT44), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n728), .B2(new_n989), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1023), .A2(new_n724), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT110), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n724), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n720), .B(new_n726), .C1(new_n721), .C2(new_n722), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1019), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT111), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1036), .B1(new_n1037), .B2(new_n717), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n718), .A2(KEYINPUT111), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1036), .A2(new_n718), .A3(KEYINPUT111), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1042), .A2(new_n750), .A3(new_n774), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1031), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1034), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1017), .B1(new_n1046), .B2(new_n776), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1016), .B1(new_n1047), .B2(new_n780), .ZN(new_n1048));
  INV_X1    g0848(.A(G317), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n399), .B1(new_n825), .B2(new_n1049), .C1(new_n820), .C2(new_n358), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n841), .A2(G97), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n876), .B2(new_n804), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1050), .B(new_n1052), .C1(G303), .C2(new_n815), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT46), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n798), .B2(new_n538), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n799), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(new_n882), .C2(new_n606), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1058), .A2(KEYINPUT112), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(KEYINPUT112), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n871), .A2(G283), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1053), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n834), .A2(new_n290), .ZN(new_n1063));
  INV_X1    g0863(.A(G143), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n804), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n811), .A2(new_n246), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(G137), .C2(new_n843), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n242), .B1(new_n266), .B2(new_n798), .C1(new_n814), .C2(new_n881), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G68), .B2(new_n821), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1067), .B(new_n1069), .C1(new_n826), .C2(new_n882), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1062), .B1(new_n1063), .B2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT47), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n794), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n781), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n228), .A2(new_n787), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n796), .B1(new_n730), .B2(new_n367), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1073), .B(new_n1077), .C1(new_n849), .C2(new_n1004), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1048), .A2(new_n1078), .ZN(G387));
  NAND3_X1  g0879(.A1(new_n775), .A2(new_n1041), .A3(new_n1040), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1080), .A2(KEYINPUT116), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(KEYINPUT116), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1082), .A2(new_n731), .A3(new_n1043), .A4(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n799), .A2(G77), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1051), .A2(new_n242), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n271), .B2(new_n823), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n290), .A2(new_n814), .B1(new_n804), .B2(new_n826), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G150), .B2(new_n843), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n820), .A2(new_n373), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G68), .B2(new_n831), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n242), .B1(new_n843), .B2(G326), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n814), .A2(new_n1049), .ZN(new_n1094));
  XOR2_X1   g0894(.A(KEYINPUT114), .B(G322), .Z(new_n1095));
  AOI21_X1  g0895(.A(new_n1094), .B1(new_n844), .B2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1096), .B1(new_n876), .B2(new_n882), .C1(new_n834), .C2(new_n529), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT48), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n821), .A2(G283), .B1(G294), .B2(new_n799), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT49), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1093), .B1(new_n538), .B2(new_n811), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1092), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT115), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n794), .A3(new_n1109), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n733), .A2(new_n730), .A3(new_n399), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n358), .B2(new_n730), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT113), .Z(new_n1113));
  NOR2_X1   g0913(.A1(new_n232), .A2(new_n506), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n370), .A2(new_n290), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT50), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n733), .B(new_n506), .C1(new_n315), .C2(new_n246), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n786), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1113), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1074), .B1(new_n1119), .B2(new_n795), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1110), .B(new_n1120), .C1(new_n723), .C2(new_n849), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1042), .A2(new_n780), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1084), .A2(new_n1124), .ZN(G393));
  INV_X1    g0925(.A(new_n1028), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n724), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n1126), .A2(new_n779), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT117), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n997), .A2(new_n793), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n237), .A2(new_n786), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n795), .B1(new_n452), .B2(new_n206), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n781), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n820), .A2(new_n246), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n399), .B1(new_n799), .B2(G68), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n825), .B2(new_n1064), .C1(new_n811), .C2(new_n636), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(G50), .C2(new_n823), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n871), .A2(new_n370), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n881), .A2(new_n804), .B1(new_n814), .B2(new_n826), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT51), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n876), .A2(new_n814), .B1(new_n804), .B2(new_n1049), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT52), .Z(new_n1144));
  INV_X1    g0944(.A(G283), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n399), .B1(new_n1145), .B2(new_n798), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1146), .B(new_n812), .C1(new_n843), .C2(new_n1095), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n821), .A2(G116), .B1(G294), .B2(new_n831), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1147), .B(new_n1148), .C1(new_n529), .C2(new_n882), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1142), .B1(new_n1144), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1134), .B1(new_n1150), .B2(new_n794), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1131), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1129), .A2(new_n1130), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1152), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT117), .B1(new_n1128), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1043), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1046), .A2(new_n731), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(G390));
  INV_X1    g0959(.A(KEYINPUT119), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n745), .A2(new_n713), .A3(new_n862), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n910), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n918), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n960), .A2(new_n956), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n773), .A2(new_n862), .A3(new_n1164), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1162), .B1(new_n704), .B2(new_n865), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n956), .B1(new_n1169), .B2(new_n1164), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1167), .B(new_n1168), .C1(new_n1170), .C2(new_n954), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n936), .A2(new_n937), .A3(new_n953), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n955), .B1(new_n913), .B2(new_n918), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1172), .A2(new_n1173), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n964), .B(G330), .C1(new_n965), .C2(new_n969), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1171), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1164), .B1(new_n773), .B2(new_n862), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1175), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1169), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1180));
  OAI211_X1 g0980(.A(G330), .B(new_n862), .C1(new_n965), .C2(new_n969), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n918), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(new_n1182), .A3(new_n1168), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1179), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n978), .A2(G330), .A3(new_n448), .ZN(new_n1185));
  AOI21_X1  g0985(.A(KEYINPUT29), .B1(new_n912), .B2(new_n713), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n746), .A2(new_n448), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n683), .B(new_n1185), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT118), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n905), .A2(KEYINPUT118), .A3(new_n683), .A4(new_n1185), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1184), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1160), .B1(new_n1176), .B2(new_n1192), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1184), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1167), .B1(new_n1170), .B2(new_n954), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n1178), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1194), .A2(KEYINPUT119), .A3(new_n1171), .A4(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1193), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n732), .B1(new_n1176), .B2(new_n1192), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1176), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1172), .A2(new_n791), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n781), .B1(new_n271), .B2(new_n869), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n799), .A2(G150), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n399), .B1(new_n1204), .B2(KEYINPUT53), .ZN(new_n1205));
  INV_X1    g1005(.A(G137), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1205), .B1(KEYINPUT53), .B2(new_n1204), .C1(new_n882), .C2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G159), .B2(new_n821), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(KEYINPUT54), .B(G143), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n871), .A2(new_n1210), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n841), .A2(G50), .B1(G128), .B2(new_n844), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n843), .A2(G125), .B1(G132), .B2(new_n815), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1208), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n834), .A2(new_n452), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n800), .A2(new_n399), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1135), .A2(new_n886), .A3(new_n1216), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n825), .A2(new_n606), .B1(new_n1145), .B2(new_n804), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G116), .B2(new_n815), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1217), .B(new_n1219), .C1(new_n358), .C2(new_n882), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1214), .B1(new_n1215), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1203), .B1(new_n1221), .B2(new_n794), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1201), .A2(new_n780), .B1(new_n1202), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1200), .A2(new_n1223), .ZN(G378));
  OAI21_X1  g1024(.A(new_n781), .B1(G50), .B2(new_n869), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n242), .A2(G41), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1085), .B(new_n1226), .C1(new_n804), .C2(new_n538), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n811), .A2(new_n266), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(G283), .C2(new_n843), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n315), .B2(new_n820), .C1(new_n373), .C2(new_n830), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n815), .A2(KEYINPUT120), .A3(G107), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT120), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n814), .B2(new_n358), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1231), .B(new_n1233), .C1(new_n882), .C2(new_n452), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1230), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT58), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n821), .A2(G150), .B1(G132), .B2(new_n823), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n1206), .B2(new_n830), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n844), .A2(G125), .B1(new_n799), .B2(new_n1210), .ZN(new_n1240));
  INV_X1    g1040(.A(G128), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1240), .B1(new_n1241), .B2(new_n814), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1239), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1244), .A2(KEYINPUT59), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(KEYINPUT59), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n332), .B(new_n497), .C1(new_n811), .C2(new_n826), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G124), .B2(new_n843), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1226), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1251), .B(new_n290), .C1(G33), .C2(G41), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1237), .A2(new_n1249), .A3(new_n1250), .A4(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1225), .B1(new_n1253), .B2(new_n794), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n293), .A2(new_n908), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n682), .B2(new_n296), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1257), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n674), .B(new_n1259), .C1(new_n680), .C2(new_n681), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1256), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n314), .A2(new_n1259), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n682), .A2(new_n296), .A3(new_n1257), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1255), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1261), .A2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1254), .B1(new_n792), .B2(new_n1265), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT121), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT122), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1265), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n751), .B(new_n1269), .C1(new_n971), .C2(new_n976), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1265), .B1(new_n977), .B2(G330), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n958), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n950), .A2(new_n951), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n975), .B1(new_n974), .B2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n975), .B1(new_n930), .B2(new_n931), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n970), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(G330), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1269), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n977), .A2(G330), .A3(new_n1265), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1278), .A2(new_n1279), .A3(new_n957), .A4(new_n933), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1272), .A2(new_n1280), .A3(KEYINPUT123), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT123), .B1(new_n1272), .B2(new_n1280), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1268), .B1(new_n1283), .B2(new_n780), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT124), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT124), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1190), .A2(new_n1191), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1198), .A2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT57), .B1(new_n1291), .B2(new_n1283), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1289), .B1(new_n1193), .B2(new_n1197), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1272), .A2(new_n1280), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(KEYINPUT57), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n731), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1284), .B1(new_n1292), .B2(new_n1296), .ZN(G375));
  AOI21_X1  g1097(.A(new_n1184), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1298));
  OR3_X1    g1098(.A1(new_n1194), .A2(new_n1298), .A3(new_n1017), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n918), .A2(new_n791), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n781), .B1(G68), .B2(new_n869), .ZN(new_n1301));
  OAI22_X1  g1101(.A1(new_n825), .A2(new_n1241), .B1(new_n1206), .B2(new_n814), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n242), .B1(new_n826), .B2(new_n798), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1302), .A2(new_n1228), .A3(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n844), .A2(KEYINPUT126), .A3(G132), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT126), .B1(new_n844), .B2(G132), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(G150), .B2(new_n831), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n821), .A2(G50), .B1(new_n823), .B2(new_n1210), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1304), .A2(new_n1305), .A3(new_n1307), .A4(new_n1308), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n823), .A2(G116), .B1(new_n844), .B2(G294), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1310), .B1(new_n834), .B2(new_n358), .ZN(new_n1311));
  XOR2_X1   g1111(.A(new_n1311), .B(KEYINPUT125), .Z(new_n1312));
  OAI22_X1  g1112(.A1(new_n825), .A2(new_n529), .B1(new_n1145), .B2(new_n814), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n399), .B1(new_n452), .B2(new_n798), .ZN(new_n1314));
  OR4_X1    g1114(.A1(new_n1066), .A2(new_n1090), .A3(new_n1313), .A4(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1309), .B1(new_n1312), .B2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1301), .B1(new_n1316), .B2(new_n794), .ZN(new_n1317));
  AOI22_X1  g1117(.A1(new_n1184), .A2(new_n780), .B1(new_n1300), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1299), .A2(new_n1318), .ZN(G381));
  AND2_X1   g1119(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(G393), .A2(G396), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1320), .A2(new_n868), .A3(new_n892), .A4(new_n1321), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1322), .A2(G387), .A3(G381), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1268), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT123), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1294), .A2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1272), .A2(new_n1280), .A3(KEYINPUT123), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1324), .B1(new_n1328), .B2(new_n779), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1295), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n732), .B1(new_n1291), .B2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT57), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1332), .B1(new_n1328), .B2(new_n1293), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1329), .B1(new_n1331), .B2(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1323), .A2(new_n1200), .A3(new_n1223), .A4(new_n1334), .ZN(G407));
  INV_X1    g1135(.A(G378), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n711), .A2(G213), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1334), .A2(new_n1336), .A3(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(G407), .A2(G213), .A3(new_n1339), .ZN(G409));
  OAI211_X1 g1140(.A(G378), .B(new_n1284), .C1(new_n1292), .C2(new_n1296), .ZN(new_n1341));
  NOR3_X1   g1141(.A1(new_n1328), .A2(new_n1293), .A3(new_n1017), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n779), .B1(new_n1272), .B2(new_n1280), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1343), .A2(new_n1267), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1336), .B1(new_n1342), .B2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1341), .A2(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1298), .B1(KEYINPUT60), .B2(new_n1192), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1285), .A2(KEYINPUT60), .A3(new_n1179), .A4(new_n1183), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n731), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1318), .B1(new_n1348), .B2(new_n1350), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1351), .A2(new_n868), .A3(new_n892), .ZN(new_n1352));
  OAI211_X1 g1152(.A(G384), .B(new_n1318), .C1(new_n1348), .C2(new_n1350), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1347), .A2(new_n1337), .A3(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(KEYINPUT62), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT61), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1338), .B1(new_n1341), .B2(new_n1346), .ZN(new_n1359));
  INV_X1    g1159(.A(KEYINPUT62), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1359), .A2(new_n1360), .A3(new_n1355), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1338), .A2(G2897), .ZN(new_n1362));
  XNOR2_X1  g1162(.A(new_n1354), .B(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1017), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1291), .A2(new_n1283), .A3(new_n1364), .ZN(new_n1365));
  AOI21_X1  g1165(.A(G378), .B1(new_n1365), .B2(new_n1344), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n1366), .B1(new_n1334), .B2(G378), .ZN(new_n1367));
  OAI21_X1  g1167(.A(new_n1363), .B1(new_n1367), .B2(new_n1338), .ZN(new_n1368));
  NAND4_X1  g1168(.A1(new_n1357), .A2(new_n1358), .A3(new_n1361), .A4(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(G387), .A2(new_n1320), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n851), .B1(new_n1084), .B2(new_n1124), .ZN(new_n1371));
  NOR2_X1   g1171(.A1(new_n1321), .A2(new_n1371), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(G390), .A2(new_n1048), .A3(new_n1078), .ZN(new_n1373));
  AND3_X1   g1173(.A1(new_n1370), .A2(new_n1372), .A3(new_n1373), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n1372), .B1(new_n1370), .B2(new_n1373), .ZN(new_n1375));
  NOR2_X1   g1175(.A1(new_n1374), .A2(new_n1375), .ZN(new_n1376));
  INV_X1    g1176(.A(new_n1376), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1369), .A2(new_n1377), .ZN(new_n1378));
  INV_X1    g1178(.A(new_n1362), .ZN(new_n1379));
  XNOR2_X1  g1179(.A(new_n1354), .B(new_n1379), .ZN(new_n1380));
  OAI211_X1 g1180(.A(new_n1376), .B(new_n1358), .C1(new_n1359), .C2(new_n1380), .ZN(new_n1381));
  INV_X1    g1181(.A(new_n1381), .ZN(new_n1382));
  AOI211_X1 g1182(.A(new_n1338), .B(new_n1354), .C1(new_n1341), .C2(new_n1346), .ZN(new_n1383));
  OAI21_X1  g1183(.A(KEYINPUT127), .B1(new_n1383), .B2(KEYINPUT63), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1383), .A2(KEYINPUT63), .ZN(new_n1385));
  INV_X1    g1185(.A(KEYINPUT127), .ZN(new_n1386));
  INV_X1    g1186(.A(KEYINPUT63), .ZN(new_n1387));
  NAND3_X1  g1187(.A1(new_n1356), .A2(new_n1386), .A3(new_n1387), .ZN(new_n1388));
  NAND4_X1  g1188(.A1(new_n1382), .A2(new_n1384), .A3(new_n1385), .A4(new_n1388), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1378), .A2(new_n1389), .ZN(G405));
  NOR2_X1   g1190(.A1(new_n1334), .A2(G378), .ZN(new_n1391));
  INV_X1    g1191(.A(new_n1391), .ZN(new_n1392));
  NAND3_X1  g1192(.A1(new_n1392), .A2(new_n1341), .A3(new_n1354), .ZN(new_n1393));
  INV_X1    g1193(.A(new_n1341), .ZN(new_n1394));
  OAI21_X1  g1194(.A(new_n1355), .B1(new_n1391), .B2(new_n1394), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1393), .A2(new_n1395), .ZN(new_n1396));
  XNOR2_X1  g1196(.A(new_n1396), .B(new_n1377), .ZN(G402));
endmodule


