//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990, new_n991;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n202));
  XOR2_X1   g001(.A(G15gat), .B(G43gat), .Z(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G227gat), .A2(G233gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT25), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT23), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT24), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  OAI221_X1 g013(.A(new_n208), .B1(KEYINPUT64), .B2(new_n210), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n209), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n220), .A2(new_n221), .B1(KEYINPUT23), .B2(new_n209), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n207), .B1(new_n215), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(KEYINPUT66), .B(G183gat), .Z(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(G190gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(new_n213), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n220), .A2(KEYINPUT25), .A3(new_n210), .A4(new_n208), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT27), .B(G183gat), .Z(new_n230));
  OAI21_X1  g029(.A(KEYINPUT28), .B1(new_n230), .B2(G190gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n216), .A2(KEYINPUT26), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT26), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n208), .B1(new_n209), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n231), .B(new_n211), .C1(new_n232), .C2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n224), .A2(KEYINPUT27), .ZN(new_n238));
  NOR2_X1   g037(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n229), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G113gat), .B(G120gat), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT1), .B1(new_n243), .B2(KEYINPUT68), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(KEYINPUT68), .B2(new_n243), .ZN(new_n245));
  NOR2_X1   g044(.A1(G127gat), .A2(G134gat), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT67), .B(G134gat), .Z(new_n247));
  AOI21_X1  g046(.A(new_n246), .B1(new_n247), .B2(G127gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G113gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G120gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT69), .B(G120gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n251), .B1(new_n252), .B2(new_n250), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n254));
  AND2_X1   g053(.A1(G127gat), .A2(G134gat), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n253), .B(new_n254), .C1(new_n255), .C2(new_n246), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n249), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n223), .A2(new_n228), .B1(new_n236), .B2(new_n240), .ZN(new_n259));
  INV_X1    g058(.A(new_n257), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n206), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n205), .B1(new_n262), .B2(KEYINPUT33), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT32), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n258), .A2(new_n261), .ZN(new_n267));
  INV_X1    g066(.A(new_n206), .ZN(new_n268));
  AOI221_X4 g067(.A(new_n264), .B1(KEYINPUT33), .B2(new_n205), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n202), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT34), .B1(new_n267), .B2(new_n268), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT34), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n258), .A2(new_n261), .A3(new_n272), .A4(new_n206), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n274), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n202), .B(new_n276), .C1(new_n266), .C2(new_n269), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G78gat), .B(G106gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT83), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT76), .B(G148gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G141gat), .ZN(new_n283));
  INV_X1    g082(.A(G148gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(G141gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT77), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n283), .A2(KEYINPUT77), .A3(new_n286), .ZN(new_n290));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT2), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n289), .A2(new_n290), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT75), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n292), .B1(new_n296), .B2(new_n291), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n296), .B2(new_n291), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n284), .A2(G141gat), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n286), .A2(new_n299), .B1(KEYINPUT75), .B2(KEYINPUT2), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT3), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT29), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G197gat), .B(G204gat), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n306), .A2(KEYINPUT72), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(KEYINPUT72), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n304), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n289), .A2(new_n290), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n294), .A2(new_n291), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n301), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n311), .A2(KEYINPUT29), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(KEYINPUT3), .ZN(new_n320));
  INV_X1    g119(.A(G228gat), .ZN(new_n321));
  INV_X1    g120(.A(G233gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n313), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n316), .A2(new_n303), .A3(new_n317), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n311), .B1(new_n329), .B2(KEYINPUT84), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT84), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n304), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n320), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n326), .B1(new_n333), .B2(new_n323), .ZN(new_n334));
  INV_X1    g133(.A(G22gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n281), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n320), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n312), .B1(new_n304), .B2(new_n331), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n329), .A2(KEYINPUT84), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI22_X1  g139(.A1(new_n340), .A2(new_n324), .B1(new_n313), .B2(new_n325), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(G22gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n280), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT83), .B1(new_n341), .B2(G22gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n334), .A2(new_n335), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n345), .A3(new_n279), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT31), .B(G50gat), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n343), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n347), .B1(new_n343), .B2(new_n346), .ZN(new_n349));
  OAI211_X1 g148(.A(KEYINPUT35), .B(new_n278), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n343), .A2(new_n346), .ZN(new_n351));
  INV_X1    g150(.A(new_n347), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n343), .A2(new_n346), .A3(new_n347), .ZN(new_n354));
  INV_X1    g153(.A(new_n266), .ZN(new_n355));
  INV_X1    g154(.A(new_n269), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n355), .A2(KEYINPUT71), .A3(new_n356), .A4(new_n274), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n274), .A2(KEYINPUT71), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT71), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n271), .A2(new_n359), .A3(new_n273), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n358), .B(new_n360), .C1(new_n266), .C2(new_n269), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT36), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n275), .A2(KEYINPUT36), .A3(new_n277), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n353), .A2(new_n354), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n257), .A2(KEYINPUT78), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n249), .A2(new_n370), .A3(new_n256), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT3), .B1(new_n295), .B2(new_n301), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n373), .A3(new_n327), .ZN(new_n374));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n318), .A2(KEYINPUT4), .A3(new_n257), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n378), .B1(new_n302), .B2(new_n260), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n368), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n302), .A2(new_n260), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT4), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n302), .A2(new_n378), .A3(new_n260), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n385), .A2(KEYINPUT79), .A3(new_n375), .A4(new_n374), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n375), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n302), .B1(new_n369), .B2(new_n371), .ZN(new_n389));
  INV_X1    g188(.A(new_n382), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT5), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n387), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n380), .A2(KEYINPUT80), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT80), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n385), .A2(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n376), .A2(KEYINPUT5), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G1gat), .B(G29gat), .ZN(new_n401));
  INV_X1    g200(.A(G85gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT0), .B(G57gat), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n403), .B(new_n404), .Z(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n394), .A2(new_n400), .A3(new_n406), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n399), .A2(new_n397), .A3(new_n395), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n392), .B1(new_n381), .B2(new_n386), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT81), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n407), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n394), .A2(new_n400), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(new_n405), .A3(new_n412), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n242), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n259), .A2(G226gat), .A3(G233gat), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n311), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(new_n420), .A3(new_n311), .ZN(new_n423));
  XOR2_X1   g222(.A(G64gat), .B(G92gat), .Z(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(KEYINPUT73), .ZN(new_n425));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  NAND3_X1  g226(.A1(new_n422), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT30), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT74), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(KEYINPUT74), .A3(new_n429), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n427), .ZN(new_n435));
  INV_X1    g234(.A(new_n423), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n435), .B1(new_n436), .B2(new_n421), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n428), .A2(new_n429), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n434), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n417), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n417), .A2(new_n439), .A3(KEYINPUT82), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n367), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n364), .A2(new_n365), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n446), .B1(new_n354), .B2(new_n353), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT37), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n437), .B1(new_n448), .B2(new_n427), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n448), .B1(new_n436), .B2(KEYINPUT86), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n422), .A2(new_n423), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n450), .B1(new_n451), .B2(KEYINPUT86), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT38), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n449), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n435), .B1(new_n451), .B2(KEYINPUT37), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n448), .B1(new_n422), .B2(new_n423), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT38), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n457), .A3(new_n428), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT87), .B1(new_n410), .B2(new_n411), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT87), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n415), .A2(new_n460), .A3(KEYINPUT6), .A4(new_n405), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n407), .A2(new_n410), .A3(new_n411), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT85), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n407), .A2(new_n410), .A3(KEYINPUT85), .A4(new_n411), .ZN(new_n465));
  AOI221_X4 g264(.A(new_n458), .B1(new_n459), .B2(new_n461), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT40), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n398), .A2(new_n374), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT39), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n469), .A3(new_n388), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n406), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n375), .B1(new_n398), .B2(new_n374), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n389), .A2(new_n390), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT39), .B1(new_n473), .B2(new_n388), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n467), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n405), .B1(new_n472), .B2(new_n469), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n477), .B(KEYINPUT40), .C1(new_n472), .C2(new_n474), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n434), .A2(new_n437), .A3(new_n438), .ZN(new_n479));
  AND4_X1   g278(.A1(new_n410), .A2(new_n476), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n447), .B1(new_n466), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT35), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n362), .B(new_n439), .C1(new_n348), .C2(new_n349), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n464), .A2(new_n465), .B1(new_n459), .B2(new_n461), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n445), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  AND2_X1   g285(.A1(G232gat), .A2(G233gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT41), .ZN(new_n488));
  INV_X1    g287(.A(G29gat), .ZN(new_n489));
  INV_X1    g288(.A(G36gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NOR3_X1   g293(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G43gat), .B(G50gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(KEYINPUT15), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(KEYINPUT88), .A2(KEYINPUT15), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n497), .B2(KEYINPUT89), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT90), .B1(new_n494), .B2(new_n495), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT14), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(new_n489), .A3(new_n490), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT90), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(new_n493), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n501), .A2(new_n492), .A3(new_n502), .A4(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT88), .ZN(new_n508));
  INV_X1    g307(.A(G50gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(G43gat), .ZN(new_n510));
  INV_X1    g309(.A(G43gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(G50gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT89), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n510), .A2(new_n512), .A3(KEYINPUT15), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n499), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n498), .B1(new_n507), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G85gat), .A2(G92gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g321(.A1(G99gat), .A2(G106gat), .ZN(new_n523));
  INV_X1    g322(.A(G92gat), .ZN(new_n524));
  AOI22_X1  g323(.A1(KEYINPUT8), .A2(new_n523), .B1(new_n402), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT101), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n522), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G99gat), .B(G106gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n530), .B(new_n522), .C1(new_n527), .C2(new_n528), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n488), .B1(new_n520), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(KEYINPUT17), .B(new_n498), .C1(new_n507), .C2(new_n518), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n504), .A2(new_n505), .A3(new_n493), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n505), .B1(new_n504), .B2(new_n493), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n511), .A2(G50gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n509), .A2(G43gat), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n514), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n491), .B1(new_n544), .B2(new_n500), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT89), .B1(new_n510), .B2(new_n512), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n516), .B(new_n499), .C1(new_n546), .C2(new_n508), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n541), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT17), .B1(new_n548), .B2(new_n498), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n538), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT102), .B1(new_n550), .B2(new_n534), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n519), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n553), .A2(KEYINPUT102), .A3(new_n534), .A4(new_n537), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n536), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(G190gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n553), .A2(new_n534), .A3(new_n537), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT102), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n554), .ZN(new_n561));
  INV_X1    g360(.A(G190gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n562), .A3(new_n536), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n557), .A2(G218gat), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(G218gat), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n562), .B1(new_n561), .B2(new_n536), .ZN(new_n566));
  AOI211_X1 g365(.A(G190gat), .B(new_n535), .C1(new_n560), .C2(new_n554), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n564), .A2(new_n568), .A3(KEYINPUT100), .ZN(new_n569));
  XOR2_X1   g368(.A(KEYINPUT98), .B(KEYINPUT99), .Z(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n487), .A2(KEYINPUT41), .ZN(new_n572));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n572), .B(new_n573), .Z(new_n574));
  INV_X1    g373(.A(new_n570), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n564), .A2(new_n568), .A3(KEYINPUT100), .A4(new_n575), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n571), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n574), .B1(new_n571), .B2(new_n576), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n580));
  XOR2_X1   g379(.A(G57gat), .B(G64gat), .Z(new_n581));
  NAND2_X1  g380(.A1(G71gat), .A2(G78gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT9), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G71gat), .ZN(new_n586));
  INV_X1    g385(.A(G78gat), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT93), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT94), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n582), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(KEYINPUT94), .A2(G71gat), .A3(G78gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n588), .A2(new_n591), .A3(new_n592), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n585), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G57gat), .B(G64gat), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT95), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT9), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n597), .A2(new_n598), .B1(new_n582), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n581), .A2(KEYINPUT95), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n596), .A2(new_n602), .A3(KEYINPUT96), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT96), .B1(new_n596), .B2(new_n602), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n580), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n605), .A2(G127gat), .ZN(new_n606));
  INV_X1    g405(.A(G155gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(G127gat), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n607), .B1(new_n606), .B2(new_n608), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(G183gat), .Z(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(G211gat), .Z(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n614), .B1(new_n609), .B2(new_n610), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT21), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n603), .A2(new_n604), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(G8gat), .ZN(new_n621));
  XOR2_X1   g420(.A(G15gat), .B(G22gat), .Z(new_n622));
  INV_X1    g421(.A(G1gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT91), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n623), .A2(KEYINPUT16), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n624), .B1(new_n622), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n626), .B(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n620), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n616), .A2(new_n632), .A3(new_n617), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n533), .A2(KEYINPUT103), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n532), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n596), .A2(new_n602), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n529), .A2(KEYINPUT103), .A3(new_n531), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n534), .B1(new_n604), .B2(new_n603), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT10), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n603), .A2(new_n604), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n650), .A2(KEYINPUT10), .A3(new_n533), .A4(new_n532), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n641), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n640), .B1(new_n646), .B2(new_n647), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n639), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n649), .A2(new_n651), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n653), .B1(new_n655), .B2(new_n640), .ZN(new_n656));
  INV_X1    g455(.A(new_n639), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT104), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n659));
  NOR4_X1   g458(.A1(new_n652), .A2(new_n659), .A3(new_n653), .A4(new_n639), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n654), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g462(.A(KEYINPUT105), .B(new_n654), .C1(new_n658), .C2(new_n660), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n579), .A2(KEYINPUT106), .A3(new_n636), .A4(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n574), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n566), .A2(new_n567), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n669), .B2(G218gat), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n575), .B1(new_n670), .B2(new_n568), .ZN(new_n671));
  INV_X1    g470(.A(new_n576), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n571), .A2(new_n574), .A3(new_n576), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n673), .A2(new_n665), .A3(new_n636), .A4(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n666), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT92), .ZN(new_n679));
  OR3_X1    g478(.A1(new_n629), .A2(new_n679), .A3(new_n519), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n629), .A2(new_n519), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n679), .B1(new_n629), .B2(new_n519), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(G229gat), .A2(G233gat), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT13), .Z(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n553), .A2(new_n537), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n681), .B(new_n684), .C1(new_n687), .C2(new_n629), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT18), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n686), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(G113gat), .B(G141gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G197gat), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT11), .B(G169gat), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT12), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n686), .A2(new_n690), .A3(new_n691), .A4(new_n697), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n486), .A2(new_n678), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n417), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g504(.A(KEYINPUT16), .B(G8gat), .Z(new_n706));
  NAND3_X1  g505(.A1(new_n702), .A2(new_n479), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(KEYINPUT42), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n702), .A2(new_n479), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n710), .B2(G8gat), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n708), .B1(new_n707), .B2(new_n711), .ZN(G1325gat));
  AOI21_X1  g511(.A(G15gat), .B1(new_n702), .B2(new_n362), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n446), .A2(G15gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT107), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n713), .B1(new_n702), .B2(new_n715), .ZN(G1326gat));
  NOR2_X1   g515(.A1(new_n348), .A2(new_n349), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT43), .B(G22gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  NAND2_X1  g519(.A1(new_n673), .A2(new_n674), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n486), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n665), .ZN(new_n723));
  INV_X1    g522(.A(new_n701), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n723), .A2(new_n636), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n489), .A3(new_n703), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT45), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n722), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n486), .A2(new_n721), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n726), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n703), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n729), .B1(new_n489), .B2(new_n737), .ZN(G1328gat));
  NAND3_X1  g537(.A1(new_n727), .A2(new_n490), .A3(new_n479), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT46), .Z(new_n740));
  NAND2_X1  g539(.A1(new_n735), .A2(new_n479), .ZN(new_n741));
  OAI21_X1  g540(.A(G36gat), .B1(new_n741), .B2(KEYINPUT109), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n741), .A2(KEYINPUT109), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n740), .B1(new_n742), .B2(new_n743), .ZN(G1329gat));
  AOI21_X1  g543(.A(new_n511), .B1(new_n735), .B2(new_n446), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n727), .ZN(new_n747));
  INV_X1    g546(.A(new_n362), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n747), .A2(G43gat), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n746), .A2(KEYINPUT47), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n745), .B2(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1330gat));
  AOI21_X1  g553(.A(new_n509), .B1(new_n735), .B2(new_n717), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n717), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n747), .A2(G50gat), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n756), .A2(KEYINPUT48), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT48), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n755), .B2(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(G1331gat));
  NAND3_X1  g562(.A1(new_n579), .A2(new_n636), .A3(new_n724), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n665), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n486), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n703), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g568(.A(new_n439), .B(new_n766), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n770));
  NOR2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1333gat));
  INV_X1    g571(.A(new_n446), .ZN(new_n773));
  OAI21_X1  g572(.A(G71gat), .B1(new_n766), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n362), .A2(new_n586), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n766), .B2(new_n775), .ZN(new_n776));
  XOR2_X1   g575(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1334gat));
  NOR2_X1   g577(.A1(new_n766), .A2(new_n757), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(new_n587), .ZN(G1335gat));
  NOR2_X1   g579(.A1(new_n636), .A2(new_n701), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n486), .A2(new_n721), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n486), .A2(KEYINPUT51), .A3(new_n721), .A4(new_n781), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(new_n703), .A3(new_n723), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n723), .A2(new_n781), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n788), .B1(new_n732), .B2(new_n734), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n417), .A2(new_n402), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n787), .A2(new_n402), .B1(new_n789), .B2(new_n790), .ZN(G1336gat));
  NOR3_X1   g590(.A1(new_n665), .A2(new_n636), .A3(new_n701), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n486), .A2(new_n721), .A3(new_n733), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n730), .B1(new_n486), .B2(new_n721), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n479), .B(new_n792), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G92gat), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n439), .A2(G92gat), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n786), .A2(new_n723), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n801), .A3(KEYINPUT52), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n796), .B(new_n798), .C1(new_n800), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1337gat));
  NAND3_X1  g604(.A1(new_n786), .A2(new_n362), .A3(new_n723), .ZN(new_n806));
  INV_X1    g605(.A(G99gat), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n773), .A2(new_n807), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n806), .A2(new_n807), .B1(new_n789), .B2(new_n808), .ZN(G1338gat));
  NAND2_X1  g608(.A1(new_n789), .A2(new_n717), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G106gat), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n757), .A2(G106gat), .A3(new_n665), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT53), .B1(new_n786), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n812), .B(KEYINPUT112), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n810), .A2(G106gat), .B1(new_n786), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(G1339gat));
  OR2_X1    g617(.A1(new_n764), .A2(new_n723), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n683), .A2(new_n685), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n687), .A2(new_n629), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n684), .B1(new_n821), .B2(new_n681), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n696), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n700), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n652), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n640), .B2(new_n655), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n657), .B1(new_n652), .B2(new_n827), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n826), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(new_n826), .A3(new_n830), .ZN(new_n833));
  INV_X1    g632(.A(new_n658), .ZN(new_n834));
  INV_X1    g633(.A(new_n660), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n832), .A2(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n721), .A2(new_n825), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n834), .A2(new_n835), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n829), .A2(new_n826), .A3(new_n830), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n701), .B(new_n838), .C1(new_n839), .C2(new_n831), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n824), .B1(new_n663), .B2(new_n664), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n674), .B(new_n673), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n837), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n636), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n417), .B1(new_n819), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n717), .A2(new_n748), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n847), .A2(new_n439), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(G113gat), .B1(new_n849), .B2(new_n724), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n757), .A2(new_n278), .A3(new_n439), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n701), .A2(new_n250), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  XOR2_X1   g653(.A(new_n854), .B(KEYINPUT113), .Z(G1340gat));
  OAI21_X1  g654(.A(G120gat), .B1(new_n849), .B2(new_n665), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n665), .A2(new_n252), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n852), .B2(new_n857), .ZN(G1341gat));
  INV_X1    g657(.A(G127gat), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n849), .A2(new_n859), .A3(new_n845), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n847), .A2(new_n636), .A3(new_n851), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n859), .B2(new_n861), .ZN(G1342gat));
  OR2_X1    g661(.A1(new_n579), .A2(new_n247), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n852), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT114), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n849), .B2(new_n579), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(G1343gat));
  NAND2_X1  g668(.A1(new_n819), .A2(new_n846), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n446), .A2(new_n417), .A3(new_n479), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n717), .A3(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(G141gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n701), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n875), .A2(KEYINPUT115), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT58), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT116), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n870), .B2(new_n717), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n764), .A2(new_n723), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n636), .B1(new_n837), .B2(new_n843), .ZN(new_n881));
  OAI211_X1 g680(.A(KEYINPUT57), .B(new_n717), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n701), .B(new_n871), .C1(new_n879), .C2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G141gat), .ZN(new_n885));
  INV_X1    g684(.A(new_n875), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n878), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI211_X1 g686(.A(KEYINPUT116), .B(new_n875), .C1(new_n884), .C2(G141gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n877), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n871), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n717), .B1(new_n880), .B2(new_n881), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n890), .B1(new_n893), .B2(new_n882), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n873), .B1(new_n894), .B2(new_n701), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT116), .B1(new_n895), .B2(new_n875), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n885), .A2(new_n878), .A3(new_n886), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n896), .A2(new_n897), .A3(KEYINPUT58), .A4(new_n876), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n889), .A2(new_n898), .ZN(G1344gat));
  INV_X1    g698(.A(new_n872), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n282), .A3(new_n723), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n903), .B(new_n836), .C1(new_n577), .C2(new_n578), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n825), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n903), .B1(new_n721), .B2(new_n836), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n843), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n907), .A2(new_n845), .B1(new_n678), .B2(new_n724), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT118), .B(new_n892), .C1(new_n908), .C2(new_n757), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n882), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n836), .B1(new_n577), .B2(new_n578), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT117), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n825), .A3(new_n904), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n636), .B1(new_n913), .B2(new_n843), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n701), .B1(new_n666), .B2(new_n677), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n717), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT118), .B1(new_n916), .B2(new_n892), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n723), .B(new_n871), .C1(new_n910), .C2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n902), .B1(new_n918), .B2(G148gat), .ZN(new_n919));
  AOI211_X1 g718(.A(KEYINPUT59), .B(new_n282), .C1(new_n894), .C2(new_n723), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n901), .B1(new_n919), .B2(new_n920), .ZN(G1345gat));
  AOI21_X1  g720(.A(G155gat), .B1(new_n900), .B2(new_n636), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n845), .A2(new_n607), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n922), .B1(new_n894), .B2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT119), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n924), .B(new_n925), .ZN(G1346gat));
  INV_X1    g725(.A(G162gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n900), .A2(new_n927), .A3(new_n721), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT120), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n894), .A2(new_n721), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(new_n927), .ZN(G1347gat));
  NOR2_X1   g730(.A1(new_n703), .A2(new_n439), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n870), .A2(new_n848), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G169gat), .B1(new_n933), .B2(new_n724), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n870), .A2(new_n757), .A3(new_n278), .A4(new_n932), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n724), .A2(G169gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n937), .B(KEYINPUT121), .Z(G1348gat));
  INV_X1    g737(.A(G176gat), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n933), .A2(new_n939), .A3(new_n665), .ZN(new_n940));
  INV_X1    g739(.A(new_n935), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n723), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n940), .B1(new_n942), .B2(new_n939), .ZN(G1349gat));
  NOR2_X1   g742(.A1(new_n845), .A2(new_n230), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT123), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n933), .A2(new_n946), .A3(new_n845), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n933), .B2(new_n845), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n224), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g750(.A(G190gat), .B1(new_n933), .B2(new_n579), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT61), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n941), .A2(new_n562), .A3(new_n721), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1351gat));
  AND2_X1   g754(.A1(new_n870), .A2(new_n932), .ZN(new_n956));
  INV_X1    g755(.A(new_n366), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n958), .A2(G197gat), .A3(new_n724), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n932), .A2(new_n773), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n701), .B(new_n963), .C1(new_n910), .C2(new_n917), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n964), .A2(KEYINPUT125), .ZN(new_n965));
  OAI21_X1  g764(.A(G197gat), .B1(new_n964), .B2(KEYINPUT125), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n961), .B1(new_n965), .B2(new_n966), .ZN(G1352gat));
  OAI211_X1 g766(.A(new_n723), .B(new_n963), .C1(new_n910), .C2(new_n917), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g769(.A(KEYINPUT126), .B(G204gat), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT118), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n907), .A2(new_n845), .ZN(new_n973));
  INV_X1    g772(.A(new_n915), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n757), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n975), .B2(KEYINPUT57), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n976), .A2(new_n882), .A3(new_n909), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n977), .A2(KEYINPUT127), .A3(new_n723), .A4(new_n963), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n970), .A2(new_n971), .A3(new_n978), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n958), .A2(new_n665), .A3(new_n971), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n979), .A2(new_n981), .ZN(G1353gat));
  OR3_X1    g781(.A1(new_n958), .A2(G211gat), .A3(new_n845), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n636), .B(new_n963), .C1(new_n910), .C2(new_n917), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n984), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT63), .B1(new_n984), .B2(G211gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(G1354gat));
  INV_X1    g786(.A(new_n958), .ZN(new_n988));
  AOI21_X1  g787(.A(G218gat), .B1(new_n988), .B2(new_n721), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n977), .A2(new_n963), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n579), .A2(new_n565), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(G1355gat));
endmodule


