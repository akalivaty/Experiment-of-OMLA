

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U553 ( .A(n664), .ZN(n649) );
  NOR2_X1 U554 ( .A1(n569), .A2(n530), .ZN(n787) );
  OR2_X1 U555 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X2 U556 ( .A1(n711), .A2(n713), .ZN(n664) );
  AND2_X2 U557 ( .A1(n580), .A2(G2104), .ZN(n883) );
  NOR2_X1 U558 ( .A1(G164), .A2(G1384), .ZN(n713) );
  XNOR2_X1 U559 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U560 ( .A(KEYINPUT5), .B(KEYINPUT75), .ZN(n533) );
  NAND2_X1 U561 ( .A1(n885), .A2(G138), .ZN(n545) );
  NOR2_X1 U562 ( .A1(n693), .A2(n692), .ZN(n694) );
  INV_X1 U563 ( .A(G2105), .ZN(n580) );
  NOR2_X1 U564 ( .A1(n605), .A2(n518), .ZN(n606) );
  NAND2_X1 U565 ( .A1(n743), .A2(n521), .ZN(n758) );
  XNOR2_X1 U566 ( .A(n537), .B(KEYINPUT76), .ZN(n538) );
  NOR2_X1 U567 ( .A1(n550), .A2(n549), .ZN(G164) );
  XNOR2_X1 U568 ( .A(n543), .B(n542), .ZN(n544) );
  AND2_X1 U569 ( .A1(n783), .A2(G43), .ZN(n518) );
  XOR2_X1 U570 ( .A(n599), .B(KEYINPUT71), .Z(n519) );
  XNOR2_X1 U571 ( .A(KEYINPUT98), .B(n757), .ZN(n520) );
  AND2_X1 U572 ( .A1(n744), .A2(n742), .ZN(n521) );
  OR2_X1 U573 ( .A1(n709), .A2(n708), .ZN(n522) );
  OR2_X1 U574 ( .A1(KEYINPUT33), .A2(n689), .ZN(n523) );
  INV_X1 U575 ( .A(KEYINPUT88), .ZN(n607) );
  XNOR2_X1 U576 ( .A(n608), .B(n607), .ZN(n609) );
  NOR2_X1 U577 ( .A1(n639), .A2(n968), .ZN(n620) );
  AND2_X1 U578 ( .A1(n644), .A2(n643), .ZN(n645) );
  INV_X1 U579 ( .A(KEYINPUT29), .ZN(n647) );
  NOR2_X1 U580 ( .A1(n659), .A2(n658), .ZN(n660) );
  INV_X1 U581 ( .A(KEYINPUT91), .ZN(n670) );
  INV_X1 U582 ( .A(n973), .ZN(n692) );
  XNOR2_X1 U583 ( .A(n705), .B(KEYINPUT95), .ZN(n710) );
  INV_X1 U584 ( .A(KEYINPUT17), .ZN(n540) );
  INV_X1 U585 ( .A(KEYINPUT81), .ZN(n542) );
  NOR2_X2 U586 ( .A1(G651), .A2(G543), .ZN(n788) );
  INV_X1 U587 ( .A(KEYINPUT7), .ZN(n537) );
  NAND2_X1 U588 ( .A1(n758), .A2(n520), .ZN(n759) );
  NAND2_X1 U589 ( .A1(n519), .A2(n606), .ZN(n977) );
  XNOR2_X1 U590 ( .A(n759), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U591 ( .A(n539), .B(n538), .ZN(G168) );
  XOR2_X1 U592 ( .A(G543), .B(KEYINPUT0), .Z(n569) );
  NOR2_X2 U593 ( .A1(G651), .A2(n569), .ZN(n783) );
  NAND2_X1 U594 ( .A1(G51), .A2(n783), .ZN(n526) );
  INV_X1 U595 ( .A(G651), .ZN(n530) );
  NOR2_X1 U596 ( .A1(G543), .A2(n530), .ZN(n524) );
  XOR2_X2 U597 ( .A(KEYINPUT1), .B(n524), .Z(n784) );
  NAND2_X1 U598 ( .A1(G63), .A2(n784), .ZN(n525) );
  NAND2_X1 U599 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U600 ( .A(KEYINPUT6), .B(n527), .ZN(n536) );
  NAND2_X1 U601 ( .A1(G89), .A2(n788), .ZN(n528) );
  XNOR2_X1 U602 ( .A(n528), .B(KEYINPUT74), .ZN(n529) );
  XNOR2_X1 U603 ( .A(n529), .B(KEYINPUT4), .ZN(n532) );
  NAND2_X1 U604 ( .A1(G76), .A2(n787), .ZN(n531) );
  NAND2_X1 U605 ( .A1(n532), .A2(n531), .ZN(n534) );
  NOR2_X1 U606 ( .A1(n536), .A2(n535), .ZN(n539) );
  NOR2_X1 U607 ( .A1(G2104), .A2(G2105), .ZN(n541) );
  XNOR2_X2 U608 ( .A(n541), .B(n540), .ZN(n885) );
  NAND2_X1 U609 ( .A1(G102), .A2(n883), .ZN(n543) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n550) );
  NOR2_X1 U611 ( .A1(G2104), .A2(n580), .ZN(n891) );
  NAND2_X1 U612 ( .A1(n891), .A2(G126), .ZN(n548) );
  NAND2_X1 U613 ( .A1(G2105), .A2(G2104), .ZN(n546) );
  XOR2_X1 U614 ( .A(KEYINPUT66), .B(n546), .Z(n714) );
  NAND2_X1 U615 ( .A1(G114), .A2(n714), .ZN(n547) );
  NAND2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U617 ( .A1(G52), .A2(n783), .ZN(n552) );
  NAND2_X1 U618 ( .A1(G64), .A2(n784), .ZN(n551) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n557) );
  NAND2_X1 U620 ( .A1(G77), .A2(n787), .ZN(n554) );
  NAND2_X1 U621 ( .A1(G90), .A2(n788), .ZN(n553) );
  NAND2_X1 U622 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U623 ( .A(KEYINPUT9), .B(n555), .Z(n556) );
  NOR2_X1 U624 ( .A1(n557), .A2(n556), .ZN(G171) );
  XNOR2_X1 U625 ( .A(KEYINPUT77), .B(KEYINPUT8), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n558), .B(G168), .ZN(G286) );
  NAND2_X1 U627 ( .A1(G75), .A2(n787), .ZN(n560) );
  NAND2_X1 U628 ( .A1(G88), .A2(n788), .ZN(n559) );
  NAND2_X1 U629 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U630 ( .A(KEYINPUT78), .B(n561), .ZN(n565) );
  NAND2_X1 U631 ( .A1(G50), .A2(n783), .ZN(n563) );
  NAND2_X1 U632 ( .A1(G62), .A2(n784), .ZN(n562) );
  NAND2_X1 U633 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U634 ( .A1(n565), .A2(n564), .ZN(G166) );
  INV_X1 U635 ( .A(G166), .ZN(G303) );
  NAND2_X1 U636 ( .A1(G49), .A2(n783), .ZN(n567) );
  NAND2_X1 U637 ( .A1(G74), .A2(G651), .ZN(n566) );
  NAND2_X1 U638 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U639 ( .A1(n784), .A2(n568), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n569), .A2(G87), .ZN(n570) );
  NAND2_X1 U641 ( .A1(n571), .A2(n570), .ZN(G288) );
  NAND2_X1 U642 ( .A1(G48), .A2(n783), .ZN(n573) );
  NAND2_X1 U643 ( .A1(G61), .A2(n784), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U645 ( .A1(G73), .A2(n787), .ZN(n574) );
  XOR2_X1 U646 ( .A(KEYINPUT2), .B(n574), .Z(n575) );
  NOR2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n788), .A2(G86), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n578), .A2(n577), .ZN(G305) );
  NAND2_X1 U650 ( .A1(G137), .A2(n885), .ZN(n584) );
  AND2_X1 U651 ( .A1(G2104), .A2(G101), .ZN(n579) );
  NAND2_X1 U652 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U653 ( .A(n581), .B(KEYINPUT65), .ZN(n582) );
  XNOR2_X1 U654 ( .A(n582), .B(KEYINPUT23), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n891), .A2(G125), .ZN(n586) );
  NAND2_X1 U657 ( .A1(G113), .A2(n714), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U659 ( .A1(n588), .A2(n587), .ZN(G160) );
  NAND2_X1 U660 ( .A1(G85), .A2(n788), .ZN(n590) );
  NAND2_X1 U661 ( .A1(G47), .A2(n783), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U663 ( .A1(G72), .A2(n787), .ZN(n591) );
  XNOR2_X1 U664 ( .A(KEYINPUT67), .B(n591), .ZN(n592) );
  NOR2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n784), .A2(G60), .ZN(n594) );
  NAND2_X1 U667 ( .A1(n595), .A2(n594), .ZN(G290) );
  AND2_X1 U668 ( .A1(G160), .A2(G40), .ZN(n711) );
  NAND2_X1 U669 ( .A1(n649), .A2(G1996), .ZN(n597) );
  XNOR2_X1 U670 ( .A(KEYINPUT26), .B(n597), .ZN(n611) );
  NAND2_X1 U671 ( .A1(G56), .A2(n784), .ZN(n598) );
  XNOR2_X1 U672 ( .A(n598), .B(KEYINPUT14), .ZN(n599) );
  NAND2_X1 U673 ( .A1(G81), .A2(n788), .ZN(n600) );
  XNOR2_X1 U674 ( .A(n600), .B(KEYINPUT72), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n601), .B(KEYINPUT12), .ZN(n603) );
  NAND2_X1 U676 ( .A1(G68), .A2(n787), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U678 ( .A(KEYINPUT13), .B(n604), .Z(n605) );
  NAND2_X1 U679 ( .A1(n664), .A2(G1341), .ZN(n608) );
  NOR2_X1 U680 ( .A1(n977), .A2(n609), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n611), .A2(n610), .ZN(n639) );
  NAND2_X1 U682 ( .A1(n784), .A2(G66), .ZN(n618) );
  NAND2_X1 U683 ( .A1(G79), .A2(n787), .ZN(n613) );
  NAND2_X1 U684 ( .A1(G92), .A2(n788), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U686 ( .A1(G54), .A2(n783), .ZN(n614) );
  XNOR2_X1 U687 ( .A(KEYINPUT73), .B(n614), .ZN(n615) );
  NOR2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U689 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U690 ( .A(KEYINPUT15), .B(n619), .Z(n968) );
  XNOR2_X1 U691 ( .A(n620), .B(KEYINPUT89), .ZN(n634) );
  NOR2_X1 U692 ( .A1(G2067), .A2(n664), .ZN(n622) );
  NOR2_X1 U693 ( .A1(n649), .A2(G1348), .ZN(n621) );
  NOR2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n632) );
  NAND2_X1 U695 ( .A1(n649), .A2(G2072), .ZN(n623) );
  XNOR2_X1 U696 ( .A(n623), .B(KEYINPUT27), .ZN(n625) );
  AND2_X1 U697 ( .A1(G1956), .A2(n664), .ZN(n624) );
  NOR2_X1 U698 ( .A1(n625), .A2(n624), .ZN(n635) );
  NAND2_X1 U699 ( .A1(G53), .A2(n783), .ZN(n627) );
  NAND2_X1 U700 ( .A1(G65), .A2(n784), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U702 ( .A1(G78), .A2(n787), .ZN(n629) );
  NAND2_X1 U703 ( .A1(G91), .A2(n788), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n980) );
  NAND2_X1 U706 ( .A1(n635), .A2(n980), .ZN(n640) );
  AND2_X1 U707 ( .A1(n632), .A2(n640), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n646) );
  NOR2_X1 U709 ( .A1(n635), .A2(n980), .ZN(n638) );
  XNOR2_X1 U710 ( .A(KEYINPUT28), .B(KEYINPUT87), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n636), .B(KEYINPUT86), .ZN(n637) );
  XNOR2_X1 U712 ( .A(n638), .B(n637), .ZN(n644) );
  NAND2_X1 U713 ( .A1(n639), .A2(n968), .ZN(n642) );
  INV_X1 U714 ( .A(n640), .ZN(n641) );
  NAND2_X1 U715 ( .A1(n646), .A2(n645), .ZN(n648) );
  XNOR2_X1 U716 ( .A(n648), .B(n647), .ZN(n653) );
  XNOR2_X1 U717 ( .A(G1961), .B(KEYINPUT85), .ZN(n995) );
  NAND2_X1 U718 ( .A1(n664), .A2(n995), .ZN(n651) );
  XNOR2_X1 U719 ( .A(G2078), .B(KEYINPUT25), .ZN(n946) );
  NAND2_X1 U720 ( .A1(n649), .A2(n946), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n657) );
  NAND2_X1 U722 ( .A1(n657), .A2(G171), .ZN(n652) );
  NAND2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n662) );
  NAND2_X1 U724 ( .A1(G8), .A2(n664), .ZN(n709) );
  NOR2_X1 U725 ( .A1(G1966), .A2(n709), .ZN(n677) );
  NOR2_X1 U726 ( .A1(G2084), .A2(n664), .ZN(n674) );
  NOR2_X1 U727 ( .A1(n677), .A2(n674), .ZN(n654) );
  NAND2_X1 U728 ( .A1(G8), .A2(n654), .ZN(n655) );
  XNOR2_X1 U729 ( .A(KEYINPUT30), .B(n655), .ZN(n656) );
  NOR2_X1 U730 ( .A1(G168), .A2(n656), .ZN(n659) );
  NOR2_X1 U731 ( .A1(G171), .A2(n657), .ZN(n658) );
  XOR2_X1 U732 ( .A(KEYINPUT31), .B(n660), .Z(n661) );
  NAND2_X1 U733 ( .A1(n662), .A2(n661), .ZN(n675) );
  NAND2_X1 U734 ( .A1(n675), .A2(G286), .ZN(n663) );
  XNOR2_X1 U735 ( .A(n663), .B(KEYINPUT90), .ZN(n669) );
  NOR2_X1 U736 ( .A1(G1971), .A2(n709), .ZN(n666) );
  NOR2_X1 U737 ( .A1(G2090), .A2(n664), .ZN(n665) );
  NOR2_X1 U738 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U739 ( .A1(n667), .A2(G303), .ZN(n668) );
  NAND2_X1 U740 ( .A1(n669), .A2(n668), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U742 ( .A1(n672), .A2(G8), .ZN(n673) );
  XNOR2_X1 U743 ( .A(KEYINPUT32), .B(n673), .ZN(n697) );
  NAND2_X1 U744 ( .A1(G8), .A2(n674), .ZN(n679) );
  INV_X1 U745 ( .A(n675), .ZN(n676) );
  NOR2_X1 U746 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U747 ( .A1(n679), .A2(n678), .ZN(n698) );
  INV_X1 U748 ( .A(n709), .ZN(n681) );
  NAND2_X1 U749 ( .A1(G288), .A2(G1976), .ZN(n680) );
  XNOR2_X1 U750 ( .A(n680), .B(KEYINPUT92), .ZN(n982) );
  AND2_X1 U751 ( .A1(n681), .A2(n982), .ZN(n683) );
  AND2_X1 U752 ( .A1(n698), .A2(n683), .ZN(n682) );
  NAND2_X1 U753 ( .A1(n697), .A2(n682), .ZN(n687) );
  INV_X1 U754 ( .A(n683), .ZN(n685) );
  NOR2_X1 U755 ( .A1(G1976), .A2(G288), .ZN(n690) );
  NOR2_X1 U756 ( .A1(G1971), .A2(G303), .ZN(n684) );
  NOR2_X1 U757 ( .A1(n690), .A2(n684), .ZN(n981) );
  OR2_X1 U758 ( .A1(n685), .A2(n981), .ZN(n686) );
  NAND2_X1 U759 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U760 ( .A(n688), .B(KEYINPUT64), .ZN(n689) );
  NAND2_X1 U761 ( .A1(n690), .A2(KEYINPUT33), .ZN(n691) );
  NOR2_X1 U762 ( .A1(n691), .A2(n709), .ZN(n693) );
  XOR2_X1 U763 ( .A(G1981), .B(G305), .Z(n973) );
  NAND2_X1 U764 ( .A1(n523), .A2(n694), .ZN(n704) );
  NAND2_X1 U765 ( .A1(G8), .A2(G166), .ZN(n695) );
  NOR2_X1 U766 ( .A1(G2090), .A2(n695), .ZN(n696) );
  XNOR2_X1 U767 ( .A(n696), .B(KEYINPUT93), .ZN(n700) );
  NAND2_X1 U768 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U769 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U770 ( .A1(n701), .A2(n709), .ZN(n702) );
  XNOR2_X1 U771 ( .A(n702), .B(KEYINPUT94), .ZN(n703) );
  NAND2_X1 U772 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U773 ( .A1(G1981), .A2(G305), .ZN(n706) );
  XOR2_X1 U774 ( .A(n706), .B(KEYINPUT24), .Z(n707) );
  XNOR2_X1 U775 ( .A(KEYINPUT84), .B(n707), .ZN(n708) );
  NAND2_X1 U776 ( .A1(n710), .A2(n522), .ZN(n743) );
  INV_X1 U777 ( .A(n711), .ZN(n712) );
  NOR2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n756) );
  NAND2_X1 U779 ( .A1(G141), .A2(n885), .ZN(n716) );
  BUF_X1 U780 ( .A(n714), .Z(n889) );
  NAND2_X1 U781 ( .A1(G117), .A2(n889), .ZN(n715) );
  NAND2_X1 U782 ( .A1(n716), .A2(n715), .ZN(n719) );
  NAND2_X1 U783 ( .A1(n883), .A2(G105), .ZN(n717) );
  XOR2_X1 U784 ( .A(KEYINPUT38), .B(n717), .Z(n718) );
  NOR2_X1 U785 ( .A1(n719), .A2(n718), .ZN(n721) );
  NAND2_X1 U786 ( .A1(n891), .A2(G129), .ZN(n720) );
  NAND2_X1 U787 ( .A1(n721), .A2(n720), .ZN(n870) );
  NAND2_X1 U788 ( .A1(G1996), .A2(n870), .ZN(n730) );
  NAND2_X1 U789 ( .A1(G131), .A2(n885), .ZN(n723) );
  NAND2_X1 U790 ( .A1(G107), .A2(n889), .ZN(n722) );
  NAND2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n726) );
  NAND2_X1 U792 ( .A1(G95), .A2(n883), .ZN(n724) );
  XNOR2_X1 U793 ( .A(KEYINPUT83), .B(n724), .ZN(n725) );
  NOR2_X1 U794 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U795 ( .A1(n891), .A2(G119), .ZN(n727) );
  NAND2_X1 U796 ( .A1(n728), .A2(n727), .ZN(n882) );
  NAND2_X1 U797 ( .A1(G1991), .A2(n882), .ZN(n729) );
  NAND2_X1 U798 ( .A1(n730), .A2(n729), .ZN(n937) );
  NAND2_X1 U799 ( .A1(n756), .A2(n937), .ZN(n744) );
  XOR2_X1 U800 ( .A(G1986), .B(G290), .Z(n979) );
  XNOR2_X1 U801 ( .A(G2067), .B(KEYINPUT37), .ZN(n753) );
  NAND2_X1 U802 ( .A1(G104), .A2(n883), .ZN(n732) );
  NAND2_X1 U803 ( .A1(G140), .A2(n885), .ZN(n731) );
  NAND2_X1 U804 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U805 ( .A(KEYINPUT34), .B(n733), .ZN(n739) );
  NAND2_X1 U806 ( .A1(n891), .A2(G128), .ZN(n735) );
  NAND2_X1 U807 ( .A1(G116), .A2(n889), .ZN(n734) );
  NAND2_X1 U808 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U809 ( .A(KEYINPUT82), .B(n736), .Z(n737) );
  XNOR2_X1 U810 ( .A(KEYINPUT35), .B(n737), .ZN(n738) );
  NOR2_X1 U811 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U812 ( .A(KEYINPUT36), .B(n740), .ZN(n898) );
  OR2_X1 U813 ( .A1(n753), .A2(n898), .ZN(n922) );
  NAND2_X1 U814 ( .A1(n979), .A2(n922), .ZN(n741) );
  NAND2_X1 U815 ( .A1(n756), .A2(n741), .ZN(n742) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n870), .ZN(n920) );
  INV_X1 U817 ( .A(n744), .ZN(n748) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n746) );
  NOR2_X1 U819 ( .A1(n882), .A2(G1991), .ZN(n745) );
  XNOR2_X1 U820 ( .A(n745), .B(KEYINPUT96), .ZN(n933) );
  NOR2_X1 U821 ( .A1(n746), .A2(n933), .ZN(n747) );
  NOR2_X1 U822 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U823 ( .A(KEYINPUT97), .B(n749), .Z(n750) );
  NOR2_X1 U824 ( .A1(n920), .A2(n750), .ZN(n751) );
  XNOR2_X1 U825 ( .A(n751), .B(KEYINPUT39), .ZN(n752) );
  NAND2_X1 U826 ( .A1(n752), .A2(n922), .ZN(n754) );
  NAND2_X1 U827 ( .A1(n753), .A2(n898), .ZN(n928) );
  NAND2_X1 U828 ( .A1(n754), .A2(n928), .ZN(n755) );
  NAND2_X1 U829 ( .A1(n756), .A2(n755), .ZN(n757) );
  AND2_X1 U830 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U831 ( .A1(G135), .A2(n885), .ZN(n761) );
  NAND2_X1 U832 ( .A1(G111), .A2(n889), .ZN(n760) );
  NAND2_X1 U833 ( .A1(n761), .A2(n760), .ZN(n764) );
  NAND2_X1 U834 ( .A1(n891), .A2(G123), .ZN(n762) );
  XOR2_X1 U835 ( .A(KEYINPUT18), .B(n762), .Z(n763) );
  NOR2_X1 U836 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U837 ( .A1(n883), .A2(G99), .ZN(n765) );
  NAND2_X1 U838 ( .A1(n766), .A2(n765), .ZN(n934) );
  XNOR2_X1 U839 ( .A(G2096), .B(n934), .ZN(n767) );
  OR2_X1 U840 ( .A1(G2100), .A2(n767), .ZN(G156) );
  INV_X1 U841 ( .A(G57), .ZN(G237) );
  INV_X1 U842 ( .A(G132), .ZN(G219) );
  NAND2_X1 U843 ( .A1(G7), .A2(G661), .ZN(n768) );
  XNOR2_X1 U844 ( .A(n768), .B(KEYINPUT70), .ZN(n769) );
  XNOR2_X1 U845 ( .A(KEYINPUT10), .B(n769), .ZN(G223) );
  INV_X1 U846 ( .A(G223), .ZN(n820) );
  NAND2_X1 U847 ( .A1(n820), .A2(G567), .ZN(n770) );
  XOR2_X1 U848 ( .A(KEYINPUT11), .B(n770), .Z(G234) );
  INV_X1 U849 ( .A(G860), .ZN(n775) );
  OR2_X1 U850 ( .A1(n977), .A2(n775), .ZN(G153) );
  INV_X1 U851 ( .A(G171), .ZN(G301) );
  NAND2_X1 U852 ( .A1(G868), .A2(G301), .ZN(n772) );
  INV_X1 U853 ( .A(G868), .ZN(n803) );
  NAND2_X1 U854 ( .A1(n968), .A2(n803), .ZN(n771) );
  NAND2_X1 U855 ( .A1(n772), .A2(n771), .ZN(G284) );
  XOR2_X1 U856 ( .A(n980), .B(KEYINPUT68), .Z(G299) );
  NAND2_X1 U857 ( .A1(G868), .A2(G286), .ZN(n774) );
  NAND2_X1 U858 ( .A1(G299), .A2(n803), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n774), .A2(n773), .ZN(G297) );
  NAND2_X1 U860 ( .A1(n775), .A2(G559), .ZN(n776) );
  INV_X1 U861 ( .A(n968), .ZN(n781) );
  NAND2_X1 U862 ( .A1(n776), .A2(n781), .ZN(n777) );
  XNOR2_X1 U863 ( .A(n777), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U864 ( .A1(G868), .A2(n977), .ZN(n780) );
  NAND2_X1 U865 ( .A1(G868), .A2(n781), .ZN(n778) );
  NOR2_X1 U866 ( .A1(G559), .A2(n778), .ZN(n779) );
  NOR2_X1 U867 ( .A1(n780), .A2(n779), .ZN(G282) );
  NAND2_X1 U868 ( .A1(n781), .A2(G559), .ZN(n801) );
  XNOR2_X1 U869 ( .A(n977), .B(n801), .ZN(n782) );
  NOR2_X1 U870 ( .A1(n782), .A2(G860), .ZN(n793) );
  NAND2_X1 U871 ( .A1(G55), .A2(n783), .ZN(n786) );
  NAND2_X1 U872 ( .A1(G67), .A2(n784), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n786), .A2(n785), .ZN(n792) );
  NAND2_X1 U874 ( .A1(G80), .A2(n787), .ZN(n790) );
  NAND2_X1 U875 ( .A1(G93), .A2(n788), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U877 ( .A1(n792), .A2(n791), .ZN(n804) );
  XNOR2_X1 U878 ( .A(n793), .B(n804), .ZN(G145) );
  XNOR2_X1 U879 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n795) );
  XNOR2_X1 U880 ( .A(G288), .B(G166), .ZN(n794) );
  XNOR2_X1 U881 ( .A(n795), .B(n794), .ZN(n798) );
  XNOR2_X1 U882 ( .A(G299), .B(n977), .ZN(n796) );
  XNOR2_X1 U883 ( .A(n796), .B(G290), .ZN(n797) );
  XNOR2_X1 U884 ( .A(n798), .B(n797), .ZN(n800) );
  XNOR2_X1 U885 ( .A(G305), .B(n804), .ZN(n799) );
  XNOR2_X1 U886 ( .A(n800), .B(n799), .ZN(n906) );
  XOR2_X1 U887 ( .A(n906), .B(n801), .Z(n802) );
  NAND2_X1 U888 ( .A1(G868), .A2(n802), .ZN(n806) );
  NAND2_X1 U889 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U890 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U891 ( .A(KEYINPUT80), .B(n807), .Z(G295) );
  NAND2_X1 U892 ( .A1(G2078), .A2(G2084), .ZN(n808) );
  XOR2_X1 U893 ( .A(KEYINPUT20), .B(n808), .Z(n809) );
  NAND2_X1 U894 ( .A1(G2090), .A2(n809), .ZN(n810) );
  XNOR2_X1 U895 ( .A(KEYINPUT21), .B(n810), .ZN(n811) );
  NAND2_X1 U896 ( .A1(n811), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U897 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U898 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  NOR2_X1 U899 ( .A1(G219), .A2(G220), .ZN(n812) );
  XOR2_X1 U900 ( .A(KEYINPUT22), .B(n812), .Z(n813) );
  NOR2_X1 U901 ( .A1(G218), .A2(n813), .ZN(n814) );
  NAND2_X1 U902 ( .A1(G96), .A2(n814), .ZN(n827) );
  NAND2_X1 U903 ( .A1(n827), .A2(G2106), .ZN(n818) );
  NAND2_X1 U904 ( .A1(G69), .A2(G120), .ZN(n815) );
  NOR2_X1 U905 ( .A1(G237), .A2(n815), .ZN(n816) );
  NAND2_X1 U906 ( .A1(G108), .A2(n816), .ZN(n828) );
  NAND2_X1 U907 ( .A1(n828), .A2(G567), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n840) );
  NAND2_X1 U909 ( .A1(G483), .A2(G661), .ZN(n819) );
  NOR2_X1 U910 ( .A1(n840), .A2(n819), .ZN(n826) );
  NAND2_X1 U911 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n820), .ZN(G217) );
  INV_X1 U913 ( .A(G661), .ZN(n822) );
  NAND2_X1 U914 ( .A1(G2), .A2(G15), .ZN(n821) );
  NOR2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U916 ( .A(KEYINPUT102), .B(n823), .Z(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n824) );
  XOR2_X1 U918 ( .A(KEYINPUT103), .B(n824), .Z(n825) );
  NAND2_X1 U919 ( .A1(n826), .A2(n825), .ZN(G188) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  XOR2_X1 U926 ( .A(G2454), .B(G2435), .Z(n830) );
  XNOR2_X1 U927 ( .A(G2438), .B(G2427), .ZN(n829) );
  XNOR2_X1 U928 ( .A(n830), .B(n829), .ZN(n837) );
  XOR2_X1 U929 ( .A(KEYINPUT99), .B(G2446), .Z(n832) );
  XNOR2_X1 U930 ( .A(G2443), .B(G2430), .ZN(n831) );
  XNOR2_X1 U931 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U932 ( .A(n833), .B(G2451), .Z(n835) );
  XNOR2_X1 U933 ( .A(G1341), .B(G1348), .ZN(n834) );
  XNOR2_X1 U934 ( .A(n835), .B(n834), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n838) );
  NAND2_X1 U936 ( .A1(n838), .A2(G14), .ZN(n839) );
  XOR2_X1 U937 ( .A(KEYINPUT100), .B(n839), .Z(n912) );
  XOR2_X1 U938 ( .A(KEYINPUT101), .B(n912), .Z(G401) );
  INV_X1 U939 ( .A(n840), .ZN(G319) );
  XOR2_X1 U940 ( .A(G2096), .B(KEYINPUT43), .Z(n842) );
  XNOR2_X1 U941 ( .A(G2090), .B(G2678), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n843), .B(KEYINPUT42), .Z(n845) );
  XNOR2_X1 U944 ( .A(G2072), .B(G2067), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U946 ( .A(KEYINPUT104), .B(G2100), .Z(n847) );
  XNOR2_X1 U947 ( .A(G2078), .B(G2084), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(G227) );
  XOR2_X1 U950 ( .A(G1986), .B(G1996), .Z(n851) );
  XNOR2_X1 U951 ( .A(G1966), .B(G1961), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U953 ( .A(G1956), .B(G1971), .Z(n853) );
  XNOR2_X1 U954 ( .A(G1981), .B(G1976), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U956 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U957 ( .A(KEYINPUT105), .B(G2474), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n859) );
  XOR2_X1 U959 ( .A(G1991), .B(KEYINPUT41), .Z(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U961 ( .A1(G124), .A2(n891), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G112), .A2(n889), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G100), .A2(n883), .ZN(n864) );
  NAND2_X1 U966 ( .A1(G136), .A2(n885), .ZN(n863) );
  NAND2_X1 U967 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U968 ( .A1(n866), .A2(n865), .ZN(G162) );
  XOR2_X1 U969 ( .A(KEYINPUT107), .B(KEYINPUT111), .Z(n868) );
  XNOR2_X1 U970 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n867) );
  XNOR2_X1 U971 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U972 ( .A(KEYINPUT46), .B(n869), .ZN(n904) );
  XNOR2_X1 U973 ( .A(G164), .B(n870), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n871), .B(n934), .ZN(n902) );
  NAND2_X1 U975 ( .A1(n891), .A2(G130), .ZN(n873) );
  NAND2_X1 U976 ( .A1(G118), .A2(n889), .ZN(n872) );
  NAND2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G106), .A2(n883), .ZN(n875) );
  NAND2_X1 U979 ( .A1(G142), .A2(n885), .ZN(n874) );
  NAND2_X1 U980 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U981 ( .A(KEYINPUT106), .B(n876), .Z(n877) );
  XNOR2_X1 U982 ( .A(KEYINPUT45), .B(n877), .ZN(n878) );
  NOR2_X1 U983 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U984 ( .A(G162), .B(n880), .Z(n881) );
  XNOR2_X1 U985 ( .A(n882), .B(n881), .ZN(n897) );
  NAND2_X1 U986 ( .A1(n883), .A2(G103), .ZN(n884) );
  XNOR2_X1 U987 ( .A(n884), .B(KEYINPUT108), .ZN(n887) );
  NAND2_X1 U988 ( .A1(G139), .A2(n885), .ZN(n886) );
  NAND2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U990 ( .A(KEYINPUT109), .B(n888), .Z(n896) );
  NAND2_X1 U991 ( .A1(G115), .A2(n889), .ZN(n890) );
  XNOR2_X1 U992 ( .A(n890), .B(KEYINPUT110), .ZN(n893) );
  NAND2_X1 U993 ( .A1(G127), .A2(n891), .ZN(n892) );
  NAND2_X1 U994 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U995 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n924) );
  XOR2_X1 U997 ( .A(n897), .B(n924), .Z(n900) );
  XOR2_X1 U998 ( .A(G160), .B(n898), .Z(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U1000 ( .A(n902), .B(n901), .Z(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U1003 ( .A(n906), .B(n968), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n907), .B(G286), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n908), .B(G171), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n909), .ZN(G397) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n910), .B(KEYINPUT49), .ZN(n911) );
  NOR2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n913), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(KEYINPUT113), .B(n914), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1014 ( .A(KEYINPUT114), .B(n917), .Z(G308) );
  INV_X1 U1015 ( .A(G308), .ZN(G225) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1017 ( .A(G2090), .B(G162), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n918), .B(KEYINPUT115), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1020 ( .A(KEYINPUT51), .B(n921), .Z(n923) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n931) );
  XOR2_X1 U1022 ( .A(G2072), .B(n924), .Z(n926) );
  XOR2_X1 U1023 ( .A(G164), .B(G2078), .Z(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(n927), .B(KEYINPUT50), .ZN(n929) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n939) );
  XOR2_X1 U1028 ( .A(G160), .B(G2084), .Z(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n940), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n941), .B(KEYINPUT116), .ZN(n942) );
  NOR2_X1 U1035 ( .A1(KEYINPUT55), .A2(n942), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(KEYINPUT117), .B(n943), .ZN(n944) );
  NAND2_X1 U1037 ( .A1(n944), .A2(G29), .ZN(n1026) );
  XOR2_X1 U1038 ( .A(G29), .B(KEYINPUT120), .Z(n965) );
  XNOR2_X1 U1039 ( .A(G2084), .B(G34), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(n945), .B(KEYINPUT54), .ZN(n962) );
  XOR2_X1 U1041 ( .A(G2090), .B(G35), .Z(n960) );
  XNOR2_X1 U1042 ( .A(G27), .B(n946), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(G1996), .B(G32), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(G26), .B(G2067), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(G33), .B(G2072), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1049 ( .A(KEYINPUT118), .B(n953), .Z(n955) );
  XNOR2_X1 U1050 ( .A(G1991), .B(G25), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n956), .A2(G28), .ZN(n957) );
  XOR2_X1 U1053 ( .A(KEYINPUT119), .B(n957), .Z(n958) );
  XNOR2_X1 U1054 ( .A(n958), .B(KEYINPUT53), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(n963), .B(KEYINPUT55), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n966), .ZN(n1024) );
  XNOR2_X1 U1060 ( .A(G16), .B(KEYINPUT56), .ZN(n994) );
  XNOR2_X1 U1061 ( .A(G171), .B(G1961), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(n967), .B(KEYINPUT122), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(G1348), .B(KEYINPUT121), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(n969), .B(n968), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(G1966), .B(G168), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1068 ( .A(KEYINPUT57), .B(n974), .Z(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n992) );
  XOR2_X1 U1070 ( .A(G1341), .B(n977), .Z(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n990) );
  XOR2_X1 U1072 ( .A(n980), .B(G1956), .Z(n987) );
  AND2_X1 U1073 ( .A1(G303), .A2(G1971), .ZN(n984) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(KEYINPUT123), .B(n985), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1078 ( .A(KEYINPUT124), .B(n988), .Z(n989) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1081 ( .A1(n994), .A2(n993), .ZN(n1022) );
  INV_X1 U1082 ( .A(G16), .ZN(n1020) );
  XNOR2_X1 U1083 ( .A(G5), .B(n995), .ZN(n1015) );
  XNOR2_X1 U1084 ( .A(G1956), .B(G20), .ZN(n1000) );
  XNOR2_X1 U1085 ( .A(G1981), .B(G6), .ZN(n997) );
  XNOR2_X1 U1086 ( .A(G1341), .B(G19), .ZN(n996) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(KEYINPUT125), .B(n998), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(KEYINPUT126), .B(n1001), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G1348), .B(KEYINPUT59), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(G4), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1005), .B(KEYINPUT60), .ZN(n1013) );
  XNOR2_X1 U1095 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n1011) );
  XNOR2_X1 U1096 ( .A(G1976), .B(G23), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(G1971), .B(G22), .ZN(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XOR2_X1 U1099 ( .A(G1986), .B(G24), .Z(n1008) );
  NAND2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1101 ( .A(n1011), .B(n1010), .Z(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(G21), .B(G1966), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

