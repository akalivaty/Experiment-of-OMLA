//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT79), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT3), .A3(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G101), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT75), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n196), .B1(new_n192), .B2(G104), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n190), .A2(KEYINPUT75), .A3(G107), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n194), .A2(new_n195), .A3(new_n197), .A4(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT76), .B1(new_n192), .B2(G104), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT76), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(new_n190), .A3(G107), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n192), .A2(G104), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G101), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT78), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT78), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n199), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G119), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G116), .ZN(new_n211));
  INV_X1    g025(.A(G116), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G119), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT5), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n211), .A2(KEYINPUT5), .ZN(new_n217));
  INV_X1    g031(.A(G113), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT2), .B(G113), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n216), .A2(new_n219), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n207), .A2(new_n209), .A3(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n192), .A2(KEYINPUT3), .A3(G104), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT3), .B1(new_n192), .B2(G104), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n197), .B(new_n198), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G101), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT4), .A3(new_n199), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n215), .A2(new_n221), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n214), .A2(new_n220), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n226), .A2(new_n232), .A3(G101), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n228), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G110), .B(G122), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n223), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G224), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G953), .ZN(new_n238));
  INV_X1    g052(.A(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G143), .ZN(new_n240));
  INV_X1    g054(.A(G143), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n239), .A2(G143), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n243), .A2(new_n244), .B1(KEYINPUT1), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n244), .A2(KEYINPUT1), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(new_n240), .A3(new_n242), .ZN(new_n248));
  AOI21_X1  g062(.A(G125), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G125), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n243), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n240), .A2(new_n242), .A3(new_n251), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n250), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n238), .B1(new_n249), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(new_n255), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G125), .ZN(new_n259));
  INV_X1    g073(.A(new_n238), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n245), .A2(KEYINPUT1), .ZN(new_n261));
  XNOR2_X1  g075(.A(G143), .B(G146), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n248), .B(new_n261), .C1(G128), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n250), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n259), .A2(new_n260), .A3(new_n264), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n257), .B(new_n265), .C1(KEYINPUT7), .C2(new_n238), .ZN(new_n266));
  OR4_X1    g080(.A1(KEYINPUT7), .A2(new_n249), .A3(new_n256), .A4(new_n238), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n236), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT80), .B(KEYINPUT8), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n235), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n223), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n222), .B1(new_n199), .B2(new_n205), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(G902), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n223), .A2(new_n234), .ZN(new_n275));
  INV_X1    g089(.A(new_n235), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(KEYINPUT6), .A3(new_n236), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n257), .A2(new_n265), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n275), .A2(new_n280), .A3(new_n276), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(G210), .B1(G237), .B2(G902), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n274), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n283), .B1(new_n274), .B2(new_n282), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n188), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(G234), .A2(G237), .ZN(new_n287));
  INV_X1    g101(.A(G953), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(G952), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT21), .B(G898), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n287), .A2(G902), .A3(G953), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n289), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n241), .A2(G128), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n244), .A2(G143), .ZN(new_n296));
  INV_X1    g110(.A(G134), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G122), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G116), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n212), .A2(G122), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G107), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n301), .A3(new_n192), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n298), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT13), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n295), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n241), .A2(KEYINPUT13), .A3(G128), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n307), .A2(new_n308), .A3(new_n296), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n305), .B1(new_n297), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n212), .A2(KEYINPUT14), .A3(G122), .ZN(new_n311));
  OAI211_X1 g125(.A(G107), .B(new_n311), .C1(new_n302), .C2(KEYINPUT14), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n297), .B1(new_n295), .B2(new_n296), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n312), .B(new_n304), .C1(new_n298), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT9), .B(G234), .ZN(new_n316));
  INV_X1    g130(.A(G217), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n316), .A2(new_n317), .A3(G953), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n310), .A2(new_n314), .A3(new_n318), .ZN(new_n321));
  AOI21_X1  g135(.A(G902), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G478), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n323), .A2(KEYINPUT15), .ZN(new_n324));
  OR2_X1    g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n324), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G902), .ZN(new_n328));
  OR2_X1    g142(.A1(KEYINPUT82), .A2(G143), .ZN(new_n329));
  NAND2_X1  g143(.A1(KEYINPUT82), .A2(G143), .ZN(new_n330));
  NOR2_X1   g144(.A1(G237), .A2(G953), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n329), .A2(new_n330), .B1(new_n331), .B2(G214), .ZN(new_n332));
  INV_X1    g146(.A(G237), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n288), .A3(G214), .ZN(new_n334));
  NOR2_X1   g148(.A1(KEYINPUT82), .A2(G143), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(G131), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G131), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n329), .A2(G214), .A3(new_n331), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT82), .B(G143), .Z(new_n340));
  INV_X1    g154(.A(new_n334), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n338), .B(new_n339), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT17), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n337), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT87), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G140), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G125), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n250), .A2(G140), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT16), .ZN(new_n350));
  OR3_X1    g164(.A1(new_n250), .A2(KEYINPUT16), .A3(G140), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n350), .A2(G146), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(G146), .B1(new_n350), .B2(new_n351), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n337), .A2(new_n342), .A3(KEYINPUT87), .A4(new_n343), .ZN(new_n355));
  OR2_X1    g169(.A1(new_n337), .A2(new_n343), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n346), .A2(new_n354), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n348), .A2(new_n349), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n239), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n348), .A2(new_n349), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G146), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT83), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(KEYINPUT18), .A3(G131), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n339), .B(new_n364), .C1(new_n340), .C2(new_n341), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(KEYINPUT18), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n362), .B(new_n365), .C1(new_n337), .C2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G113), .B(G122), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(new_n190), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(KEYINPUT86), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n357), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n369), .B1(new_n357), .B2(new_n367), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n328), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT88), .B(G475), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n337), .A2(new_n342), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n350), .A2(new_n351), .A3(G146), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT19), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n348), .B(new_n349), .C1(KEYINPUT84), .C2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n382), .B(new_n239), .C1(new_n358), .C2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n379), .A2(new_n380), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n367), .ZN(new_n386));
  INV_X1    g200(.A(new_n369), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n378), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI211_X1 g202(.A(KEYINPUT85), .B(new_n369), .C1(new_n385), .C2(new_n367), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n371), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n391));
  NOR2_X1   g205(.A1(G475), .A2(G902), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  XOR2_X1   g207(.A(KEYINPUT81), .B(KEYINPUT20), .Z(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(new_n390), .B2(new_n392), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n327), .B(new_n377), .C1(new_n393), .C2(new_n395), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n286), .A2(new_n294), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT29), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT11), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n297), .B2(G137), .ZN(new_n400));
  INV_X1    g214(.A(G137), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT11), .A3(G134), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n297), .A2(G137), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G131), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n400), .A2(new_n402), .A3(new_n338), .A4(new_n403), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n258), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n297), .A2(G137), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n401), .A2(G134), .ZN(new_n410));
  OAI21_X1  g224(.A(G131), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n263), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n408), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT30), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n414), .A2(new_n415), .B1(new_n230), .B2(new_n229), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n412), .A2(KEYINPUT66), .B1(new_n246), .B2(new_n248), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT66), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n406), .A2(new_n411), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n405), .A2(KEYINPUT65), .A3(new_n406), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT65), .B1(new_n405), .B2(new_n406), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OR2_X1    g237(.A1(KEYINPUT0), .A2(G128), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n240), .A2(new_n242), .B1(new_n424), .B2(new_n251), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n240), .A2(new_n242), .A3(new_n251), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT64), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT64), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n252), .A2(new_n253), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n255), .B(new_n428), .C1(new_n429), .C2(new_n262), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(KEYINPUT30), .B(new_n420), .C1(new_n423), .C2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT65), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n407), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n405), .A2(KEYINPUT65), .A3(new_n406), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n431), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n436), .A2(new_n437), .B1(new_n419), .B2(new_n417), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n231), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n229), .A2(KEYINPUT67), .A3(new_n230), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n416), .A2(new_n432), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  XOR2_X1   g257(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n444));
  NAND2_X1  g258(.A1(new_n331), .A2(G210), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n444), .B(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT26), .B(G101), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n446), .B(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n398), .B1(new_n443), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT28), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n442), .B(new_n420), .C1(new_n423), .C2(new_n431), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n414), .A2(new_n231), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT28), .B1(new_n438), .B2(new_n442), .ZN(new_n454));
  INV_X1    g268(.A(new_n448), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n328), .B1(new_n449), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n440), .A2(new_n441), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n431), .B1(new_n435), .B2(new_n434), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n412), .A2(KEYINPUT66), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n460), .A2(new_n419), .A3(new_n263), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n458), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(KEYINPUT69), .A3(new_n451), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT69), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n438), .A2(new_n464), .A3(new_n442), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n463), .A2(KEYINPUT28), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n454), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n455), .A2(new_n398), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(G472), .B1(new_n457), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT32), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n455), .B1(new_n453), .B2(new_n454), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n406), .A2(new_n411), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n407), .A2(new_n258), .B1(new_n473), .B2(new_n263), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n231), .B1(new_n474), .B2(KEYINPUT30), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n438), .B2(KEYINPUT30), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n451), .A2(new_n448), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT31), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n416), .A2(new_n432), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT31), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n479), .A2(new_n480), .A3(new_n451), .A4(new_n448), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n472), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(G472), .A2(G902), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n471), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n482), .A2(new_n471), .A3(new_n483), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n470), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT73), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT23), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(new_n210), .B2(G128), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n244), .A2(KEYINPUT23), .A3(G119), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n210), .A2(G128), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  XOR2_X1   g306(.A(KEYINPUT24), .B(G110), .Z(new_n493));
  XNOR2_X1  g307(.A(G119), .B(G128), .ZN(new_n494));
  OAI22_X1  g308(.A1(new_n492), .A2(G110), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n380), .A3(new_n359), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n493), .A2(new_n494), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n352), .B2(new_n353), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n492), .A2(KEYINPUT70), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT70), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n489), .A2(new_n490), .A3(new_n500), .A4(new_n491), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n499), .A2(G110), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n496), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT71), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n499), .A2(G110), .A3(new_n501), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n505), .B(new_n497), .C1(new_n353), .C2(new_n352), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT71), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(new_n496), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT22), .B(G137), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n288), .A2(G221), .A3(G234), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n504), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n511), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n503), .A2(KEYINPUT71), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n317), .B1(G234), .B2(new_n328), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(G902), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(G902), .B1(new_n512), .B2(new_n514), .ZN(new_n519));
  XOR2_X1   g333(.A(KEYINPUT72), .B(KEYINPUT25), .Z(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  OR2_X1    g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n516), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT25), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n523), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  AOI211_X1 g339(.A(new_n487), .B(new_n518), .C1(new_n522), .C2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n515), .A2(new_n524), .A3(new_n328), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(new_n516), .C1(new_n519), .C2(new_n521), .ZN(new_n528));
  INV_X1    g342(.A(new_n518), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT73), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G221), .ZN(new_n532));
  INV_X1    g346(.A(new_n316), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n532), .B1(new_n533), .B2(new_n328), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n407), .A2(KEYINPUT12), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n263), .B1(new_n207), .B2(new_n209), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n262), .A2(KEYINPUT77), .A3(new_n247), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT77), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n248), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n246), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(new_n199), .A3(new_n205), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n535), .B1(new_n536), .B2(new_n542), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n199), .A2(new_n205), .A3(new_n208), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n208), .B1(new_n199), .B2(new_n205), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n413), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n423), .B1(new_n546), .B2(new_n541), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n543), .B1(new_n547), .B2(KEYINPUT12), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n228), .A2(new_n427), .A3(new_n430), .A4(new_n233), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT10), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n550), .B1(new_n246), .B2(new_n248), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n207), .A2(new_n209), .A3(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n246), .A2(new_n537), .A3(new_n539), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n550), .B1(new_n553), .B2(new_n206), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n549), .A2(new_n552), .A3(new_n423), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n548), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(G110), .B(G140), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT74), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n288), .A2(G227), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n549), .A2(new_n552), .A3(new_n554), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n436), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n555), .A2(new_n560), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n556), .A2(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(G469), .B1(new_n565), .B2(G902), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n563), .A2(new_n555), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n561), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n548), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G469), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n571), .A3(new_n328), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n534), .B1(new_n566), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n397), .A2(new_n486), .A3(new_n531), .A4(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(G101), .ZN(G3));
  OR2_X1    g389(.A1(new_n526), .A2(new_n530), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n482), .A2(new_n483), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G472), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n482), .B2(new_n328), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(G469), .A2(G902), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n556), .A2(new_n561), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n564), .A2(new_n563), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(G469), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n572), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n534), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n576), .A2(new_n582), .A3(new_n589), .ZN(new_n590));
  OR3_X1    g404(.A1(new_n322), .A2(KEYINPUT91), .A3(G478), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT91), .B1(new_n322), .B2(G478), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT33), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n315), .B2(KEYINPUT89), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(new_n321), .A3(new_n320), .ZN(new_n596));
  INV_X1    g410(.A(new_n321), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n318), .B1(new_n310), .B2(new_n314), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT89), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n310), .B2(new_n314), .ZN(new_n600));
  OAI22_X1  g414(.A1(new_n597), .A2(new_n598), .B1(new_n600), .B2(new_n594), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n323), .A2(G902), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n596), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT90), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n593), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n377), .B1(new_n393), .B2(new_n395), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n608), .A3(new_n293), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n187), .B1(new_n284), .B2(new_n285), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n590), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT92), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  AOI22_X1  g429(.A1(new_n374), .A2(new_n376), .B1(new_n325), .B2(new_n326), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n293), .B(KEYINPUT93), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n390), .A2(new_n392), .ZN(new_n618));
  INV_X1    g432(.A(new_n394), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n616), .B(new_n617), .C1(new_n620), .C2(new_n395), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n610), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n590), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT94), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT35), .B(G107), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  NOR2_X1   g440(.A1(new_n511), .A2(KEYINPUT36), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n503), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n517), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n528), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n397), .A2(new_n573), .A3(new_n581), .A4(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT37), .B(G110), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT95), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n631), .B(new_n633), .ZN(G12));
  AND2_X1   g448(.A1(new_n528), .A2(new_n629), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n577), .A2(KEYINPUT32), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n482), .A2(new_n471), .A3(new_n483), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n635), .B1(new_n638), .B2(new_n470), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n289), .B(KEYINPUT96), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n640), .B1(G900), .B2(new_n292), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n616), .B(new_n641), .C1(new_n620), .C2(new_n395), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n610), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n639), .A2(new_n643), .A3(new_n573), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  INV_X1    g460(.A(new_n285), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n274), .A2(new_n282), .A3(new_n283), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(KEYINPUT38), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n641), .B(KEYINPUT39), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n589), .A2(KEYINPUT40), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n325), .A2(new_n326), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n608), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n635), .A2(new_n187), .ZN(new_n656));
  NOR4_X1   g470(.A1(new_n650), .A2(new_n653), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(KEYINPUT40), .B1(new_n589), .B2(new_n652), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n463), .A2(new_n465), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n455), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n455), .B1(new_n479), .B2(new_n451), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n661), .A2(KEYINPUT97), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT97), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n448), .B1(new_n463), .B2(new_n465), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n665), .B1(new_n666), .B2(new_n662), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n664), .A2(new_n328), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT98), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n669), .A3(G472), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n638), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n669), .B1(new_n668), .B2(G472), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n659), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(new_n241), .ZN(G45));
  NAND3_X1  g489(.A1(new_n607), .A2(new_n608), .A3(new_n641), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n639), .A2(new_n573), .A3(new_n644), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  NAND3_X1  g493(.A1(new_n611), .A2(new_n486), .A3(new_n531), .ZN(new_n680));
  AOI21_X1  g494(.A(G902), .B1(new_n568), .B2(new_n569), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT99), .ZN(new_n682));
  OAI21_X1  g496(.A(G469), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n561), .A2(new_n567), .B1(new_n564), .B2(new_n548), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n684), .A2(KEYINPUT99), .A3(G902), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT100), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n681), .A2(new_n682), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT99), .B1(new_n684), .B2(G902), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT100), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n687), .A2(new_n688), .A3(new_n689), .A4(G469), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n686), .A2(new_n588), .A3(new_n572), .A4(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n680), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT41), .B(G113), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND3_X1  g508(.A1(new_n486), .A2(new_n622), .A3(new_n531), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n691), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n212), .ZN(G18));
  NOR2_X1   g511(.A1(new_n396), .A2(new_n294), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n486), .A2(new_n698), .A3(new_n644), .A4(new_n630), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n691), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n210), .ZN(G21));
  XOR2_X1   g515(.A(new_n483), .B(KEYINPUT101), .Z(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n466), .A2(new_n467), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n455), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n478), .A2(new_n481), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n703), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n528), .A2(new_n529), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n708), .A2(new_n709), .A3(new_n580), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n610), .A2(new_n655), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n711), .A3(new_n617), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n691), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT102), .B(G122), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G24));
  AND3_X1   g529(.A1(new_n686), .A2(new_n572), .A3(new_n690), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n448), .B1(new_n466), .B2(new_n467), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n702), .B1(new_n717), .B2(new_n706), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n482), .A2(new_n328), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n630), .B(new_n718), .C1(new_n719), .C2(new_n579), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n676), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n716), .A2(new_n588), .A3(new_n644), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G125), .ZN(G27));
  INV_X1    g537(.A(new_n709), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n486), .A2(new_n677), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n647), .A2(new_n648), .A3(new_n187), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n573), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT42), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n589), .A2(new_n726), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n676), .A2(KEYINPUT42), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n730), .A2(new_n486), .A3(new_n531), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n338), .ZN(G33));
  XNOR2_X1  g548(.A(new_n642), .B(KEYINPUT103), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n735), .A2(new_n730), .A3(new_n486), .A4(new_n531), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G134), .ZN(G36));
  NAND2_X1  g551(.A1(new_n618), .A2(new_n619), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n738), .A2(new_n739), .B1(new_n374), .B2(new_n376), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n607), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n742), .B1(new_n743), .B2(KEYINPUT43), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n744), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n582), .A3(new_n630), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n727), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n565), .A2(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n565), .A2(KEYINPUT45), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(G469), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT46), .B1(new_n755), .B2(new_n583), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n756), .B1(new_n571), .B2(new_n681), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n583), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n588), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n652), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n747), .A2(new_n748), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n749), .A2(KEYINPUT105), .A3(new_n727), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n752), .A2(new_n761), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  XOR2_X1   g579(.A(new_n760), .B(KEYINPUT47), .Z(new_n766));
  NOR4_X1   g580(.A1(new_n486), .A2(new_n531), .A3(new_n676), .A4(new_n726), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  INV_X1    g583(.A(new_n640), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n746), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT110), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n588), .A2(new_n686), .A3(new_n572), .A4(new_n690), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n772), .A2(new_n773), .A3(new_n727), .ZN(new_n774));
  OR3_X1    g588(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n479), .A2(new_n451), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT29), .B1(new_n776), .B2(new_n455), .ZN(new_n777));
  AOI21_X1  g591(.A(G902), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n579), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n780), .B1(new_n636), .B2(new_n637), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n709), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n774), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT48), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n576), .A2(new_n289), .ZN(new_n785));
  AND4_X1   g599(.A1(new_n673), .A2(new_n773), .A3(new_n727), .A4(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n608), .A3(new_n607), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n288), .A2(G952), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n772), .A2(new_n710), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n691), .A2(new_n610), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n784), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n720), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n607), .A2(new_n608), .ZN(new_n794));
  AOI22_X1  g608(.A1(new_n774), .A2(new_n793), .B1(new_n786), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT111), .ZN(new_n797));
  INV_X1    g611(.A(new_n650), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n798), .A2(new_n187), .A3(new_n691), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n789), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n797), .B1(new_n789), .B2(new_n799), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n795), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n716), .A2(new_n534), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n766), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n789), .A2(new_n727), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n802), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  XOR2_X1   g621(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n808));
  NAND2_X1  g622(.A1(new_n802), .A2(KEYINPUT112), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n804), .A2(new_n806), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(KEYINPUT51), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n802), .A2(KEYINPUT112), .ZN(new_n812));
  OAI221_X1 g626(.A(new_n792), .B1(new_n807), .B2(new_n808), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n699), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n710), .A2(new_n711), .A3(new_n617), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n773), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n781), .A2(new_n576), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n817), .B(new_n773), .C1(new_n611), .C2(new_n622), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT106), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n816), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n691), .B1(new_n699), .B2(new_n712), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n691), .B1(new_n680), .B2(new_n695), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT106), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n396), .B1(new_n740), .B2(new_n607), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n188), .B(new_n617), .C1(new_n284), .C2(new_n285), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(new_n531), .A3(new_n573), .A4(new_n581), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n574), .A3(new_n631), .ZN(new_n828));
  INV_X1    g642(.A(new_n721), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n620), .A2(new_n395), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n327), .A2(new_n377), .A3(new_n641), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n486), .A2(new_n630), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n728), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n828), .A2(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n729), .A2(new_n736), .A3(new_n732), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n820), .A2(new_n823), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT107), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n729), .A2(new_n736), .A3(new_n732), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n839), .A2(new_n834), .A3(new_n828), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT107), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n841), .A3(new_n823), .A4(new_n820), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n486), .A2(new_n573), .A3(new_n644), .A4(new_n630), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n790), .A2(new_n721), .B1(new_n843), .B2(new_n643), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n588), .A2(new_n587), .A3(new_n635), .A4(new_n641), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n846), .B(new_n711), .C1(new_n672), .C2(new_n671), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n844), .A2(new_n845), .A3(new_n678), .A4(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n722), .A2(new_n645), .A3(new_n678), .A4(new_n847), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT52), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n838), .A2(new_n842), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n821), .A2(new_n822), .A3(new_n853), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n722), .A2(new_n645), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT52), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n840), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n848), .A2(new_n850), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n854), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(KEYINPUT54), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n859), .B1(KEYINPUT107), .B2(new_n837), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n857), .A2(new_n853), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n842), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n864), .B1(new_n854), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT108), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n854), .A2(new_n867), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT54), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT108), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n871), .B(new_n872), .C1(KEYINPUT54), .C2(new_n862), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  OAI22_X1  g688(.A1(new_n813), .A2(new_n874), .B1(G952), .B2(G953), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n724), .A2(new_n742), .A3(new_n588), .A4(new_n188), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n650), .A3(new_n673), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n716), .B(KEYINPUT49), .Z(new_n878));
  OAI21_X1  g692(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(G75));
  AND2_X1   g693(.A1(new_n278), .A2(new_n281), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n279), .ZN(new_n881));
  XNOR2_X1  g695(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n881), .B(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n862), .A2(G902), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT114), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n860), .B1(new_n852), .B2(new_n853), .ZN(new_n887));
  OR3_X1    g701(.A1(new_n887), .A2(KEYINPUT114), .A3(new_n328), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n884), .B1(new_n889), .B2(new_n283), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n288), .A2(G952), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT56), .ZN(new_n892));
  INV_X1    g706(.A(G210), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n892), .B1(new_n885), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n891), .B1(new_n894), .B2(new_n883), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n890), .A2(new_n895), .ZN(G51));
  XNOR2_X1  g710(.A(new_n887), .B(new_n864), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n583), .B(KEYINPUT57), .Z(new_n898));
  AOI21_X1  g712(.A(new_n684), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n755), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n886), .A2(new_n900), .A3(new_n888), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n899), .B1(KEYINPUT115), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n901), .A2(KEYINPUT115), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n891), .B1(new_n902), .B2(new_n903), .ZN(G54));
  AND2_X1   g718(.A1(KEYINPUT58), .A2(G475), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n886), .A2(new_n888), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n390), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n891), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n886), .A2(new_n390), .A3(new_n888), .A4(new_n905), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT116), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT116), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n908), .A2(new_n913), .A3(new_n909), .A4(new_n910), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(G60));
  AND2_X1   g729(.A1(new_n596), .A2(new_n601), .ZN(new_n916));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT59), .Z(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n891), .B1(new_n897), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n918), .B1(new_n869), .B2(new_n873), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(new_n916), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT117), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT117), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n925), .B(new_n921), .C1(new_n922), .C2(new_n916), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(G63));
  INV_X1    g741(.A(new_n515), .ZN(new_n928));
  XNOR2_X1  g742(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n317), .A2(new_n328), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n928), .B1(new_n887), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT53), .B1(new_n865), .B2(new_n842), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n628), .B(new_n931), .C1(new_n934), .C2(new_n860), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n935), .A3(new_n909), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n936), .A2(KEYINPUT119), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT119), .B1(new_n936), .B2(new_n937), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n933), .A2(new_n935), .A3(KEYINPUT61), .A4(new_n909), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT120), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT121), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n862), .A2(new_n931), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n891), .B1(new_n944), .B2(new_n928), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n945), .A2(KEYINPUT120), .A3(KEYINPUT61), .A4(new_n935), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT120), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n941), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT121), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n949), .B(new_n950), .C1(new_n939), .C2(new_n938), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n943), .A2(new_n951), .ZN(G66));
  AOI21_X1  g766(.A(new_n288), .B1(new_n291), .B2(G224), .ZN(new_n953));
  INV_X1    g767(.A(new_n828), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n820), .A2(new_n823), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n953), .B1(new_n955), .B2(new_n288), .ZN(new_n956));
  INV_X1    g770(.A(G898), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n880), .B1(new_n957), .B2(G953), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n956), .B(new_n958), .ZN(G69));
  INV_X1    g773(.A(KEYINPUT123), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n844), .A2(new_n678), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n782), .A2(new_n711), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n839), .B1(new_n761), .B2(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n768), .A2(new_n764), .A3(new_n962), .A4(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n965), .A2(G953), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n432), .B1(KEYINPUT30), .B2(new_n474), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT122), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n382), .B1(new_n358), .B2(new_n383), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n968), .B(new_n969), .Z(new_n970));
  INV_X1    g784(.A(G900), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(new_n288), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n768), .A2(new_n764), .ZN(new_n973));
  OAI21_X1  g787(.A(KEYINPUT62), .B1(new_n674), .B2(new_n961), .ZN(new_n974));
  OR3_X1    g788(.A1(new_n674), .A2(KEYINPUT62), .A3(new_n961), .ZN(new_n975));
  INV_X1    g789(.A(new_n824), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n817), .A2(new_n651), .A3(new_n730), .A4(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n977), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n978), .A2(new_n288), .ZN(new_n979));
  OAI221_X1 g793(.A(new_n960), .B1(new_n966), .B2(new_n972), .C1(new_n979), .C2(new_n970), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n288), .B1(G227), .B2(G900), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G72));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n978), .B2(new_n955), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT124), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n663), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n986), .B2(new_n985), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n776), .A2(new_n448), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n990), .A2(new_n663), .A3(new_n984), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT126), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n870), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT127), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT125), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n995), .B(new_n984), .C1(new_n965), .C2(new_n955), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n996), .A2(new_n989), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n984), .B1(new_n965), .B2(new_n955), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(KEYINPUT125), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n891), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n988), .A2(new_n994), .A3(new_n1000), .ZN(G57));
endmodule


