//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  INV_X1    g0011(.A(new_n201), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n208), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n211), .B(new_n218), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n202), .A2(G68), .ZN(new_n242));
  INV_X1    g0042(.A(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n241), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT79), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G50), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n215), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n254), .B1(new_n250), .B2(G20), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n252), .B1(new_n255), .B2(G50), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n203), .A2(G20), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G58), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT8), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT8), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G58), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n263), .A2(new_n265), .A3(KEYINPUT65), .ZN(new_n266));
  AOI21_X1  g0066(.A(KEYINPUT65), .B1(new_n263), .B2(new_n265), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n216), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n261), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n254), .ZN(new_n272));
  OAI211_X1 g0072(.A(KEYINPUT9), .B(new_n256), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT9), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT65), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT65), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n264), .A2(G58), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n262), .A2(KEYINPUT8), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n276), .A2(new_n280), .A3(new_n270), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n259), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n272), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n256), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n274), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT64), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n215), .ZN(new_n289));
  NAND3_X1  g0089(.A1(KEYINPUT64), .A2(G33), .A3(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G41), .ZN(new_n292));
  INV_X1    g0092(.A(G45), .ZN(new_n293));
  AOI21_X1  g0093(.A(G1), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(G274), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n294), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n291), .A2(new_n296), .A3(G226), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT3), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT3), .ZN(new_n302));
  INV_X1    g0102(.A(G1698), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n300), .A2(new_n302), .A3(G222), .A4(new_n303), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n300), .A2(new_n302), .A3(G223), .A4(G1698), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n300), .A2(new_n302), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n304), .B(new_n305), .C1(new_n306), .C2(new_n220), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n289), .A2(new_n286), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G190), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n298), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(G200), .B1(new_n298), .B2(new_n310), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n273), .B(new_n285), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT10), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n298), .A2(new_n310), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n298), .A2(new_n310), .A3(new_n311), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT10), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(new_n285), .A4(new_n273), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n300), .A2(new_n302), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G107), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n300), .A2(new_n302), .A3(G238), .A4(G1698), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n300), .A2(new_n302), .A3(G232), .A4(new_n303), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT66), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT66), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n325), .A2(new_n330), .A3(new_n326), .A4(new_n327), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n309), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n291), .A2(new_n296), .A3(G244), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n295), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(G169), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n255), .A2(G77), .ZN(new_n337));
  INV_X1    g0137(.A(new_n251), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n220), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT15), .B(G87), .ZN(new_n341));
  OR3_X1    g0141(.A1(new_n341), .A2(KEYINPUT67), .A3(new_n269), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT67), .B1(new_n341), .B2(new_n269), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n263), .A2(new_n265), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n340), .B1(new_n346), .B2(new_n254), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT68), .B1(new_n336), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n254), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(new_n339), .A3(new_n337), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT68), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n331), .A2(new_n309), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n334), .B1(new_n352), .B2(new_n329), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n350), .B(new_n351), .C1(new_n353), .C2(G169), .ZN(new_n354));
  INV_X1    g0154(.A(G179), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n348), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n350), .B1(new_n353), .B2(G190), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n317), .B2(new_n353), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n316), .A2(G179), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n283), .A2(new_n284), .ZN(new_n361));
  AOI21_X1  g0161(.A(G169), .B1(new_n298), .B2(new_n310), .ZN(new_n362));
  NOR3_X1   g0162(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n323), .A2(new_n357), .A3(new_n359), .A4(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT69), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n363), .B1(new_n315), .B2(new_n322), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n368), .A2(KEYINPUT69), .A3(new_n357), .A4(new_n359), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT70), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n259), .A2(G50), .B1(G20), .B2(new_n243), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n220), .B2(new_n269), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n254), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT11), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n374), .A2(new_n375), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n371), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n378), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(KEYINPUT70), .A3(new_n376), .ZN(new_n381));
  OR3_X1    g0181(.A1(new_n251), .A2(KEYINPUT12), .A3(G68), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT12), .B1(new_n251), .B2(G68), .ZN(new_n383));
  AOI22_X1  g0183(.A1(G68), .A2(new_n255), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n379), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT14), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT13), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n300), .A2(new_n302), .A3(G232), .A4(G1698), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n300), .A2(new_n302), .A3(G226), .A4(new_n303), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G97), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n309), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n291), .A2(new_n296), .A3(G238), .ZN(new_n393));
  AND4_X1   g0193(.A1(new_n387), .A2(new_n392), .A3(new_n295), .A4(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n295), .A2(new_n393), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n387), .B1(new_n395), .B2(new_n392), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n386), .B(G169), .C1(new_n394), .C2(new_n396), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n391), .A2(new_n309), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n295), .A2(new_n393), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT13), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n395), .A2(new_n387), .A3(new_n392), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(G179), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n400), .A2(new_n401), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n386), .B1(new_n404), .B2(G169), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n385), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n385), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(G200), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n400), .A2(G190), .A3(new_n401), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT71), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT71), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n406), .A2(new_n413), .A3(new_n410), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n370), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n301), .A2(KEYINPUT72), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT72), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G33), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n419), .A3(KEYINPUT3), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT73), .B1(new_n301), .B2(KEYINPUT3), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT73), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n417), .A2(new_n419), .A3(new_n424), .A4(KEYINPUT3), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G226), .A2(G1698), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n303), .A2(G223), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n427), .B1(new_n428), .B2(KEYINPUT77), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G87), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n431), .B(KEYINPUT78), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT77), .ZN(new_n434));
  INV_X1    g0234(.A(new_n428), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n434), .B1(new_n426), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n309), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n291), .A2(new_n296), .A3(G232), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n437), .A2(G179), .A3(new_n295), .A4(new_n438), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT72), .B(G33), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n421), .B1(new_n440), .B2(KEYINPUT3), .ZN(new_n441));
  AND4_X1   g0241(.A1(new_n424), .A2(new_n417), .A3(new_n419), .A4(KEYINPUT3), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT77), .B1(new_n443), .B2(new_n428), .ZN(new_n444));
  INV_X1    g0244(.A(new_n432), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n426), .B2(new_n429), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n308), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n295), .A2(new_n438), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(G169), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n439), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n262), .A2(new_n243), .ZN(new_n452));
  OAI21_X1  g0252(.A(G20), .B1(new_n452), .B2(new_n201), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT74), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT74), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n455), .B(G20), .C1(new_n452), .C2(new_n201), .ZN(new_n456));
  INV_X1    g0256(.A(G159), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n454), .B(new_n456), .C1(new_n457), .C2(new_n260), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n302), .B1(new_n440), .B2(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n216), .A2(KEYINPUT7), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT7), .B1(new_n324), .B2(new_n216), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n458), .B1(G68), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n254), .B1(new_n466), .B2(KEYINPUT16), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n423), .A2(new_n216), .A3(new_n425), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT7), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT7), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n423), .A2(new_n470), .A3(new_n216), .A4(new_n425), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(G68), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n458), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(KEYINPUT16), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT75), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n243), .B1(new_n468), .B2(KEYINPUT7), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n458), .B1(new_n476), .B2(new_n471), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT75), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT16), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n467), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n268), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n251), .ZN(new_n482));
  INV_X1    g0282(.A(new_n255), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n268), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT76), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n451), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT18), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n463), .B1(new_n459), .B2(new_n461), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n473), .B1(new_n243), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT16), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n272), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AND4_X1   g0292(.A1(new_n478), .A2(new_n472), .A3(KEYINPUT16), .A4(new_n473), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n478), .B1(new_n477), .B2(KEYINPUT16), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n317), .B1(new_n447), .B2(new_n448), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n437), .A2(new_n295), .A3(new_n438), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(G190), .ZN(new_n498));
  INV_X1    g0298(.A(new_n486), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n495), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT17), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT18), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n451), .B(new_n503), .C1(new_n480), .C2(new_n486), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n495), .A2(new_n498), .A3(KEYINPUT17), .A4(new_n499), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n488), .A2(new_n502), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n249), .B1(new_n416), .B2(new_n506), .ZN(new_n507));
  AND4_X1   g0307(.A1(new_n488), .A2(new_n502), .A3(new_n504), .A4(new_n505), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n508), .A2(KEYINPUT79), .A3(new_n415), .A4(new_n370), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT24), .ZN(new_n511));
  INV_X1    g0311(.A(G87), .ZN(new_n512));
  NOR4_X1   g0312(.A1(new_n324), .A2(KEYINPUT22), .A3(G20), .A4(new_n512), .ZN(new_n513));
  AOI211_X1 g0313(.A(G20), .B(new_n512), .C1(new_n423), .C2(new_n425), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT22), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT85), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n216), .B(G87), .C1(new_n441), .C2(new_n442), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT85), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT22), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n513), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n222), .A2(G20), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n521), .A2(KEYINPUT23), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(KEYINPUT23), .ZN(new_n523));
  INV_X1    g0323(.A(G116), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n440), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n522), .B(new_n523), .C1(new_n526), .C2(G20), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n511), .B1(new_n520), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n513), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT22), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n518), .B1(new_n517), .B2(KEYINPUT22), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n527), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n532), .A2(KEYINPUT24), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n528), .A2(new_n254), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n338), .A2(new_n222), .ZN(new_n536));
  NOR2_X1   g0336(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n537));
  OR2_X1    g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n536), .B2(new_n537), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n250), .A2(G33), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n272), .A2(new_n251), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n538), .A2(new_n540), .B1(new_n543), .B2(G107), .ZN(new_n544));
  INV_X1    g0344(.A(G250), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n303), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(G257), .B2(new_n303), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n423), .B2(new_n425), .ZN(new_n548));
  INV_X1    g0348(.A(G294), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n440), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n309), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n291), .A2(G274), .ZN(new_n552));
  AND2_X1   g0352(.A1(KEYINPUT5), .A2(G41), .ZN(new_n553));
  NOR2_X1   g0353(.A1(KEYINPUT5), .A2(G41), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n250), .B(G45), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  OR2_X1    g0355(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n555), .A2(new_n291), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G264), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n551), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n317), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(G190), .B2(new_n559), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n535), .A2(new_n544), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n544), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n532), .A2(new_n533), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n272), .B1(new_n564), .B2(new_n511), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n563), .B1(new_n565), .B2(new_n534), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n559), .A2(G179), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n450), .B2(new_n559), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n562), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n557), .A2(G257), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n556), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(KEYINPUT4), .A2(G244), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n300), .A2(new_n302), .A3(new_n575), .A4(new_n303), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n300), .A2(new_n302), .A3(G250), .A4(G1698), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G283), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n221), .A2(G1698), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n423), .B2(new_n425), .ZN(new_n583));
  XOR2_X1   g0383(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n580), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT81), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n309), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n581), .B1(new_n441), .B2(new_n442), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n584), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT81), .B1(new_n590), .B2(new_n580), .ZN(new_n591));
  OAI211_X1 g0391(.A(G190), .B(new_n574), .C1(new_n588), .C2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(G97), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n338), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n542), .B2(new_n593), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n222), .A2(KEYINPUT6), .A3(G97), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n593), .A2(new_n222), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n597), .A2(new_n205), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n598), .B2(KEYINPUT6), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n599), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n489), .B2(new_n222), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n595), .B1(new_n601), .B2(new_n254), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n592), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n574), .B1(new_n588), .B2(new_n591), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n317), .B1(new_n604), .B2(KEYINPUT82), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT82), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n606), .B(new_n574), .C1(new_n588), .C2(new_n591), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n603), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n355), .B(new_n574), .C1(new_n588), .C2(new_n591), .ZN(new_n609));
  INV_X1    g0409(.A(new_n602), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n579), .B1(new_n589), .B2(new_n584), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n308), .B1(new_n611), .B2(KEYINPUT81), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n586), .A2(new_n587), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n573), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n609), .B(new_n610), .C1(new_n614), .C2(G169), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n221), .A2(G1698), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(G238), .B2(G1698), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n423), .B2(new_n425), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n309), .B1(new_n619), .B2(new_n525), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n545), .B1(new_n293), .B2(G1), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n250), .A2(G45), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n291), .B(new_n621), .C1(G274), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G169), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n620), .A2(G179), .A3(new_n623), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n341), .A2(new_n338), .ZN(new_n628));
  INV_X1    g0428(.A(new_n341), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n543), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(G20), .B1(new_n423), .B2(new_n425), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n205), .A2(new_n512), .B1(new_n390), .B2(new_n216), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT19), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n270), .A2(new_n633), .A3(G97), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n631), .A2(G68), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n628), .B(new_n630), .C1(new_n636), .C2(new_n272), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT83), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n628), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n216), .B(G68), .C1(new_n441), .C2(new_n442), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n634), .A2(new_n635), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n640), .B1(new_n643), .B2(new_n254), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n644), .A2(KEYINPUT83), .A3(new_n630), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n627), .A2(new_n639), .A3(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n620), .A2(G190), .A3(new_n623), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n317), .B1(new_n620), .B2(new_n623), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n542), .A2(new_n512), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n628), .B(new_n651), .C1(new_n636), .C2(new_n272), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n646), .A2(new_n654), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n608), .A2(new_n616), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n223), .A2(G1698), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(G257), .B2(G1698), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n423), .B2(new_n425), .ZN(new_n659));
  INV_X1    g0459(.A(G303), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n306), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n309), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n555), .A2(new_n291), .A3(G270), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT84), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n555), .A2(new_n291), .A3(KEYINPUT84), .A4(G270), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n662), .A2(new_n556), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n578), .B(new_n216), .C1(G33), .C2(new_n593), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n670), .B(new_n254), .C1(new_n216), .C2(G116), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT20), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n251), .A2(G116), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n543), .B2(G116), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n669), .A2(G179), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n450), .B1(new_n673), .B2(new_n675), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT21), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n678), .A2(new_n668), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n679), .B1(new_n678), .B2(new_n668), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n677), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n669), .A2(G190), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n676), .B1(new_n668), .B2(G200), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  AND4_X1   g0486(.A1(new_n510), .A2(new_n571), .A3(new_n656), .A4(new_n686), .ZN(G372));
  AOI21_X1  g0487(.A(new_n610), .B1(new_n614), .B2(G190), .ZN(new_n688));
  OAI21_X1  g0488(.A(G200), .B1(new_n614), .B2(new_n606), .ZN(new_n689));
  INV_X1    g0489(.A(new_n607), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n625), .A2(new_n626), .B1(new_n644), .B2(new_n630), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT87), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n652), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n644), .A2(KEYINPUT87), .A3(new_n651), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n692), .B1(new_n696), .B2(new_n649), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n562), .A2(new_n691), .A3(new_n615), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n535), .A2(new_n544), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n682), .B1(new_n699), .B2(new_n568), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n692), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT26), .B1(new_n616), .B2(new_n697), .ZN(new_n703));
  XNOR2_X1  g0503(.A(KEYINPUT88), .B(KEYINPUT26), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n655), .A2(new_n615), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n702), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n510), .B1(new_n701), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n406), .A2(new_n357), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n505), .A2(new_n502), .A3(new_n410), .A4(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n488), .A2(new_n504), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n363), .B1(new_n711), .B2(new_n323), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n707), .A2(new_n712), .ZN(G369));
  INV_X1    g0513(.A(G13), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n714), .A2(G1), .A3(G20), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(KEYINPUT89), .A3(KEYINPUT27), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(KEYINPUT89), .B1(new_n716), .B2(KEYINPUT27), .ZN(new_n719));
  OAI221_X1 g0519(.A(G213), .B1(KEYINPUT27), .B2(new_n716), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(G343), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n571), .B1(new_n566), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n699), .A2(new_n568), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n724), .B1(new_n725), .B2(new_n723), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n722), .A2(new_n676), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n686), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n682), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n728), .B1(new_n729), .B2(new_n727), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G330), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n729), .A2(new_n722), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n571), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n733), .B(new_n735), .C1(new_n725), .C2(new_n722), .ZN(G399));
  INV_X1    g0536(.A(new_n209), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G41), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n739), .A2(G1), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(new_n213), .B2(new_n739), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  INV_X1    g0543(.A(G330), .ZN(new_n744));
  XOR2_X1   g0544(.A(KEYINPUT90), .B(KEYINPUT30), .Z(new_n745));
  NAND2_X1  g0545(.A1(new_n551), .A2(new_n558), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n626), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n669), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n745), .B1(new_n748), .B2(new_n604), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n614), .A2(KEYINPUT30), .A3(new_n669), .A4(new_n747), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n559), .A2(new_n355), .A3(new_n624), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n751), .A2(new_n604), .A3(new_n668), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n722), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(KEYINPUT31), .B1(new_n753), .B2(new_n722), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n682), .A2(new_n685), .A3(new_n722), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n656), .A2(new_n725), .A3(new_n562), .A4(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n744), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n723), .B1(new_n701), .B2(new_n706), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT29), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n702), .B1(new_n698), .B2(new_n700), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT91), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n765), .B(new_n704), .C1(new_n655), .C2(new_n615), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n616), .A2(KEYINPUT26), .A3(new_n697), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n602), .B1(new_n604), .B2(new_n450), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n769), .A2(new_n646), .A3(new_n654), .A4(new_n609), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n765), .B1(new_n770), .B2(new_n704), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g0572(.A(KEYINPUT29), .B(new_n723), .C1(new_n764), .C2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n760), .B1(new_n763), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n743), .B1(new_n774), .B2(G1), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT92), .Z(G364));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT93), .Z(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n216), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT94), .Z(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n215), .B1(G20), .B2(new_n450), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n426), .A2(new_n737), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n214), .A2(new_n293), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n786), .B(new_n787), .C1(new_n247), .C2(new_n293), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n737), .A2(new_n324), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n789), .A2(G355), .B1(new_n524), .B2(new_n737), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n785), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n714), .A2(G20), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n250), .B1(new_n792), .B2(G45), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n738), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n783), .ZN(new_n797));
  NOR4_X1   g0597(.A1(new_n216), .A2(new_n355), .A3(new_n311), .A4(G200), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G322), .ZN(new_n800));
  INV_X1    g0600(.A(G311), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n216), .A2(G190), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n802), .A2(G179), .A3(new_n317), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n799), .A2(new_n800), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G179), .A2(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n306), .B(new_n804), .C1(G329), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n216), .A2(new_n355), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n809), .A2(G190), .A3(G200), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT96), .Z(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(KEYINPUT97), .B(G326), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n216), .A2(G179), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n815), .A2(G190), .A3(G200), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n216), .B1(new_n805), .B2(G190), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n817), .A2(G303), .B1(new_n819), .B2(G294), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n809), .A2(G200), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(G190), .ZN(new_n822));
  XNOR2_X1  g0622(.A(KEYINPUT33), .B(G317), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n815), .A2(new_n311), .A3(G200), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n822), .A2(new_n823), .B1(new_n825), .B2(G283), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n808), .A2(new_n814), .A3(new_n820), .A4(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n822), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n828), .A2(new_n243), .B1(new_n818), .B2(new_n593), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n807), .A2(G159), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n830), .A2(KEYINPUT32), .B1(new_n512), .B2(new_n816), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n803), .A2(KEYINPUT95), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n803), .A2(KEYINPUT95), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(G77), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n306), .B1(new_n799), .B2(new_n262), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(G107), .B2(new_n825), .ZN(new_n839));
  INV_X1    g0639(.A(new_n810), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n830), .A2(KEYINPUT32), .B1(new_n840), .B2(G50), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n832), .A2(new_n837), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n797), .B1(new_n827), .B2(new_n842), .ZN(new_n843));
  NOR3_X1   g0643(.A1(new_n791), .A2(new_n796), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n730), .B2(new_n781), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n731), .A2(new_n796), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n730), .A2(G330), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(G396));
  NOR2_X1   g0648(.A1(new_n783), .A2(new_n777), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n796), .B1(new_n220), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(G283), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n828), .A2(new_n851), .B1(new_n810), .B2(new_n660), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G116), .B2(new_n836), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT98), .Z(new_n854));
  OAI221_X1 g0654(.A(new_n324), .B1(new_n806), .B2(new_n801), .C1(new_n222), .C2(new_n816), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n798), .A2(G294), .B1(new_n819), .B2(G97), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT99), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n855), .B(new_n857), .C1(G87), .C2(new_n825), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n840), .A2(G137), .B1(new_n798), .B2(G143), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n859), .B1(new_n828), .B2(new_n258), .C1(new_n835), .C2(new_n457), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT34), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n825), .A2(G68), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n202), .B2(new_n816), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n863), .A2(KEYINPUT100), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(KEYINPUT100), .ZN(new_n865));
  INV_X1    g0665(.A(G132), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n866), .A2(new_n806), .B1(new_n818), .B2(new_n262), .ZN(new_n867));
  NOR4_X1   g0667(.A1(new_n864), .A2(new_n865), .A3(new_n443), .A4(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n854), .A2(new_n858), .B1(new_n861), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n723), .A2(new_n347), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n357), .B2(new_n359), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n357), .A2(new_n870), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n850), .B1(new_n797), .B2(new_n869), .C1(new_n873), .C2(new_n778), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n729), .B1(new_n566), .B2(new_n569), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT87), .B1(new_n644), .B2(new_n651), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n272), .B1(new_n641), .B2(new_n642), .ZN(new_n878));
  NOR4_X1   g0678(.A1(new_n878), .A2(new_n693), .A3(new_n640), .A4(new_n650), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n649), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n702), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n608), .A2(new_n616), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n876), .A2(new_n882), .A3(new_n562), .ZN(new_n883));
  OR3_X1    g0683(.A1(new_n655), .A2(new_n615), .A3(new_n704), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT26), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n881), .B2(new_n615), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n692), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n722), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n873), .ZN(new_n889));
  INV_X1    g0689(.A(new_n873), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n761), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n760), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(new_n795), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n889), .A2(new_n891), .A3(new_n760), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n875), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(G384));
  OR2_X1    g0696(.A1(new_n599), .A2(KEYINPUT35), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n599), .A2(KEYINPUT35), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n897), .A2(G116), .A3(new_n217), .A4(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n899), .B(KEYINPUT36), .Z(new_n900));
  OR3_X1    g0700(.A1(new_n213), .A2(new_n220), .A3(new_n452), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n250), .B(G13), .C1(new_n901), .C2(new_n242), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n720), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n710), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n254), .B1(new_n477), .B2(KEYINPUT16), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n479), .B2(new_n475), .ZN(new_n907));
  INV_X1    g0707(.A(new_n485), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n451), .B1(new_n907), .B2(new_n908), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(new_n910), .A3(new_n500), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT37), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n904), .B1(new_n480), .B2(new_n486), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT37), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n487), .A2(new_n913), .A3(new_n500), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n909), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n506), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT38), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n915), .A2(new_n912), .B1(new_n506), .B2(new_n917), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT38), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n357), .A2(new_n722), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT101), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n889), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n385), .A2(new_n722), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n411), .B(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n487), .A2(new_n913), .A3(new_n500), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT37), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n915), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT102), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT102), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n934), .A2(new_n937), .A3(new_n915), .ZN(new_n938));
  INV_X1    g0738(.A(new_n913), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n506), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n936), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n920), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT39), .B1(new_n922), .B2(KEYINPUT38), .ZN(new_n943));
  AOI22_X1  g0743(.A1(KEYINPUT39), .A2(new_n924), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n406), .A2(new_n722), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n905), .B1(new_n925), .B2(new_n932), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n510), .A2(new_n763), .A3(new_n773), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n712), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n946), .B(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n942), .A2(new_n923), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n753), .A2(new_n722), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT31), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n655), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n758), .A2(new_n691), .A3(new_n615), .A4(new_n954), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n953), .B(new_n754), .C1(new_n955), .C2(new_n570), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n956), .A2(new_n873), .A3(new_n931), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n957), .A2(KEYINPUT40), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n919), .A2(new_n920), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT38), .B1(new_n916), .B2(new_n918), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT40), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n950), .A2(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n963), .A2(new_n510), .A3(new_n956), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n950), .A2(new_n958), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n961), .A2(new_n962), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n510), .A2(new_n956), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n964), .A2(new_n969), .A3(G330), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n949), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n250), .B2(new_n792), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n949), .A2(new_n970), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n903), .B1(new_n972), .B2(new_n973), .ZN(G367));
  NOR2_X1   g0774(.A1(new_n608), .A2(new_n616), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n610), .A2(new_n722), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n975), .A2(new_n976), .B1(new_n616), .B2(new_n722), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n735), .A2(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT42), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(KEYINPUT42), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n615), .B1(new_n725), .B2(new_n608), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n979), .A2(new_n980), .B1(new_n723), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n696), .A2(new_n723), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n692), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n881), .B2(new_n983), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT43), .ZN(new_n986));
  OR3_X1    g0786(.A1(new_n982), .A2(KEYINPUT103), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(KEYINPUT103), .B1(new_n982), .B2(new_n986), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n982), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n987), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n733), .A2(new_n977), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n738), .B(KEYINPUT41), .Z(new_n994));
  OAI21_X1  g0794(.A(new_n735), .B1(new_n725), .B2(new_n722), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n995), .A2(new_n977), .ZN(new_n996));
  XOR2_X1   g0796(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n996), .B(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n995), .A2(new_n977), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT44), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n733), .A2(KEYINPUT105), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1003), .B(new_n1004), .Z(new_n1005));
  OAI21_X1  g0805(.A(new_n735), .B1(new_n726), .B2(new_n734), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(new_n732), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n774), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n994), .B1(new_n1010), .B2(new_n774), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n993), .B1(new_n1011), .B2(new_n794), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n784), .B1(new_n209), .B2(new_n341), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n786), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1014), .A2(new_n237), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n795), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n817), .A2(G58), .B1(new_n807), .B2(G137), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n812), .A2(G143), .B1(KEYINPUT107), .B2(new_n1017), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n824), .A2(new_n220), .B1(new_n818), .B2(new_n243), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n306), .B1(new_n799), .B2(new_n258), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(G159), .C2(new_n822), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n836), .A2(G50), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1017), .A2(KEYINPUT107), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1018), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n824), .A2(new_n593), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G317), .A2(new_n807), .B1(new_n798), .B2(G303), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n222), .B2(new_n818), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1025), .B(new_n1027), .C1(G294), .C2(new_n822), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n426), .B1(new_n836), .B2(G283), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(new_n801), .C2(new_n811), .ZN(new_n1030));
  AOI21_X1  g0830(.A(KEYINPUT106), .B1(new_n817), .B2(G116), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT46), .Z(new_n1032));
  OAI21_X1  g0832(.A(new_n1024), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT47), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1016), .B1(new_n1034), .B2(new_n783), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n985), .B2(new_n781), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1012), .A2(new_n1036), .ZN(G387));
  OR2_X1    g0837(.A1(new_n726), .A2(new_n781), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n789), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1039), .A2(new_n740), .B1(G107), .B2(new_n209), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n234), .A2(new_n293), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n740), .B(new_n293), .C1(new_n243), .C2(new_n220), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT50), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n275), .B2(G50), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n344), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1042), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1046), .A2(new_n1014), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1040), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n795), .B1(new_n785), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n810), .A2(new_n457), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT108), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n816), .A2(new_n220), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n818), .A2(new_n341), .ZN(new_n1053));
  NOR4_X1   g0853(.A1(new_n1051), .A2(new_n1025), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n799), .A2(new_n202), .B1(new_n806), .B2(new_n258), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n803), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n443), .B(new_n1055), .C1(G68), .C2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1054), .B(new_n1057), .C1(new_n481), .C2(new_n828), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n817), .A2(G294), .B1(new_n819), .B2(G283), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n822), .A2(G311), .B1(G317), .B2(new_n798), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n835), .B2(new_n660), .C1(new_n811), .C2(new_n800), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT109), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT49), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1068), .A2(KEYINPUT110), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n825), .A2(G116), .B1(new_n807), .B2(new_n813), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT110), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n443), .B(new_n1070), .C1(new_n1067), .C2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1058), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1049), .B1(new_n1073), .B2(new_n783), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1007), .A2(new_n794), .B1(new_n1038), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1008), .A2(new_n738), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1007), .A2(new_n774), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(G393));
  XNOR2_X1  g0878(.A(new_n1003), .B(new_n733), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1010), .B(new_n738), .C1(new_n1009), .C2(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n836), .A2(new_n344), .B1(G50), .B2(new_n822), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1081), .A2(KEYINPUT113), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n819), .A2(G77), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(KEYINPUT113), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT114), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n840), .A2(G150), .B1(new_n798), .B2(G159), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT51), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n807), .A2(G143), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n243), .B2(new_n816), .C1(new_n512), .C2(new_n824), .ZN(new_n1090));
  NOR4_X1   g0890(.A1(new_n1086), .A2(new_n443), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n840), .A2(G317), .B1(new_n798), .B2(G311), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT52), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n324), .B1(new_n806), .B2(new_n800), .C1(new_n549), .C2(new_n803), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n828), .A2(new_n660), .B1(new_n222), .B2(new_n824), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n816), .A2(new_n851), .B1(new_n818), .B2(new_n524), .ZN(new_n1096));
  NOR4_X1   g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n783), .B1(new_n1091), .B2(new_n1097), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n784), .B1(new_n593), .B2(new_n209), .C1(new_n241), .C2(new_n1014), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n795), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT112), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT115), .Z(new_n1103));
  NAND2_X1  g0903(.A1(new_n977), .A2(new_n782), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1104), .A2(KEYINPUT111), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(KEYINPUT111), .ZN(new_n1106));
  NOR3_X1   g0906(.A1(new_n1103), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n1079), .B2(new_n794), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1080), .A2(new_n1108), .ZN(G390));
  INV_X1    g0909(.A(new_n927), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n888), .B2(new_n873), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n945), .B1(new_n1111), .B2(new_n930), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n942), .A2(new_n943), .ZN(new_n1113));
  OAI21_X1  g0913(.A(KEYINPUT39), .B1(new_n959), .B2(new_n960), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n956), .A2(G330), .A3(new_n873), .A4(new_n931), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n723), .B(new_n873), .C1(new_n764), .C2(new_n772), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n926), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n931), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n950), .A2(new_n1122), .A3(new_n945), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1115), .A2(new_n1119), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n945), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n942), .B2(new_n923), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n944), .A2(new_n1112), .B1(new_n1126), .B2(new_n1122), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1116), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1124), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n510), .A2(new_n760), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n947), .A2(new_n712), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(KEYINPUT117), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT117), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n947), .A2(new_n1130), .A3(new_n1133), .A4(new_n712), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1116), .A2(KEYINPUT118), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n956), .A2(G330), .A3(new_n873), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n930), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(KEYINPUT118), .A3(new_n930), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n931), .B1(new_n760), .B2(new_n873), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1142), .A2(new_n1121), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1141), .A2(new_n928), .B1(new_n1118), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1135), .A2(new_n1144), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1129), .A2(new_n1145), .A3(KEYINPUT119), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT119), .B1(new_n1129), .B2(new_n1145), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n738), .B1(new_n1129), .B2(new_n1145), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n849), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n862), .B1(new_n549), .B2(new_n806), .C1(new_n524), .C2(new_n799), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1083), .B1(new_n851), .B2(new_n810), .C1(new_n828), .C2(new_n222), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(G97), .C2(new_n836), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n324), .B1(new_n816), .B2(new_n512), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT121), .Z(new_n1154));
  NAND2_X1  g0954(.A1(new_n822), .A2(G137), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT54), .B(G143), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1155), .B1(new_n835), .B2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT120), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n817), .A2(G150), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT53), .ZN(new_n1160));
  INV_X1    g0960(.A(G125), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n306), .B1(new_n806), .B2(new_n1161), .C1(new_n799), .C2(new_n866), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n825), .A2(G50), .B1(new_n819), .B2(G159), .ZN(new_n1163));
  INV_X1    g0963(.A(G128), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n810), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n1160), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1152), .A2(new_n1154), .B1(new_n1158), .B2(new_n1166), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n795), .B1(new_n268), .B2(new_n1149), .C1(new_n1167), .C2(new_n797), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n944), .B2(new_n779), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n1129), .B2(new_n794), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1148), .A2(new_n1170), .ZN(G378));
  NOR2_X1   g0971(.A1(new_n361), .A2(new_n720), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n368), .B(new_n1172), .Z(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1173), .B(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n963), .B2(G330), .ZN(new_n1177));
  AND4_X1   g0977(.A1(G330), .A2(new_n965), .A3(new_n966), .A4(new_n1176), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n946), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1175), .B1(new_n967), .B2(new_n744), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n905), .B1(new_n932), .B2(new_n925), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n944), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1181), .B1(new_n1182), .B2(new_n1125), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n963), .A2(G330), .A3(new_n1176), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT123), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1179), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1183), .B1(new_n1184), .B2(new_n1180), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT123), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1187), .A2(new_n1189), .A3(new_n794), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n795), .B1(G50), .B2(new_n1149), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT122), .Z(new_n1192));
  NOR2_X1   g0992(.A1(new_n824), .A2(new_n262), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G97), .B2(new_n822), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n524), .B2(new_n810), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n426), .A2(G41), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1056), .A2(new_n629), .B1(new_n798), .B2(G107), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n851), .B2(new_n806), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n816), .A2(new_n220), .B1(new_n818), .B2(new_n243), .ZN(new_n1200));
  NOR4_X1   g1000(.A1(new_n1195), .A2(new_n1197), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  AOI211_X1 g1001(.A(G50), .B(new_n1196), .C1(new_n301), .C2(new_n292), .ZN(new_n1202));
  OAI21_X1  g1002(.A(KEYINPUT58), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n828), .A2(new_n866), .B1(new_n810), .B2(new_n1161), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1056), .A2(G137), .B1(new_n798), .B2(G128), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n816), .B2(new_n1156), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(G150), .C2(new_n819), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n825), .A2(G159), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G33), .B(G41), .C1(new_n807), .C2(G124), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1203), .B1(KEYINPUT58), .B2(new_n1201), .C1(new_n1212), .C2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1192), .B1(new_n1214), .B2(new_n783), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1176), .B2(new_n778), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1190), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT119), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1115), .A2(new_n1119), .A3(new_n1123), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1128), .B1(new_n1115), .B2(new_n1123), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1118), .A2(new_n1143), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1111), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1132), .B(new_n1134), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1218), .B1(new_n1221), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1129), .A2(new_n1145), .A3(KEYINPUT119), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1135), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1185), .ZN(new_n1228));
  OAI21_X1  g1028(.A(KEYINPUT57), .B1(new_n1228), .B2(new_n1188), .ZN(new_n1229));
  OAI211_X1 g1029(.A(KEYINPUT124), .B(new_n738), .C1(new_n1227), .C2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT57), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1231), .B1(new_n1227), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1230), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1135), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1231), .B1(new_n1179), .B2(new_n1185), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT124), .B1(new_n1238), .B2(new_n738), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1217), .B1(new_n1234), .B2(new_n1239), .ZN(G375));
  NAND2_X1  g1040(.A1(new_n1135), .A2(new_n1144), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1242), .A2(new_n1145), .A3(new_n994), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1056), .A2(G150), .B1(new_n798), .B2(G137), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1164), .B2(new_n806), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1193), .B(new_n1245), .C1(G132), .C2(new_n840), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n828), .A2(new_n1156), .B1(new_n202), .B2(new_n818), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G159), .B2(new_n817), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1246), .A2(new_n426), .A3(new_n1248), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n828), .A2(new_n524), .B1(new_n816), .B2(new_n593), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G294), .B2(new_n840), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n836), .A2(G107), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n324), .B1(new_n806), .B2(new_n660), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G283), .B2(new_n798), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1053), .B1(G77), .B2(new_n825), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1251), .A2(new_n1252), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n797), .B1(new_n1249), .B2(new_n1256), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n796), .B(new_n1257), .C1(new_n243), .C2(new_n849), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n777), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1258), .B1(new_n931), .B2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1144), .B2(new_n793), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1243), .A2(new_n1261), .ZN(G381));
  OR4_X1    g1062(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1263), .A2(G387), .A3(G381), .ZN(new_n1264));
  INV_X1    g1064(.A(G378), .ZN(new_n1265));
  INV_X1    g1065(.A(G375), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(G407));
  NAND2_X1  g1067(.A1(new_n721), .A2(G213), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1268), .B(KEYINPUT125), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1265), .A3(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(G407), .A2(G213), .A3(new_n1270), .ZN(G409));
  OAI211_X1 g1071(.A(G378), .B(new_n1217), .C1(new_n1234), .C2(new_n1239), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1227), .A2(new_n1232), .A3(new_n994), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n794), .B1(new_n1228), .B2(new_n1188), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1216), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1265), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1272), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1135), .A2(KEYINPUT60), .A3(new_n1144), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1278), .A2(new_n738), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT60), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1241), .B1(new_n1145), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1261), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1282), .A2(G384), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(G384), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1277), .A2(new_n1268), .A3(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n721), .A2(G213), .A3(G2897), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1285), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT127), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1269), .A2(G2897), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1290), .A2(new_n1291), .A3(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1291), .B1(new_n1290), .B2(new_n1293), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1277), .A2(new_n1268), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1269), .B1(new_n1272), .B2(new_n1276), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(KEYINPUT63), .A3(new_n1285), .ZN(new_n1300));
  XOR2_X1   g1100(.A(G393), .B(G396), .Z(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1012), .A2(new_n1036), .A3(G390), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(G390), .B1(new_n1012), .B2(new_n1036), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1302), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1305), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1307), .A2(new_n1301), .A3(new_n1303), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT61), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1306), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1288), .A2(new_n1298), .A3(new_n1300), .A4(new_n1310), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1309), .B1(new_n1299), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT62), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1286), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1299), .A2(KEYINPUT62), .A3(new_n1285), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1313), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1311), .B1(new_n1317), .B2(new_n1319), .ZN(G405));
  NAND2_X1  g1120(.A1(G375), .A2(new_n1265), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1272), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1285), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1322), .A2(new_n1285), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1318), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1325), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1327), .A2(new_n1319), .A3(new_n1323), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1326), .A2(new_n1328), .ZN(G402));
endmodule


