//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n440, new_n446, new_n448, new_n450, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n579, new_n580,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(new_n440));
  INV_X1    g015(.A(new_n440), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  INV_X1    g024(.A(G567), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT67), .Z(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g028(.A1(G218), .A2(G219), .A3(G221), .A4(G220), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NAND4_X1  g030(.A1(new_n440), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G325));
  XOR2_X1   g034(.A(new_n458), .B(KEYINPUT69), .Z(G261));
  NOR2_X1   g035(.A1(new_n457), .A2(new_n450), .ZN(new_n461));
  INV_X1    g036(.A(new_n455), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(G2106), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n468), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT70), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n468), .A2(G137), .A3(new_n474), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n470), .A2(G101), .A3(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n475), .A2(new_n478), .ZN(G160));
  INV_X1    g054(.A(new_n474), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n468), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  INV_X1    g058(.A(new_n468), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n474), .C2(G112), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND3_X1  g064(.A1(new_n468), .A2(G138), .A3(new_n474), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n468), .A2(KEYINPUT4), .A3(G138), .A4(new_n474), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n468), .A2(G126), .A3(G2105), .ZN(new_n495));
  OR2_X1    g070(.A1(KEYINPUT71), .A2(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT71), .A2(G114), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n496), .A2(G2105), .A3(new_n497), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n498), .A2(G2104), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT72), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n495), .A2(new_n500), .A3(KEYINPUT72), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n494), .B1(new_n502), .B2(new_n503), .ZN(G164));
  AND2_X1   g079(.A1(KEYINPUT73), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT73), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT75), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G62), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT78), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n508), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n519), .B(KEYINPUT6), .C1(new_n505), .C2(new_n506), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT73), .A2(G651), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT74), .B1(new_n523), .B2(KEYINPUT6), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n520), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(new_n513), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT76), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n528), .A2(new_n531), .A3(new_n513), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n530), .A2(G88), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT77), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n528), .A2(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G50), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n534), .B1(new_n533), .B2(new_n536), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n518), .B1(new_n537), .B2(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  AND3_X1   g115(.A1(new_n528), .A2(new_n531), .A3(new_n513), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n531), .B1(new_n528), .B2(new_n513), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G89), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n535), .A2(G51), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT7), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n544), .A2(new_n545), .A3(new_n547), .A4(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  AOI22_X1  g125(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n508), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n528), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G52), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(new_n543), .B2(G90), .ZN(G171));
  AOI22_X1  g131(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n508), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n530), .A2(G81), .A3(new_n532), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n535), .A2(G43), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n560), .A2(KEYINPUT79), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(KEYINPUT79), .B1(new_n560), .B2(new_n561), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT80), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n566));
  INV_X1    g141(.A(G81), .ZN(new_n567));
  NOR3_X1   g142(.A1(new_n541), .A2(new_n542), .A3(new_n567), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n535), .A2(G43), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n560), .A2(KEYINPUT79), .A3(new_n561), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n572), .A2(new_n573), .A3(new_n559), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n565), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G860), .ZN(G153));
  AND3_X1   g151(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G36), .ZN(G176));
  NAND2_X1  g153(.A1(G1), .A2(G3), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT8), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(G188));
  NAND3_X1  g156(.A1(new_n530), .A2(G91), .A3(new_n532), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n583), .A2(new_n523), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT9), .ZN(new_n585));
  INV_X1    g160(.A(G53), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n553), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n535), .A2(KEYINPUT9), .A3(G53), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n582), .A2(new_n584), .A3(new_n587), .A4(new_n588), .ZN(G299));
  INV_X1    g164(.A(G171), .ZN(G301));
  OAI21_X1  g165(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n535), .A2(G49), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n530), .A2(new_n532), .ZN(new_n593));
  INV_X1    g168(.A(G87), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n591), .B(new_n592), .C1(new_n593), .C2(new_n594), .ZN(G288));
  AND2_X1   g170(.A1(new_n513), .A2(G61), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT81), .Z(new_n598));
  OAI21_X1  g173(.A(new_n507), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT82), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT82), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n601), .B(new_n507), .C1(new_n596), .C2(new_n598), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n530), .A2(G86), .A3(new_n532), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n535), .A2(G48), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(G305));
  NAND2_X1  g181(.A1(new_n543), .A2(G85), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n513), .A2(G60), .ZN(new_n608));
  INV_X1    g183(.A(G72), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n510), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n535), .A2(G47), .B1(new_n507), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n607), .A2(new_n611), .ZN(G290));
  NAND2_X1  g187(.A1(G301), .A2(G868), .ZN(new_n613));
  XOR2_X1   g188(.A(KEYINPUT83), .B(KEYINPUT10), .Z(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n593), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n543), .A2(G92), .A3(new_n614), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT84), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n620), .A2(G651), .B1(G54), .B2(new_n535), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n617), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n613), .B1(new_n623), .B2(G868), .ZN(G321));
  XNOR2_X1  g199(.A(G321), .B(KEYINPUT85), .ZN(G284));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(G299), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G168), .B2(new_n626), .ZN(G297));
  OAI21_X1  g203(.A(new_n627), .B1(G168), .B2(new_n626), .ZN(G280));
  INV_X1    g204(.A(G860), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n622), .B1(G559), .B2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT86), .Z(G148));
  NOR2_X1   g207(.A1(new_n622), .A2(G559), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n575), .B2(G868), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g212(.A1(new_n470), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  INV_X1    g214(.A(G2100), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT87), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  AOI22_X1  g218(.A1(G123), .A2(new_n482), .B1(new_n485), .B2(G135), .ZN(new_n644));
  INV_X1    g219(.A(G2096), .ZN(new_n645));
  OR3_X1    g220(.A1(new_n474), .A2(KEYINPUT88), .A3(G111), .ZN(new_n646));
  OAI21_X1  g221(.A(KEYINPUT88), .B1(new_n474), .B2(G111), .ZN(new_n647));
  OR2_X1    g222(.A1(G99), .A2(G2105), .ZN(new_n648));
  NAND4_X1  g223(.A1(new_n646), .A2(new_n647), .A3(G2104), .A4(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n644), .A2(new_n645), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n644), .A2(new_n649), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G2096), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n643), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT89), .Z(G156));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2435), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2438), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT14), .ZN(new_n659));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n659), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1341), .B(G1348), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n664), .B(new_n665), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(G14), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2067), .B(G2678), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT90), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2072), .B(G2078), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(new_n671), .B2(new_n672), .ZN(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n672), .B(KEYINPUT17), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n674), .B(new_n676), .C1(new_n669), .C2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT91), .Z(new_n680));
  NAND3_X1  g255(.A1(new_n670), .A2(new_n675), .A3(new_n672), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT18), .Z(new_n682));
  NAND3_X1  g257(.A1(new_n678), .A2(new_n675), .A3(new_n669), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(new_n645), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(new_n640), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G227));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n688), .A2(new_n689), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n691), .A2(new_n693), .A3(new_n695), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n698), .B(new_n699), .C1(new_n697), .C2(new_n696), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT21), .B(G1986), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G1991), .B(G1996), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT92), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT22), .B(G1981), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n705), .B(new_n706), .Z(G229));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G33), .ZN(new_n709));
  NAND2_X1  g284(.A1(G115), .A2(G2104), .ZN(new_n710));
  INV_X1    g285(.A(G127), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n484), .B2(new_n711), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n712), .A2(new_n480), .B1(new_n485), .B2(G139), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT25), .Z(new_n715));
  AND2_X1   g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n709), .B1(new_n716), .B2(new_n708), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G2072), .ZN(new_n718));
  NAND2_X1  g293(.A1(G299), .A2(G16), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n720), .A2(KEYINPUT23), .A3(G20), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT23), .ZN(new_n722));
  INV_X1    g297(.A(G20), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(G16), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n719), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT100), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1956), .ZN(new_n727));
  OR2_X1    g302(.A1(KEYINPUT24), .A2(G34), .ZN(new_n728));
  NAND2_X1  g303(.A1(KEYINPUT24), .A2(G34), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n728), .A2(new_n708), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G160), .B2(new_n708), .ZN(new_n731));
  INV_X1    g306(.A(G2084), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n485), .A2(G141), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT96), .Z(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT26), .Z(new_n737));
  NAND3_X1  g312(.A1(new_n470), .A2(G105), .A3(G2104), .ZN(new_n738));
  INV_X1    g313(.A(G129), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n737), .B(new_n738), .C1(new_n481), .C2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G29), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G29), .B2(G32), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT27), .B(G1996), .ZN(new_n744));
  OAI22_X1  g319(.A1(new_n743), .A2(new_n744), .B1(new_n717), .B2(G2072), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n708), .A2(G35), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G162), .B2(new_n708), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT29), .B(G2090), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  AND4_X1   g325(.A1(new_n718), .A2(new_n727), .A3(new_n733), .A4(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n708), .B1(new_n752), .B2(G28), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(KEYINPUT98), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(G28), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(KEYINPUT98), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT31), .B(G11), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n757), .B(new_n758), .C1(new_n651), .C2(new_n708), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT99), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n720), .A2(G21), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G168), .B2(new_n720), .ZN(new_n762));
  INV_X1    g337(.A(G1966), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G5), .A2(G16), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G171), .B2(G16), .ZN(new_n766));
  INV_X1    g341(.A(G1961), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT28), .ZN(new_n770));
  INV_X1    g345(.A(G26), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(G29), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(G29), .ZN(new_n773));
  AOI22_X1  g348(.A1(G128), .A2(new_n482), .B1(new_n485), .B2(G140), .ZN(new_n774));
  OAI221_X1 g349(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n474), .C2(G116), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n773), .B1(new_n776), .B2(G29), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n772), .B1(new_n777), .B2(new_n770), .ZN(new_n778));
  AOI211_X1 g353(.A(new_n760), .B(new_n769), .C1(G2067), .C2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G19), .ZN(new_n780));
  OAI21_X1  g355(.A(KEYINPUT95), .B1(new_n780), .B2(G16), .ZN(new_n781));
  OR3_X1    g356(.A1(new_n780), .A2(KEYINPUT95), .A3(G16), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n781), .B(new_n782), .C1(new_n575), .C2(new_n720), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G1341), .Z(new_n784));
  OR2_X1    g359(.A1(new_n778), .A2(G2067), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n751), .A2(new_n779), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT34), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n720), .A2(G22), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G303), .B2(G16), .ZN(new_n790));
  INV_X1    g365(.A(G1971), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n603), .A2(new_n604), .A3(G16), .A4(new_n605), .ZN(new_n794));
  OR2_X1    g369(.A1(G6), .A2(G16), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(KEYINPUT32), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT32), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n794), .A2(new_n798), .A3(new_n795), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n797), .A2(G1981), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n797), .A2(new_n799), .ZN(new_n801));
  INV_X1    g376(.A(G1981), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n792), .A2(new_n793), .A3(new_n800), .A4(new_n803), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n720), .A2(G23), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G288), .B2(G16), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT33), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  AOI211_X1 g384(.A(KEYINPUT33), .B(new_n805), .C1(G288), .C2(G16), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n809), .A2(G1976), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G1976), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n808), .B2(new_n810), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n787), .B1(new_n804), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n812), .A2(new_n814), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n790), .B(G1971), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n803), .A2(new_n800), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n817), .A2(new_n818), .A3(new_n819), .A4(KEYINPUT34), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n720), .A2(G24), .ZN(new_n822));
  INV_X1    g397(.A(G290), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(new_n720), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(G1986), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(G1986), .ZN(new_n826));
  AOI22_X1  g401(.A1(G119), .A2(new_n482), .B1(new_n485), .B2(G131), .ZN(new_n827));
  OAI221_X1 g402(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n474), .C2(G107), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  MUX2_X1   g404(.A(G25), .B(new_n829), .S(G29), .Z(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT35), .B(G1991), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n830), .B(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n825), .A2(new_n826), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n821), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT93), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT93), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n821), .A2(new_n838), .A3(new_n835), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n837), .A2(KEYINPUT36), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT36), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n838), .B1(new_n821), .B2(new_n835), .ZN(new_n842));
  AOI211_X1 g417(.A(KEYINPUT93), .B(new_n834), .C1(new_n816), .C2(new_n820), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n786), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n743), .A2(new_n744), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT97), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n708), .A2(G27), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(G164), .B2(new_n708), .ZN(new_n849));
  INV_X1    g424(.A(G2078), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(G4), .A2(G16), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(new_n623), .B2(G16), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT94), .ZN(new_n854));
  INV_X1    g429(.A(G1348), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n845), .A2(new_n847), .A3(new_n851), .A4(new_n856), .ZN(G150));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n858));
  NAND2_X1  g433(.A1(G150), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n856), .ZN(new_n860));
  AOI211_X1 g435(.A(new_n860), .B(new_n786), .C1(new_n840), .C2(new_n844), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n861), .A2(KEYINPUT101), .A3(new_n847), .A4(new_n851), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(G311));
  AND2_X1   g438(.A1(new_n543), .A2(G93), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n535), .A2(G55), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT102), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n867), .B2(new_n508), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n869), .A2(new_n630), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT104), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT37), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n623), .A2(G559), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT39), .ZN(new_n874));
  XNOR2_X1  g449(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n869), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n573), .B1(new_n572), .B2(new_n559), .ZN(new_n878));
  AOI211_X1 g453(.A(KEYINPUT80), .B(new_n558), .C1(new_n570), .C2(new_n571), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n564), .A2(new_n869), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n876), .B(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n872), .B1(new_n883), .B2(G860), .ZN(G145));
  NAND2_X1  g459(.A1(new_n495), .A2(new_n500), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n492), .A2(new_n887), .A3(new_n493), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n887), .B1(new_n492), .B2(new_n493), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n776), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n716), .A2(KEYINPUT106), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n741), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  AOI22_X1  g470(.A1(G130), .A2(new_n482), .B1(new_n485), .B2(G142), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n474), .A2(G118), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT107), .ZN(new_n898));
  OAI21_X1  g473(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n639), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(new_n829), .Z(new_n902));
  XOR2_X1   g477(.A(new_n895), .B(new_n902), .Z(new_n903));
  XNOR2_X1  g478(.A(new_n651), .B(G160), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(G162), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G37), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n895), .B(new_n909), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n906), .B(new_n907), .C1(new_n905), .C2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g487(.A1(new_n877), .A2(new_n626), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n622), .A2(G299), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n622), .A2(G299), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n915), .B2(new_n916), .ZN(new_n919));
  INV_X1    g494(.A(new_n916), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n920), .A2(KEYINPUT41), .A3(new_n914), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n882), .B(new_n634), .ZN(new_n924));
  MUX2_X1   g499(.A(new_n917), .B(new_n923), .S(new_n924), .Z(new_n925));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n926));
  INV_X1    g501(.A(G288), .ZN(new_n927));
  NAND2_X1  g502(.A1(G303), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n518), .B(G288), .C1(new_n537), .C2(new_n538), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n928), .A2(G290), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(G290), .B1(new_n928), .B2(new_n929), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n930), .A2(new_n931), .A3(G305), .ZN(new_n932));
  INV_X1    g507(.A(G305), .ZN(new_n933));
  INV_X1    g508(.A(new_n929), .ZN(new_n934));
  INV_X1    g509(.A(G88), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n541), .A2(new_n542), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n536), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT77), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(G288), .B1(new_n940), .B2(new_n518), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n823), .B1(new_n934), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n928), .A2(G290), .A3(new_n929), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n933), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n926), .B1(new_n932), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(G305), .B1(new_n930), .B2(new_n931), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(new_n933), .A3(new_n943), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n946), .A2(KEYINPUT109), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT109), .B1(new_n946), .B2(new_n947), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n945), .B1(new_n950), .B2(new_n926), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n925), .B(new_n951), .Z(new_n952));
  OAI21_X1  g527(.A(new_n913), .B1(new_n952), .B2(new_n626), .ZN(G295));
  OAI21_X1  g528(.A(new_n913), .B1(new_n952), .B2(new_n626), .ZN(G331));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n869), .B1(new_n565), .B2(new_n574), .ZN(new_n956));
  XNOR2_X1  g531(.A(G286), .B(G171), .ZN(new_n957));
  INV_X1    g532(.A(new_n881), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(G286), .B(G301), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n880), .B2(new_n881), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n923), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n959), .A2(new_n961), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n962), .A2(KEYINPUT110), .B1(new_n963), .B2(new_n917), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n957), .B1(new_n956), .B2(new_n958), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n880), .A2(new_n881), .A3(new_n960), .ZN(new_n966));
  AOI211_X1 g541(.A(KEYINPUT110), .B(new_n922), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n964), .A2(new_n950), .A3(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n965), .A2(new_n917), .A3(new_n966), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n922), .B1(new_n965), .B2(new_n966), .ZN(new_n971));
  OAI22_X1  g546(.A1(new_n948), .A2(new_n949), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n907), .B1(new_n972), .B2(new_n973), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT113), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n932), .B2(new_n944), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n946), .A2(KEYINPUT109), .A3(new_n947), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n965), .A2(new_n966), .A3(new_n917), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n979), .A2(new_n980), .B1(new_n962), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(G37), .B1(new_n982), .B2(KEYINPUT112), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n983), .A2(new_n984), .A3(new_n974), .A4(new_n969), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n955), .B1(new_n977), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n979), .A2(new_n980), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n981), .B1(new_n971), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n987), .B1(new_n989), .B2(new_n967), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n969), .A2(new_n907), .A3(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n991), .A2(new_n955), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT44), .B1(new_n986), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT111), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n983), .A2(new_n955), .A3(new_n974), .A4(new_n969), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n991), .A2(new_n997), .A3(KEYINPUT43), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n993), .A2(new_n1001), .ZN(G397));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n890), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  AND2_X1   g580(.A1(G160), .A2(G40), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1996), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n1011), .A2(new_n1012), .A3(new_n741), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  INV_X1    g591(.A(G2067), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n776), .B(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n741), .A2(new_n1012), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1011), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1015), .A2(new_n1016), .A3(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n829), .B(new_n832), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1021), .B1(new_n1011), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1011), .ZN(new_n1024));
  XNOR2_X1  g599(.A(G290), .B(G1986), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1006), .A2(new_n890), .A3(new_n1003), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1027), .A2(G8), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G288), .A2(new_n813), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT52), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G305), .A2(G1981), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(G305), .A2(G1981), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1032), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1035), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(KEYINPUT49), .A3(new_n1033), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1036), .A2(new_n1038), .A3(new_n1028), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT52), .B1(G288), .B2(new_n813), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1028), .B(new_n1040), .C1(new_n813), .C2(G288), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1031), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n890), .A2(KEYINPUT45), .A3(new_n1003), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n495), .A2(KEYINPUT72), .A3(new_n500), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(new_n501), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1003), .B1(new_n1045), .B2(new_n494), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n1005), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1047), .A3(new_n1006), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n791), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1006), .B1(new_n1046), .B2(KEYINPUT50), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1051), .B1(new_n890), .B2(new_n1003), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1049), .B1(new_n1053), .B2(G2090), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G303), .A2(G8), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT55), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n1057));
  NAND3_X1  g632(.A1(G303), .A2(new_n1057), .A3(G8), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1054), .A2(G8), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1042), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n890), .A2(new_n1051), .A3(new_n1003), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1006), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1049), .B1(G2090), .B2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1064), .A2(G8), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1060), .A2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT58), .B(G1341), .Z(new_n1067));
  NAND2_X1  g642(.A1(new_n1027), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n1048), .B2(G1996), .ZN(new_n1069));
  AND2_X1   g644(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n575), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1070), .B1(new_n575), .B2(new_n1069), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1027), .A2(G2067), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1075), .A2(new_n1076), .B1(new_n1063), .B2(new_n855), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT120), .B1(new_n1027), .B2(G2067), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n622), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1076), .A2(new_n1075), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1063), .A2(new_n855), .ZN(new_n1081));
  AND4_X1   g656(.A1(new_n622), .A2(new_n1080), .A3(new_n1081), .A4(new_n1078), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT60), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n1084));
  AND4_X1   g659(.A1(new_n1084), .A2(new_n1080), .A3(new_n1081), .A4(new_n1078), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n582), .A2(new_n584), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n588), .A2(new_n587), .ZN(new_n1087));
  NAND2_X1  g662(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1088));
  OR2_X1    g663(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(G299), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n1094));
  INV_X1    g669(.A(G1956), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1043), .A2(new_n1047), .A3(new_n1006), .A4(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1093), .A2(new_n1094), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1085), .A2(new_n623), .B1(new_n1099), .B2(KEYINPUT61), .ZN(new_n1100));
  NOR2_X1   g675(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1093), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(new_n1092), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1101), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1074), .A2(new_n1083), .A3(new_n1100), .A4(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1092), .B(KEYINPUT121), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1103), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1079), .B1(new_n1103), .B2(new_n1092), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1048), .B2(G2078), .ZN(new_n1112));
  NAND2_X1  g687(.A1(G160), .A2(G40), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1046), .A2(new_n1005), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1114), .A2(KEYINPUT53), .A3(new_n850), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1063), .A2(new_n767), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1112), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(G171), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1114), .A2(KEYINPUT53), .A3(new_n850), .A4(new_n1043), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1112), .A2(new_n1122), .A3(G301), .A4(new_n1117), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1118), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT54), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1121), .A2(new_n1125), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1118), .A2(G301), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1112), .A2(new_n1122), .A3(new_n1117), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1129), .B(KEYINPUT54), .C1(G301), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT51), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n763), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1063), .A2(G2084), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(G8), .B(new_n1135), .C1(new_n1139), .C2(G286), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1135), .ZN(new_n1141));
  NAND2_X1  g716(.A1(G286), .A2(G8), .ZN(new_n1142));
  AOI21_X1  g717(.A(G1966), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1063), .A2(G2084), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(G8), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1141), .B(new_n1142), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1140), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1139), .A2(G8), .A3(G286), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1110), .A2(new_n1132), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(KEYINPUT62), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1149), .A2(new_n1155), .A3(new_n1150), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1153), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1066), .B1(new_n1152), .B2(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1031), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1054), .A2(G8), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1145), .A2(new_n1146), .A3(G286), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1159), .A2(new_n1162), .A3(new_n1163), .A4(new_n1065), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT118), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT118), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1060), .A2(new_n1166), .A3(new_n1065), .A4(new_n1163), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT63), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT116), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1042), .B(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1064), .A2(G8), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1168), .B1(new_n1172), .B2(new_n1161), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1171), .A2(new_n1065), .A3(new_n1163), .A4(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1169), .A2(new_n1174), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1028), .B(KEYINPUT117), .Z(new_n1176));
  AND3_X1   g751(.A1(new_n1039), .A2(new_n813), .A3(new_n927), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1176), .B1(new_n1177), .B2(new_n1035), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1065), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1171), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1175), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1026), .B1(new_n1158), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(KEYINPUT127), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1184), .B(new_n1026), .C1(new_n1158), .C2(new_n1181), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1021), .A2(new_n832), .A3(new_n827), .A4(new_n828), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n774), .A2(new_n1017), .A3(new_n775), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1011), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n1011), .A2(G1986), .A3(G290), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT48), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1023), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1011), .B1(new_n741), .B2(new_n1018), .ZN(new_n1193));
  OR3_X1    g768(.A1(new_n1011), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1194));
  OAI21_X1  g769(.A(KEYINPUT46), .B1(new_n1011), .B2(G1996), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT47), .ZN(new_n1197));
  NOR3_X1   g772(.A1(new_n1189), .A2(new_n1192), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1186), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g774(.A(G229), .ZN(new_n1201));
  AND3_X1   g775(.A1(new_n911), .A2(G319), .A3(new_n667), .ZN(new_n1202));
  AND4_X1   g776(.A1(new_n686), .A2(new_n999), .A3(new_n1201), .A4(new_n1202), .ZN(G308));
  NAND4_X1  g777(.A1(new_n999), .A2(new_n686), .A3(new_n1201), .A4(new_n1202), .ZN(G225));
endmodule


