//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1027, new_n1028, new_n1029;
  XNOR2_X1  g000(.A(KEYINPUT88), .B(G29gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G36gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT89), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT89), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n202), .A2(new_n205), .A3(G36gat), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT14), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT14), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n204), .A2(new_n206), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  INV_X1    g014(.A(G43gat), .ZN(new_n216));
  INV_X1    g015(.A(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G43gat), .A2(G50gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n215), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n212), .A2(KEYINPUT90), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT90), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n211), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n218), .A2(new_n215), .A3(new_n219), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n223), .A2(new_n221), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI22_X1  g026(.A1(new_n214), .A2(new_n221), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(G15gat), .B(G22gat), .Z(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT91), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT92), .ZN(new_n232));
  XNOR2_X1  g031(.A(G15gat), .B(G22gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT91), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G1gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT16), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n231), .A2(new_n239), .A3(new_n235), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n231), .A2(new_n232), .A3(G1gat), .A4(new_n235), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n238), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G8gat), .ZN(new_n243));
  INV_X1    g042(.A(G8gat), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n238), .A2(new_n240), .A3(new_n244), .A4(new_n241), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n229), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT18), .ZN(new_n247));
  NAND2_X1  g046(.A1(G229gat), .A2(G233gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n246), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT17), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n228), .A2(new_n251), .ZN(new_n252));
  OAI221_X1 g051(.A(KEYINPUT17), .B1(new_n222), .B2(new_n227), .C1(new_n214), .C2(new_n221), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n252), .A2(new_n243), .A3(new_n253), .A4(new_n245), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT93), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n254), .A2(new_n255), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n250), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n243), .A2(new_n245), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n229), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n228), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n248), .B(KEYINPUT13), .Z(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n259), .A2(KEYINPUT93), .A3(new_n252), .A4(new_n253), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n255), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n246), .A2(new_n249), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G113gat), .B(G141gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT11), .ZN(new_n275));
  INV_X1    g074(.A(G169gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(G197gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT12), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n266), .A2(new_n273), .A3(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n272), .B1(new_n256), .B2(new_n257), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n267), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n271), .A2(new_n250), .B1(new_n263), .B2(new_n264), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n279), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT36), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT68), .B(G71gat), .ZN(new_n288));
  INV_X1    g087(.A(G99gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G15gat), .B(G43gat), .Z(new_n291));
  XOR2_X1   g090(.A(new_n290), .B(new_n291), .Z(new_n292));
  NAND2_X1  g091(.A1(G227gat), .A2(G233gat), .ZN(new_n293));
  INV_X1    g092(.A(G120gat), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT66), .B1(new_n294), .B2(G113gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n296));
  INV_X1    g095(.A(G113gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n296), .A2(new_n297), .A3(G120gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(G113gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n295), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G134gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G127gat), .ZN(new_n302));
  INV_X1    g101(.A(G127gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G134gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT1), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n297), .A2(G120gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n294), .A2(G113gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n302), .A2(new_n304), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n300), .A2(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT27), .B(G183gat), .ZN(new_n312));
  INV_X1    g111(.A(G190gat), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT28), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G183gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT27), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT27), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G183gat), .ZN(new_n318));
  AND4_X1   g117(.A1(KEYINPUT28), .A2(new_n316), .A3(new_n318), .A4(new_n313), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR3_X1   g123(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT65), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n316), .A2(new_n318), .A3(new_n313), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n312), .A2(KEYINPUT28), .A3(new_n313), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n326), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT65), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT24), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n315), .A2(new_n313), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G176gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n276), .A2(new_n343), .A3(KEYINPUT23), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(G169gat), .B2(G176gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n346), .A3(new_n323), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n336), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n344), .A2(new_n346), .A3(new_n323), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT64), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n339), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n351), .A2(new_n340), .A3(new_n338), .A4(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n349), .A2(new_n353), .A3(KEYINPUT25), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  AND4_X1   g154(.A1(new_n311), .A2(new_n327), .A3(new_n335), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n309), .A2(new_n310), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n306), .A2(new_n300), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n326), .B1(new_n330), .B2(new_n331), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n344), .A2(new_n346), .A3(KEYINPUT25), .A4(new_n323), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n351), .A2(new_n340), .A3(new_n338), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n361), .B1(new_n362), .B2(new_n352), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT25), .B1(new_n349), .B2(new_n341), .ZN(new_n364));
  OAI22_X1  g163(.A1(new_n360), .A2(new_n334), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n335), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n359), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n356), .B1(KEYINPUT67), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT67), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n369), .B(new_n359), .C1(new_n365), .C2(new_n366), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n293), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n292), .B1(new_n371), .B2(KEYINPUT33), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n367), .A2(KEYINPUT67), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n332), .A2(new_n333), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n374), .A2(KEYINPUT65), .B1(new_n348), .B2(new_n354), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(new_n311), .A3(new_n335), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n373), .A2(new_n370), .A3(new_n293), .A4(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT69), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT34), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT34), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n377), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n372), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n292), .ZN(new_n384));
  INV_X1    g183(.A(new_n293), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n311), .B1(new_n375), .B2(new_n335), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n376), .B1(new_n386), .B2(new_n369), .ZN(new_n387));
  INV_X1    g186(.A(new_n370), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT33), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n384), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n377), .A2(new_n378), .A3(new_n381), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n381), .B1(new_n377), .B2(new_n378), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n389), .A2(KEYINPUT32), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n383), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n396), .B1(new_n383), .B2(new_n394), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n287), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n394), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n395), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n394), .A3(new_n396), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(KEYINPUT36), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n405));
  AND2_X1   g204(.A1(G141gat), .A2(G148gat), .ZN(new_n406));
  NOR2_X1   g205(.A1(G141gat), .A2(G148gat), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT73), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(G141gat), .ZN(new_n409));
  INV_X1    g208(.A(G148gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT73), .ZN(new_n412));
  NAND2_X1  g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT2), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n408), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(G155gat), .A2(G162gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(G155gat), .A2(G162gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT74), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n420), .B1(new_n417), .B2(new_n418), .ZN(new_n421));
  INV_X1    g220(.A(G155gat), .ZN(new_n422));
  INV_X1    g221(.A(G162gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G155gat), .A2(G162gat), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(KEYINPUT74), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G141gat), .B(G148gat), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n415), .B1(G155gat), .B2(G162gat), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n416), .A2(new_n419), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT3), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT29), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(G211gat), .B(G218gat), .Z(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(G211gat), .A2(G218gat), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT22), .ZN(new_n437));
  INV_X1    g236(.A(G197gat), .ZN(new_n438));
  INV_X1    g237(.A(G204gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G197gat), .A2(G204gat), .ZN(new_n441));
  AOI221_X4 g240(.A(KEYINPUT70), .B1(new_n436), .B2(new_n437), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT70), .ZN(new_n443));
  XNOR2_X1  g242(.A(G197gat), .B(G204gat), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n443), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n435), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(G197gat), .A2(G204gat), .ZN(new_n449));
  NOR2_X1   g248(.A1(G197gat), .A2(G204gat), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT70), .B1(new_n451), .B2(new_n445), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n444), .A2(new_n443), .A3(new_n446), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n434), .A3(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT77), .B1(new_n433), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT29), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n448), .A2(new_n457), .A3(new_n454), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n432), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n416), .A2(new_n419), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n427), .A2(new_n430), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n432), .A3(new_n461), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n457), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT77), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n448), .A2(new_n454), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n456), .A2(new_n463), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(G228gat), .A2(G233gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(G22gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n465), .A2(new_n467), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT78), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n470), .B1(new_n459), .B2(new_n462), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT78), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n465), .A2(new_n476), .A3(new_n467), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n471), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT80), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n473), .A2(KEYINPUT77), .B1(new_n459), .B2(new_n462), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n481), .A2(new_n468), .B1(G228gat), .B2(G233gat), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n483));
  OAI21_X1  g282(.A(G22gat), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G78gat), .B(G106gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT31), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(new_n217), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n471), .A2(new_n472), .A3(new_n478), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT80), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n480), .A2(new_n484), .A3(new_n488), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n484), .A2(new_n489), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT79), .B1(new_n493), .B2(new_n487), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT79), .ZN(new_n495));
  AOI211_X1 g294(.A(new_n495), .B(new_n488), .C1(new_n484), .C2(new_n489), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n405), .B(new_n492), .C1(new_n494), .C2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n472), .B1(new_n471), .B2(new_n478), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n487), .B1(new_n479), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n495), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n493), .A2(KEYINPUT79), .A3(new_n487), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n405), .B1(new_n503), .B2(new_n492), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G8gat), .B(G36gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(G64gat), .ZN(new_n507));
  INV_X1    g306(.A(G92gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G226gat), .ZN(new_n510));
  INV_X1    g309(.A(G233gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT71), .B1(new_n365), .B2(new_n366), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT71), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n327), .A2(new_n515), .A3(new_n335), .A4(new_n355), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n513), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n360), .B1(new_n348), .B2(new_n354), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n518), .A2(KEYINPUT29), .A3(new_n512), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n517), .A2(new_n467), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n512), .A2(KEYINPUT29), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n514), .A2(new_n516), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n518), .A2(new_n512), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n455), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n509), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT72), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT30), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n520), .ZN(new_n531));
  INV_X1    g330(.A(new_n524), .ZN(new_n532));
  INV_X1    g331(.A(new_n509), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT5), .ZN(new_n537));
  INV_X1    g336(.A(new_n419), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT2), .B1(new_n428), .B2(KEYINPUT73), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(new_n414), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n411), .B(new_n413), .C1(new_n417), .C2(new_n415), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n541), .B1(new_n421), .B2(new_n426), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n359), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n311), .A2(new_n460), .A3(new_n461), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G225gat), .A2(G233gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT75), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n537), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(KEYINPUT4), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n431), .A2(KEYINPUT4), .A3(new_n311), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n464), .A2(new_n359), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n431), .A2(new_n432), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n551), .B(new_n552), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(new_n359), .A3(new_n464), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT4), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n548), .A2(KEYINPUT5), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n558), .A2(new_n552), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G57gat), .B(G85gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(G1gat), .B(G29gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT6), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n562), .A3(new_n568), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n563), .A2(KEYINPUT6), .A3(new_n569), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n536), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n404), .B1(new_n505), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n503), .A2(new_n492), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n560), .B(new_n552), .C1(new_n553), .C2(new_n554), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT82), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n580), .A2(new_n581), .A3(new_n548), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n580), .B2(new_n548), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n584), .B(KEYINPUT39), .C1(new_n548), .C2(new_n545), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT83), .B(KEYINPUT39), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(new_n582), .B2(new_n583), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n587), .A2(KEYINPUT84), .A3(new_n568), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT84), .B1(new_n587), .B2(new_n568), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT40), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(KEYINPUT40), .B(new_n585), .C1(new_n588), .C2(new_n589), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n592), .A2(new_n535), .A3(new_n570), .A4(new_n593), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n573), .A2(new_n574), .A3(new_n525), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT86), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT85), .B(KEYINPUT37), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(new_n520), .B2(new_n524), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n467), .B1(new_n517), .B2(new_n519), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n522), .A2(new_n523), .A3(new_n455), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(KEYINPUT37), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT38), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n598), .A2(new_n601), .A3(new_n602), .A4(new_n533), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n595), .A2(new_n596), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n596), .B1(new_n595), .B2(new_n603), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n531), .A2(KEYINPUT37), .A3(new_n532), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n607), .A2(new_n598), .A3(new_n533), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT38), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT87), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT87), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n608), .A2(new_n611), .A3(KEYINPUT38), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n579), .B(new_n594), .C1(new_n606), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n578), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n535), .A2(new_n575), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n401), .A2(new_n402), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n617), .A3(new_n579), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT35), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT35), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n616), .A2(new_n617), .A3(new_n620), .A4(new_n579), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n286), .B1(new_n615), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n625));
  AND2_X1   g424(.A1(G71gat), .A2(G78gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(G71gat), .A2(G78gat), .ZN(new_n627));
  OAI22_X1  g426(.A1(new_n624), .A2(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(G57gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(G64gat), .ZN(new_n630));
  INV_X1    g429(.A(G64gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(G57gat), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n624), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n628), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(KEYINPUT21), .ZN(new_n637));
  XOR2_X1   g436(.A(G127gat), .B(G155gat), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G211gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(KEYINPUT21), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n243), .A2(new_n245), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(G183gat), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n243), .A2(new_n315), .A3(new_n245), .A4(new_n641), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n645));
  NAND2_X1  g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n643), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n643), .B2(new_n644), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n640), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n643), .A2(new_n644), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n647), .ZN(new_n653));
  INV_X1    g452(.A(G211gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n639), .B(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n643), .A2(new_n644), .A3(new_n648), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n653), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G134gat), .B(G162gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT96), .ZN(new_n660));
  NAND2_X1  g459(.A1(G232gat), .A2(G233gat), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n660), .B(new_n663), .Z(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(G85gat), .A2(G92gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT7), .ZN(new_n667));
  NAND2_X1  g466(.A1(G99gat), .A2(G106gat), .ZN(new_n668));
  INV_X1    g467(.A(G85gat), .ZN(new_n669));
  AOI22_X1  g468(.A1(KEYINPUT8), .A2(new_n668), .B1(new_n669), .B2(new_n508), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(G99gat), .B(G106gat), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n672), .B1(new_n667), .B2(new_n670), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n252), .A2(new_n253), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(G190gat), .B(G218gat), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT97), .ZN(new_n681));
  OAI22_X1  g480(.A1(new_n680), .A2(KEYINPUT97), .B1(new_n662), .B2(new_n661), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n228), .B2(new_n676), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n678), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n681), .B1(new_n678), .B2(new_n683), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n665), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n678), .A2(new_n683), .ZN(new_n687));
  INV_X1    g486(.A(new_n681), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n678), .A2(new_n681), .A3(new_n683), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(new_n664), .A3(new_n690), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n658), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT98), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT98), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n658), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(G230gat), .A2(G233gat), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n672), .A2(KEYINPUT99), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n671), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n671), .A2(new_n701), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n636), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n635), .B(new_n634), .C1(new_n674), .C2(new_n675), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT10), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n676), .A2(KEYINPUT10), .A3(new_n636), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n700), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n704), .A2(new_n705), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n700), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(G120gat), .B(G148gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G176gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(new_n439), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n711), .A2(new_n714), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n698), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n623), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n576), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(new_n237), .ZN(G1324gat));
  NAND3_X1  g520(.A1(new_n623), .A2(new_n535), .A3(new_n718), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT100), .B(KEYINPUT16), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(new_n244), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n725), .A2(KEYINPUT42), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(KEYINPUT42), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n722), .A2(G8gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(G1325gat));
  AND2_X1   g528(.A1(new_n399), .A2(new_n403), .ZN(new_n730));
  OAI21_X1  g529(.A(G15gat), .B1(new_n719), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n617), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n732), .A2(G15gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n719), .B2(new_n733), .ZN(G1326gat));
  INV_X1    g533(.A(new_n505), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n719), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT43), .B(G22gat), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1327gat));
  INV_X1    g537(.A(new_n692), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n579), .A2(KEYINPUT81), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(new_n577), .A3(new_n497), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n614), .A2(KEYINPUT101), .A3(new_n741), .A4(new_n730), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n622), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT101), .B1(new_n578), .B2(new_n614), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n739), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n615), .A2(new_n622), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n748), .A2(KEYINPUT44), .A3(new_n739), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n280), .B1(new_n266), .B2(new_n273), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n283), .A2(new_n279), .A3(new_n284), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n658), .ZN(new_n754));
  INV_X1    g553(.A(new_n717), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n750), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n202), .B1(new_n758), .B2(new_n576), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n658), .A2(new_n692), .A3(new_n717), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n623), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n761), .A2(new_n576), .A3(new_n202), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT45), .Z(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n763), .ZN(G1328gat));
  OAI21_X1  g563(.A(G36gat), .B1(new_n758), .B2(new_n536), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n761), .A2(G36gat), .A3(new_n536), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT46), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1329gat));
  NOR2_X1   g567(.A1(new_n730), .A2(new_n216), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n757), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n623), .A2(new_n617), .A3(new_n760), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT102), .B1(new_n771), .B2(new_n216), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n770), .A2(KEYINPUT47), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT47), .B1(new_n770), .B2(new_n772), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(G1330gat));
  NAND4_X1  g574(.A1(new_n623), .A2(new_n217), .A3(new_n505), .A4(new_n760), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n757), .A2(new_n505), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(G50gat), .ZN(new_n779));
  INV_X1    g578(.A(new_n579), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n217), .B1(new_n757), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n776), .A2(KEYINPUT48), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n779), .A2(KEYINPUT48), .B1(new_n781), .B2(new_n782), .ZN(G1331gat));
  OR2_X1    g582(.A1(new_n743), .A2(new_n744), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n698), .A2(new_n753), .A3(new_n755), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n575), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g588(.A(new_n536), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n792));
  XOR2_X1   g591(.A(new_n791), .B(new_n792), .Z(G1333gat));
  OAI21_X1  g592(.A(G71gat), .B1(new_n786), .B2(new_n730), .ZN(new_n794));
  INV_X1    g593(.A(G71gat), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n617), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n786), .B2(new_n796), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n797), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g597(.A1(new_n787), .A2(new_n505), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g599(.A1(new_n753), .A2(new_n658), .A3(new_n755), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n747), .A2(new_n749), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT103), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n747), .A2(KEYINPUT103), .A3(new_n749), .A4(new_n801), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n805), .A2(new_n807), .A3(new_n576), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n753), .A2(new_n658), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n784), .A2(KEYINPUT51), .A3(new_n739), .A4(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n811));
  INV_X1    g610(.A(new_n809), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n745), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n717), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n575), .A2(new_n669), .ZN(new_n816));
  OAI22_X1  g615(.A1(new_n808), .A2(new_n669), .B1(new_n815), .B2(new_n816), .ZN(G1336gat));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n818), .B(G92gat), .C1(new_n802), .C2(new_n536), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n535), .A2(new_n508), .A3(new_n717), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT104), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n814), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n819), .B(new_n823), .C1(KEYINPUT105), .C2(new_n818), .ZN(new_n824));
  AOI211_X1 g623(.A(KEYINPUT105), .B(new_n821), .C1(new_n810), .C2(new_n813), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n804), .A2(new_n535), .A3(new_n806), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n826), .B2(G92gat), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n824), .B1(new_n827), .B2(new_n818), .ZN(G1337gat));
  NOR3_X1   g627(.A1(new_n805), .A2(new_n807), .A3(new_n730), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n617), .A2(new_n289), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n829), .A2(new_n289), .B1(new_n815), .B2(new_n830), .ZN(G1338gat));
  OR3_X1    g630(.A1(new_n579), .A2(G106gat), .A3(new_n755), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT106), .Z(new_n833));
  NAND3_X1  g632(.A1(new_n814), .A2(KEYINPUT107), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G106gat), .B1(new_n802), .B2(new_n579), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT53), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n804), .A2(new_n505), .A3(new_n806), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(KEYINPUT53), .A3(G106gat), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n814), .A2(new_n833), .B1(KEYINPUT107), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n836), .B1(new_n838), .B2(new_n840), .ZN(G1339gat));
  NAND2_X1  g640(.A1(new_n707), .A2(new_n708), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n699), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n707), .A2(new_n700), .A3(new_n708), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(KEYINPUT54), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n714), .B1(new_n709), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(KEYINPUT55), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n716), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT55), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n845), .A2(new_n847), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n753), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n248), .B1(new_n271), .B2(new_n262), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n263), .A2(new_n264), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n278), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n752), .A2(new_n856), .A3(new_n717), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n739), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n752), .A2(new_n856), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n739), .A3(new_n852), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n754), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n286), .A2(new_n694), .A3(new_n696), .A4(new_n755), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n505), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n535), .A2(new_n576), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n617), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n867), .A2(new_n297), .A3(new_n286), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n864), .A2(new_n576), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n732), .A2(new_n780), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT108), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n536), .A3(new_n753), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n868), .B1(new_n873), .B2(new_n297), .ZN(G1340gat));
  NOR3_X1   g673(.A1(new_n867), .A2(new_n294), .A3(new_n755), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n872), .A2(new_n536), .A3(new_n717), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(new_n294), .ZN(G1341gat));
  OAI21_X1  g676(.A(G127gat), .B1(new_n867), .B2(new_n754), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n872), .A2(new_n536), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n658), .A2(new_n303), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(G1342gat));
  NOR2_X1   g680(.A1(new_n692), .A2(G134gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n872), .A2(new_n536), .A3(new_n882), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n884));
  OAI21_X1  g683(.A(G134gat), .B1(new_n867), .B2(new_n692), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(G1343gat));
  INV_X1    g686(.A(new_n863), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT112), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT110), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT55), .B1(new_n851), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT111), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n845), .A2(KEYINPUT110), .A3(new_n847), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n892), .B1(new_n891), .B2(new_n893), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n849), .B1(new_n751), .B2(new_n752), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n896), .A2(new_n897), .B1(new_n859), .B2(new_n717), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n889), .B1(new_n898), .B2(new_n739), .ZN(new_n899));
  INV_X1    g698(.A(new_n849), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n900), .B1(new_n281), .B2(new_n285), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n851), .A2(new_n890), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n850), .A3(new_n893), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT111), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n857), .B1(new_n901), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(KEYINPUT112), .A3(new_n692), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n899), .A2(new_n860), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n888), .B1(new_n909), .B2(new_n754), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n735), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT113), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT113), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n907), .A2(new_n692), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n861), .B1(new_n916), .B2(new_n889), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n658), .B1(new_n917), .B2(new_n908), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n915), .B(new_n912), .C1(new_n918), .C2(new_n888), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n911), .B1(new_n864), .B2(new_n579), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n914), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n730), .A2(new_n866), .ZN(new_n922));
  XOR2_X1   g721(.A(new_n922), .B(KEYINPUT109), .Z(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n753), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G141gat), .ZN(new_n925));
  AND4_X1   g724(.A1(new_n536), .A2(new_n869), .A3(new_n780), .A4(new_n730), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n753), .A2(new_n409), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT114), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT115), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n931), .A2(KEYINPUT58), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(KEYINPUT58), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT116), .Z(new_n935));
  NAND3_X1  g734(.A1(new_n930), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n935), .ZN(new_n937));
  AOI22_X1  g736(.A1(new_n924), .A2(G141gat), .B1(new_n926), .B2(new_n928), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n932), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n939), .ZN(G1344gat));
  NAND3_X1  g739(.A1(new_n926), .A2(new_n410), .A3(new_n717), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT117), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n923), .A2(new_n717), .ZN(new_n944));
  AOI211_X1 g743(.A(new_n911), .B(new_n579), .C1(new_n862), .C2(new_n863), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n658), .B1(new_n916), .B2(new_n860), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n863), .B(KEYINPUT119), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n505), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n911), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n945), .B1(new_n949), .B2(KEYINPUT120), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT120), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n948), .A2(new_n951), .A3(new_n911), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n944), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n943), .B(KEYINPUT59), .C1(new_n953), .C2(new_n410), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n921), .A2(new_n717), .A3(new_n923), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT118), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n410), .A2(KEYINPUT59), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT119), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n863), .B(new_n959), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n753), .A2(new_n900), .A3(new_n905), .A4(new_n904), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n739), .B1(new_n961), .B2(new_n857), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n754), .B1(new_n962), .B2(new_n861), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n735), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(KEYINPUT120), .B1(new_n964), .B2(KEYINPUT57), .ZN(new_n965));
  INV_X1    g764(.A(new_n945), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n965), .A2(new_n952), .A3(new_n966), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n923), .A2(new_n717), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n410), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT59), .ZN(new_n970));
  OAI21_X1  g769(.A(KEYINPUT121), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n954), .A2(new_n958), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n956), .B1(new_n955), .B2(new_n957), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n942), .B1(new_n972), .B2(new_n973), .ZN(G1345gat));
  NAND2_X1  g773(.A1(new_n921), .A2(new_n923), .ZN(new_n975));
  OAI21_X1  g774(.A(G155gat), .B1(new_n975), .B2(new_n754), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n926), .A2(new_n422), .A3(new_n658), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1346gat));
  OAI21_X1  g777(.A(G162gat), .B1(new_n975), .B2(new_n692), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n926), .A2(new_n423), .A3(new_n739), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(G1347gat));
  NOR2_X1   g780(.A1(new_n864), .A2(new_n575), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n870), .A2(new_n535), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g785(.A(G169gat), .B1(new_n986), .B2(new_n753), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n865), .A2(new_n576), .A3(new_n535), .A4(new_n617), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n988), .A2(new_n276), .A3(new_n286), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n987), .A2(new_n989), .ZN(G1348gat));
  OAI21_X1  g789(.A(G176gat), .B1(new_n988), .B2(new_n755), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n717), .A2(new_n343), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n991), .B1(new_n985), .B2(new_n992), .ZN(G1349gat));
  OAI21_X1  g792(.A(G183gat), .B1(new_n988), .B2(new_n754), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n658), .A2(new_n312), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n994), .B1(new_n985), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n997));
  XOR2_X1   g796(.A(new_n996), .B(new_n997), .Z(G1350gat));
  OAI21_X1  g797(.A(G190gat), .B1(new_n988), .B2(new_n692), .ZN(new_n999));
  XOR2_X1   g798(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n1000));
  XNOR2_X1  g799(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n313), .A3(new_n739), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(G1351gat));
  NAND3_X1  g802(.A1(new_n730), .A2(new_n535), .A3(new_n780), .ZN(new_n1004));
  OR2_X1    g803(.A1(new_n1004), .A2(KEYINPUT124), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(KEYINPUT124), .ZN(new_n1006));
  AND3_X1   g805(.A1(new_n982), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  XOR2_X1   g806(.A(new_n1007), .B(KEYINPUT125), .Z(new_n1008));
  NAND3_X1  g807(.A1(new_n1008), .A2(new_n438), .A3(new_n753), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n404), .A2(new_n575), .A3(new_n536), .ZN(new_n1010));
  AND2_X1   g809(.A1(new_n967), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1011), .A2(KEYINPUT126), .A3(new_n753), .ZN(new_n1012));
  INV_X1    g811(.A(KEYINPUT126), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n967), .A2(new_n1010), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1013), .B1(new_n1014), .B2(new_n286), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1012), .A2(G197gat), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1009), .A2(new_n1016), .ZN(G1352gat));
  NAND3_X1  g816(.A1(new_n1007), .A2(new_n439), .A3(new_n717), .ZN(new_n1018));
  XOR2_X1   g817(.A(new_n1018), .B(KEYINPUT62), .Z(new_n1019));
  OAI21_X1  g818(.A(G204gat), .B1(new_n1014), .B2(new_n755), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1019), .A2(new_n1020), .ZN(G1353gat));
  NAND3_X1  g820(.A1(new_n1008), .A2(new_n654), .A3(new_n658), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1011), .A2(new_n658), .ZN(new_n1023));
  AND3_X1   g822(.A1(new_n1023), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1024));
  AOI21_X1  g823(.A(KEYINPUT63), .B1(new_n1023), .B2(G211gat), .ZN(new_n1025));
  OAI21_X1  g824(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(G1354gat));
  INV_X1    g825(.A(G218gat), .ZN(new_n1027));
  NOR3_X1   g826(.A1(new_n1014), .A2(new_n1027), .A3(new_n692), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1008), .A2(new_n739), .ZN(new_n1029));
  AOI21_X1  g828(.A(new_n1028), .B1(new_n1029), .B2(new_n1027), .ZN(G1355gat));
endmodule


