//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n569, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n606, new_n608, new_n609, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  OR2_X1    g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n467), .A2(new_n464), .A3(G101), .A4(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n463), .A2(G137), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n470), .B1(new_n461), .B2(new_n462), .ZN(new_n471));
  AND2_X1   g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n463), .A2(G136), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT69), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n464), .B1(new_n461), .B2(new_n462), .ZN(new_n481));
  AOI211_X1 g056(.A(new_n478), .B(new_n480), .C1(G124), .C2(new_n481), .ZN(G162));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI211_X1 g059(.A(G126), .B(G2105), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(new_n488), .A3(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n483), .B2(new_n484), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n492), .B(new_n495), .C1(new_n484), .C2(new_n483), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n490), .B1(new_n494), .B2(new_n496), .ZN(G164));
  AND2_X1   g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  NOR2_X1   g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G50), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n503), .B(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n507));
  XNOR2_X1  g082(.A(new_n506), .B(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n510), .A2(new_n500), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n504), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n508), .A2(new_n509), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n513), .A2(new_n518), .ZN(G166));
  OR2_X1    g094(.A1(new_n498), .A2(new_n499), .ZN(new_n520));
  XOR2_X1   g095(.A(KEYINPUT73), .B(G89), .Z(new_n521));
  NAND3_X1  g096(.A1(new_n515), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n502), .A2(G51), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n522), .A2(new_n523), .A3(new_n526), .A4(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  AOI22_X1  g104(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n514), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n502), .A2(G52), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n515), .A2(new_n520), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n531), .A2(new_n535), .ZN(G171));
  NAND4_X1  g111(.A1(new_n508), .A2(G81), .A3(new_n509), .A4(new_n520), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n520), .A2(G543), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n510), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G651), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n540), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n543), .A2(KEYINPUT74), .A3(G651), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI211_X1 g132(.A(new_n555), .B(new_n556), .C1(new_n539), .C2(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n508), .A2(G91), .A3(new_n509), .A4(new_n520), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n557), .B1(KEYINPUT75), .B2(KEYINPUT9), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n502), .B(new_n560), .C1(KEYINPUT75), .C2(KEYINPUT9), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n508), .A2(G65), .A3(new_n509), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n514), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  AOI22_X1  g143(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n504), .B(new_n512), .C1(new_n569), .C2(new_n514), .ZN(G303));
  NAND4_X1  g145(.A1(new_n508), .A2(G87), .A3(new_n509), .A4(new_n520), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n502), .A2(G49), .ZN(new_n572));
  AOI21_X1  g147(.A(G74), .B1(new_n508), .B2(new_n509), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n514), .ZN(G288));
  NAND3_X1  g149(.A1(new_n508), .A2(G61), .A3(new_n509), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n508), .A2(G86), .A3(new_n509), .A4(new_n520), .ZN(new_n579));
  OAI211_X1 g154(.A(G48), .B(G543), .C1(new_n498), .C2(new_n499), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT76), .Z(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(new_n502), .A2(G47), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n533), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n515), .A2(G60), .ZN(new_n586));
  NAND2_X1  g161(.A1(G72), .A2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n514), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n585), .A2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  XOR2_X1   g165(.A(KEYINPUT77), .B(KEYINPUT10), .Z(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n533), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n511), .A2(G92), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n502), .A2(G54), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n514), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n590), .B1(G868), .B2(new_n600), .ZN(G284));
  XNOR2_X1  g176(.A(G284), .B(KEYINPUT78), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n566), .ZN(G297));
  OAI21_X1  g179(.A(new_n603), .B1(G868), .B2(new_n566), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n600), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n600), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g185(.A(KEYINPUT79), .B(KEYINPUT11), .ZN(new_n611));
  XNOR2_X1  g186(.A(G323), .B(new_n611), .ZN(G282));
  XNOR2_X1  g187(.A(KEYINPUT3), .B(G2104), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n464), .A2(G2104), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  XOR2_X1   g193(.A(KEYINPUT80), .B(G2100), .Z(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n463), .A2(G135), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n481), .A2(G123), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n464), .A2(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  NAND3_X1  g202(.A1(new_n620), .A2(new_n621), .A3(new_n627), .ZN(G156));
  XOR2_X1   g203(.A(KEYINPUT15), .B(G2435), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2438), .ZN(new_n630));
  XOR2_X1   g205(.A(G2427), .B(G2430), .Z(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT82), .B(KEYINPUT14), .Z(new_n633));
  NAND2_X1  g208(.A1(new_n630), .A2(new_n631), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n635), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(G14), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT83), .Z(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT84), .Z(G401));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT85), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT17), .Z(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT87), .ZN(new_n655));
  INV_X1    g230(.A(new_n651), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n649), .B2(new_n652), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n657), .A2(KEYINPUT86), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(KEYINPUT86), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n658), .B(new_n659), .C1(new_n650), .C2(new_n653), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT18), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n655), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2096), .B(G2100), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT20), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n667), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n667), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1991), .B(G1996), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(G229));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G23), .ZN(new_n686));
  INV_X1    g261(.A(G288), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n685), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT33), .B(G1976), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n688), .B(new_n689), .Z(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(KEYINPUT91), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(KEYINPUT91), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n685), .A2(G22), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G166), .B2(new_n685), .ZN(new_n694));
  INV_X1    g269(.A(G1971), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(G6), .A2(G16), .ZN(new_n697));
  INV_X1    g272(.A(G305), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(G16), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND4_X1  g276(.A1(new_n691), .A2(new_n692), .A3(new_n696), .A4(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(KEYINPUT34), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(KEYINPUT34), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n685), .A2(G24), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n585), .A2(new_n588), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n685), .ZN(new_n707));
  INV_X1    g282(.A(G1986), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G25), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n463), .A2(G131), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT88), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n717));
  INV_X1    g292(.A(G107), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(G2105), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G119), .B2(new_n481), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n714), .B1(new_n722), .B2(new_n713), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT89), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n723), .B(new_n725), .ZN(new_n726));
  NOR3_X1   g301(.A1(new_n711), .A2(new_n712), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n703), .A2(new_n704), .A3(new_n727), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT36), .Z(new_n729));
  INV_X1    g304(.A(G34), .ZN(new_n730));
  AOI21_X1  g305(.A(G29), .B1(new_n730), .B2(KEYINPUT24), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(KEYINPUT24), .B2(new_n730), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n474), .B2(new_n713), .ZN(new_n733));
  INV_X1    g308(.A(G2084), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT31), .B(G11), .Z(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT30), .B(G28), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n736), .B1(new_n713), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT25), .Z(new_n740));
  INV_X1    g315(.A(G139), .ZN(new_n741));
  INV_X1    g316(.A(new_n463), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n613), .A2(G127), .ZN(new_n744));
  NAND2_X1  g319(.A1(G115), .A2(G2104), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n464), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G29), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G29), .B2(G33), .ZN(new_n749));
  INV_X1    g324(.A(G2072), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n738), .B1(new_n713), .B2(new_n626), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n735), .B(new_n751), .C1(new_n750), .C2(new_n749), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n713), .A2(G26), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT28), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n463), .A2(G140), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n481), .A2(G128), .ZN(new_n756));
  OR2_X1    g331(.A1(G104), .A2(G2105), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n757), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n754), .B1(new_n760), .B2(new_n713), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2067), .ZN(new_n762));
  NOR2_X1   g337(.A1(G168), .A2(new_n685), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n685), .B2(G21), .ZN(new_n764));
  INV_X1    g339(.A(G1966), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G171), .A2(new_n685), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G5), .B2(new_n685), .ZN(new_n768));
  INV_X1    g343(.A(G1961), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n733), .A2(new_n734), .ZN(new_n771));
  NAND2_X1  g346(.A1(G164), .A2(G29), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G27), .B2(G29), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT95), .B(G2078), .Z(new_n774));
  OAI21_X1  g349(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n773), .B2(new_n774), .ZN(new_n776));
  AND4_X1   g351(.A1(new_n752), .A2(new_n766), .A3(new_n770), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G29), .A2(G32), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n615), .A2(G105), .ZN(new_n779));
  INV_X1    g354(.A(G141), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n742), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g356(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT26), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n481), .A2(G129), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT93), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n778), .B1(new_n787), .B2(G29), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT27), .B(G1996), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OAI22_X1  g365(.A1(new_n768), .A2(new_n769), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n790), .B2(new_n788), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n764), .A2(new_n765), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT94), .ZN(new_n794));
  NOR2_X1   g369(.A1(G4), .A2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n600), .B2(G16), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT92), .B(G1348), .Z(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n777), .A2(new_n792), .A3(new_n794), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n713), .A2(G35), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G162), .B2(new_n713), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2090), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n685), .A2(G19), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n549), .B2(new_n685), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(G1341), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n685), .A2(G20), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT23), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n566), .B2(new_n685), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1956), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n796), .B2(new_n797), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n804), .A2(new_n807), .A3(new_n812), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n729), .A2(new_n799), .A3(new_n813), .ZN(G311));
  INV_X1    g389(.A(G311), .ZN(G150));
  NAND3_X1  g390(.A1(new_n508), .A2(G67), .A3(new_n509), .ZN(new_n816));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n514), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n508), .A2(G93), .A3(new_n509), .A4(new_n520), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT98), .B(G55), .Z(new_n820));
  NAND2_X1  g395(.A1(new_n502), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(G860), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT37), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(KEYINPUT99), .B1(new_n818), .B2(new_n822), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n548), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n546), .A2(new_n828), .A3(new_n547), .A4(new_n829), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n600), .A2(G559), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n836));
  XOR2_X1   g411(.A(new_n835), .B(new_n836), .Z(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n824), .B1(new_n838), .B2(KEYINPUT39), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n826), .B1(new_n839), .B2(new_n840), .ZN(G145));
  XNOR2_X1  g416(.A(new_n721), .B(new_n617), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n463), .A2(G142), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n481), .A2(G130), .ZN(new_n844));
  OR2_X1    g419(.A1(G106), .A2(G2105), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n845), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n842), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n494), .A2(new_n496), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n485), .A2(new_n489), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n760), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(G164), .A2(new_n759), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(KEYINPUT100), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n853), .B2(new_n854), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n856), .A2(new_n787), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n787), .B1(new_n856), .B2(new_n858), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n747), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n855), .A2(new_n786), .ZN(new_n862));
  INV_X1    g437(.A(new_n786), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n853), .B2(new_n854), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n862), .B(new_n864), .C1(new_n746), .C2(new_n743), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n849), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n626), .B(new_n474), .ZN(new_n867));
  XNOR2_X1  g442(.A(G162), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n861), .A2(new_n849), .A3(new_n865), .ZN(new_n871));
  AOI21_X1  g446(.A(G37), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n866), .B2(KEYINPUT101), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n861), .A2(new_n849), .A3(new_n874), .A4(new_n865), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT102), .B1(new_n876), .B2(new_n869), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  AOI211_X1 g453(.A(new_n878), .B(new_n868), .C1(new_n873), .C2(new_n875), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n872), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g456(.A(G868), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n818), .B2(new_n822), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n596), .A2(new_n599), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G299), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n600), .A2(new_n566), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(KEYINPUT41), .A3(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n608), .B(KEYINPUT103), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n833), .ZN(new_n893));
  MUX2_X1   g468(.A(new_n891), .B(new_n887), .S(new_n893), .Z(new_n894));
  NAND2_X1  g469(.A1(G290), .A2(G288), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n706), .A2(new_n687), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT104), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n706), .A2(new_n687), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n585), .A2(new_n588), .A3(G288), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n698), .B(G303), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n897), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(G303), .B(G305), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n904), .A2(KEYINPUT104), .A3(new_n895), .A4(new_n896), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT42), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n903), .A2(KEYINPUT105), .A3(new_n905), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT105), .B1(new_n903), .B2(new_n905), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n906), .B1(new_n909), .B2(KEYINPUT42), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n894), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n883), .B1(new_n911), .B2(new_n882), .ZN(G295));
  OAI21_X1  g487(.A(new_n883), .B1(new_n911), .B2(new_n882), .ZN(G331));
  AND3_X1   g488(.A1(new_n831), .A2(G301), .A3(new_n832), .ZN(new_n914));
  AOI21_X1  g489(.A(G301), .B1(new_n831), .B2(new_n832), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n914), .A2(new_n915), .A3(G286), .ZN(new_n916));
  INV_X1    g491(.A(new_n832), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n547), .A2(new_n546), .B1(new_n828), .B2(new_n829), .ZN(new_n918));
  OAI21_X1  g493(.A(G171), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n831), .A2(G301), .A3(new_n832), .ZN(new_n920));
  AOI21_X1  g495(.A(G168), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n891), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(G286), .B1(new_n914), .B2(new_n915), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(G168), .A3(new_n920), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n887), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(KEYINPUT106), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n909), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n907), .A2(new_n908), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n929), .A2(new_n922), .A3(KEYINPUT106), .A4(new_n925), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n927), .A2(new_n933), .A3(new_n928), .A4(new_n930), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n935), .B(new_n938), .Z(G397));
  NAND3_X1  g514(.A1(new_n469), .A2(new_n473), .A3(G40), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n469), .A2(new_n473), .A3(KEYINPUT109), .A4(G40), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G1384), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n852), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n949), .A2(G1996), .A3(new_n863), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n950), .B(KEYINPUT110), .Z(new_n951));
  INV_X1    g526(.A(G1996), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n787), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n759), .B(G2067), .Z(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n949), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n951), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT111), .ZN(new_n958));
  INV_X1    g533(.A(new_n949), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n721), .B(new_n724), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n960), .B2(KEYINPUT112), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(KEYINPUT112), .B2(new_n960), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n706), .B(G1986), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n964), .B1(new_n959), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT124), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT122), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n969));
  NAND2_X1  g544(.A1(G286), .A2(G8), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT121), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n974));
  INV_X1    g549(.A(new_n496), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n495), .B1(new_n613), .B2(new_n492), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n974), .B(new_n945), .C1(new_n977), .C2(new_n490), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n973), .A2(KEYINPUT113), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n946), .A2(new_n980), .A3(KEYINPUT50), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT115), .B(G2084), .Z(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n942), .A2(new_n943), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(G164), .B2(G1384), .ZN(new_n989));
  INV_X1    g564(.A(new_n947), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n852), .A2(new_n945), .A3(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n989), .A2(new_n991), .A3(new_n942), .A4(new_n943), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n765), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n987), .A2(new_n993), .ZN(new_n994));
  OAI211_X1 g569(.A(G8), .B(new_n972), .C1(new_n994), .C2(G286), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT45), .B1(new_n852), .B2(new_n945), .ZN(new_n996));
  AOI211_X1 g571(.A(G1384), .B(new_n947), .C1(new_n850), .C2(new_n851), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n942), .A2(new_n943), .ZN(new_n999));
  AOI21_X1  g574(.A(G1966), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n985), .B1(new_n979), .B2(new_n981), .ZN(new_n1001));
  OAI21_X1  g576(.A(G8), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n970), .A2(new_n971), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT51), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n970), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n995), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n970), .B1(new_n987), .B2(new_n993), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n968), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  AOI211_X1 g584(.A(KEYINPUT122), .B(new_n1007), .C1(new_n995), .C2(new_n1005), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1009), .A2(new_n1010), .A3(KEYINPUT62), .ZN(new_n1011));
  OAI21_X1  g586(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1012), .A2(G1976), .A3(new_n571), .A4(new_n572), .ZN(new_n1013));
  NOR2_X1   g588(.A1(G164), .A2(G1384), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(new_n942), .A3(new_n943), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(new_n1015), .A3(G8), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT52), .ZN(new_n1017));
  INV_X1    g592(.A(G1976), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT52), .B1(G288), .B2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1019), .A2(new_n1013), .A3(new_n1015), .A4(G8), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n581), .A2(new_n579), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n514), .B1(new_n575), .B2(new_n576), .ZN(new_n1023));
  OAI21_X1  g598(.A(G1981), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1981), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n578), .A2(new_n1025), .A3(new_n579), .A4(new_n581), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1024), .A2(new_n1026), .A3(KEYINPUT49), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1024), .A2(new_n1026), .A3(KEYINPUT114), .A4(KEYINPUT49), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT49), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1015), .A2(G8), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1021), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n944), .B1(new_n979), .B2(new_n981), .ZN(new_n1036));
  INV_X1    g611(.A(G2090), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1014), .A2(KEYINPUT45), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n999), .A2(new_n948), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n695), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n1043));
  INV_X1    g618(.A(G8), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(G166), .B2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(KEYINPUT55), .B(G8), .C1(new_n513), .C2(new_n518), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1042), .A2(new_n1047), .A3(G8), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1046), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n973), .A2(new_n978), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1052), .A2(new_n944), .A3(G2090), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(new_n695), .B2(new_n1040), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1051), .B1(new_n1054), .B2(new_n1044), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1035), .A2(new_n1048), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n1040), .B2(G2078), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n982), .B2(new_n999), .ZN(new_n1061));
  AOI211_X1 g636(.A(KEYINPUT117), .B(new_n944), .C1(new_n979), .C2(new_n981), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1059), .B1(new_n1063), .B2(new_n769), .ZN(new_n1064));
  OR3_X1    g639(.A1(new_n992), .A2(KEYINPUT123), .A3(G2078), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT123), .B1(new_n992), .B2(G2078), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(KEYINPUT53), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(G301), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1056), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n967), .B1(new_n1011), .B2(new_n1069), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1002), .A2(new_n970), .A3(new_n1004), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1004), .B1(new_n1002), .B2(new_n970), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1008), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT122), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT62), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1006), .A2(new_n968), .A3(new_n1008), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1056), .A2(new_n1068), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(KEYINPUT124), .A3(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT62), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT125), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1082), .B(KEYINPUT62), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1070), .A2(new_n1079), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n687), .A2(new_n1018), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1026), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1033), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1048), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1087), .A2(new_n1088), .B1(new_n1089), .B2(new_n1035), .ZN(new_n1090));
  OAI211_X1 g665(.A(G8), .B(G168), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1035), .A2(new_n1048), .A3(new_n1055), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT63), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1042), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1051), .B1(new_n1096), .B2(new_n1044), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n1048), .A2(new_n1097), .A3(new_n1035), .A4(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1090), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1101), .A2(KEYINPUT57), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(KEYINPUT57), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n566), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1101), .B(KEYINPUT57), .C1(new_n562), .C2(new_n565), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G1956), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n1052), .B2(new_n944), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n999), .A2(new_n948), .A3(new_n1039), .A4(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1112), .A2(KEYINPUT118), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1110), .A2(new_n1108), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(KEYINPUT118), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1113), .A2(KEYINPUT119), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G1348), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1063), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1015), .A2(G2067), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n884), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1111), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1122), .A2(KEYINPUT60), .A3(new_n1124), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT60), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1127), .A2(new_n1128), .A3(new_n884), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1111), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1106), .A2(KEYINPUT61), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1131), .A2(new_n1132), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1122), .A2(KEYINPUT60), .A3(new_n884), .A4(new_n1124), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT58), .B(G1341), .Z(new_n1136));
  NAND2_X1  g711(.A1(new_n1015), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1040), .B2(G1996), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT120), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1140), .B(new_n1137), .C1(new_n1040), .C2(G1996), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1135), .B1(new_n1142), .B2(new_n549), .ZN(new_n1143));
  AOI211_X1 g718(.A(KEYINPUT59), .B(new_n548), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1133), .B(new_n1134), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1126), .B1(new_n1129), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1147));
  XOR2_X1   g722(.A(G171), .B(KEYINPUT54), .Z(new_n1148));
  NOR3_X1   g723(.A1(new_n940), .A2(new_n1057), .A3(G2078), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1039), .A2(new_n948), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1148), .B1(new_n1064), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1061), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1062), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(new_n1153), .A3(new_n769), .ZN(new_n1154));
  AND4_X1   g729(.A1(new_n1154), .A2(new_n1148), .A3(new_n1058), .A4(new_n1067), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1056), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1147), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1100), .B1(new_n1146), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n966), .B1(new_n1084), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n706), .A2(new_n949), .A3(new_n708), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT48), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n964), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT111), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n957), .B(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n722), .A2(new_n724), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n759), .A2(G2067), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n949), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n949), .B1(new_n955), .B2(new_n863), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n959), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT46), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1171), .B1(new_n949), .B2(new_n952), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1169), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT47), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1162), .A2(new_n1168), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(KEYINPUT126), .B1(new_n1159), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1079), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1177));
  AOI21_X1  g752(.A(KEYINPUT124), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1158), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n966), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1162), .A2(new_n1168), .A3(new_n1174), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1176), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g760(.A1(G227), .A2(new_n459), .ZN(new_n1187));
  OAI211_X1 g761(.A(new_n1187), .B(new_n646), .C1(new_n682), .C2(new_n683), .ZN(new_n1188));
  INV_X1    g762(.A(new_n1188), .ZN(new_n1189));
  AND2_X1   g763(.A1(new_n880), .A2(new_n1189), .ZN(new_n1190));
  AND3_X1   g764(.A1(new_n1190), .A2(new_n935), .A3(KEYINPUT127), .ZN(new_n1191));
  AOI21_X1  g765(.A(KEYINPUT127), .B1(new_n1190), .B2(new_n935), .ZN(new_n1192));
  NOR2_X1   g766(.A1(new_n1191), .A2(new_n1192), .ZN(G308));
  NAND2_X1  g767(.A1(new_n1190), .A2(new_n935), .ZN(G225));
endmodule


