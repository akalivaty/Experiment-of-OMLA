//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT64), .B(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G58), .A2(G232), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n206), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  AND2_X1   g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G20), .ZN(new_n220));
  OAI21_X1  g0020(.A(G50), .B1(G58), .B2(G68), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n209), .B1(KEYINPUT1), .B2(new_n218), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XNOR2_X1  g0023(.A(G238), .B(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT2), .B(G226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(G264), .B(G270), .Z(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n228), .B(new_n231), .Z(G358));
  XOR2_X1   g0032(.A(G58), .B(G77), .Z(new_n233));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G351));
  XNOR2_X1  g0039(.A(KEYINPUT3), .B(G33), .ZN(new_n240));
  INV_X1    g0040(.A(G1698), .ZN(new_n241));
  NAND3_X1  g0041(.A1(new_n240), .A2(G222), .A3(new_n241), .ZN(new_n242));
  NAND3_X1  g0042(.A1(new_n240), .A2(G223), .A3(G1698), .ZN(new_n243));
  OAI211_X1 g0043(.A(new_n242), .B(new_n243), .C1(new_n210), .C2(new_n240), .ZN(new_n244));
  NAND2_X1  g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n245), .A2(G1), .A3(G13), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  INV_X1    g0049(.A(G41), .ZN(new_n250));
  INV_X1    g0050(.A(G45), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI22_X1  g0052(.A1(new_n249), .A2(new_n252), .B1(new_n219), .B2(new_n245), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n254), .B1(new_n219), .B2(new_n245), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1), .B1(new_n250), .B2(new_n251), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n253), .A2(G226), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n248), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G169), .ZN(new_n259));
  INV_X1    g0059(.A(G179), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(new_n258), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT8), .B(G58), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT66), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G58), .ZN(new_n267));
  OR3_X1    g0067(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT8), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G20), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n263), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G1), .A2(G13), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(new_n206), .B2(new_n270), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT65), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n275), .B(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n275), .B(KEYINPUT65), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n249), .A2(G13), .A3(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT67), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT67), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n282), .A2(new_n249), .A3(G13), .A4(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n249), .A2(G20), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n279), .A2(G50), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT68), .ZN(new_n287));
  INV_X1    g0087(.A(new_n284), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n202), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n287), .B1(new_n286), .B2(new_n289), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n278), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n261), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n248), .A2(G190), .A3(new_n257), .ZN(new_n294));
  INV_X1    g0094(.A(G200), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n294), .B1(new_n258), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT9), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n296), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(KEYINPUT9), .B(new_n278), .C1(new_n290), .C2(new_n291), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT71), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n299), .A2(new_n300), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n305), .B(new_n298), .C1(new_n301), .C2(new_n302), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n293), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n269), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n285), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n279), .A2(new_n284), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n309), .A2(new_n310), .B1(new_n308), .B2(new_n284), .ZN(new_n311));
  INV_X1    g0111(.A(new_n275), .ZN(new_n312));
  AND2_X1   g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  NOR2_X1   g0113(.A1(KEYINPUT3), .A2(G33), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G20), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT7), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT7), .ZN(new_n318));
  NOR4_X1   g0118(.A1(new_n313), .A2(new_n314), .A3(new_n318), .A4(G20), .ZN(new_n319));
  OAI21_X1  g0119(.A(G68), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G68), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n267), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(G20), .B1(new_n322), .B2(new_n201), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n262), .A2(G159), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT16), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n312), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n320), .A2(KEYINPUT16), .A3(new_n326), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n311), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OR2_X1    g0131(.A1(G223), .A2(G1698), .ZN(new_n332));
  INV_X1    g0132(.A(G226), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G1698), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n332), .B(new_n334), .C1(new_n313), .C2(new_n314), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G87), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n247), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n253), .A2(G232), .B1(new_n255), .B2(new_n256), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(KEYINPUT76), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT76), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n246), .B1(new_n335), .B2(new_n336), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n256), .A2(new_n246), .A3(G274), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n246), .A2(G232), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n341), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n340), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n295), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n342), .A2(new_n346), .ZN(new_n350));
  INV_X1    g0150(.A(G190), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT77), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT17), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n331), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n318), .B1(new_n240), .B2(G20), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n315), .A2(KEYINPUT7), .A3(new_n316), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n321), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n328), .B1(new_n359), .B2(new_n325), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(new_n330), .A3(new_n275), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n269), .B1(new_n249), .B2(G20), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n277), .A2(new_n288), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n362), .A2(new_n363), .B1(new_n269), .B2(new_n288), .ZN(new_n364));
  AOI21_X1  g0164(.A(G200), .B1(new_n340), .B2(new_n347), .ZN(new_n365));
  INV_X1    g0165(.A(new_n352), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n361), .B(new_n364), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  XOR2_X1   g0167(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n356), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G107), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n246), .B1(new_n315), .B2(new_n371), .ZN(new_n372));
  MUX2_X1   g0172(.A(G232), .B(G238), .S(G1698), .Z(new_n373));
  OAI21_X1  g0173(.A(new_n372), .B1(new_n315), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n253), .A2(G244), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n343), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G200), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n351), .B2(new_n376), .ZN(new_n378));
  INV_X1    g0178(.A(new_n210), .ZN(new_n379));
  XOR2_X1   g0179(.A(KEYINPUT15), .B(G87), .Z(new_n380));
  AOI22_X1  g0180(.A1(new_n379), .A2(G20), .B1(new_n380), .B2(new_n271), .ZN(new_n381));
  INV_X1    g0181(.A(new_n262), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n382), .A2(KEYINPUT69), .ZN(new_n383));
  INV_X1    g0183(.A(new_n264), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT69), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n384), .B1(new_n385), .B2(new_n262), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n381), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(new_n275), .B1(new_n210), .B2(new_n288), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n275), .B1(new_n281), .B2(new_n283), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(G77), .A3(new_n285), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n378), .B1(KEYINPUT70), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT70), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(new_n393), .A3(new_n390), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n361), .A2(new_n364), .ZN(new_n396));
  INV_X1    g0196(.A(G169), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n348), .A2(new_n397), .B1(new_n260), .B2(new_n350), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT18), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT18), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n396), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n376), .A2(G179), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n376), .A2(new_n397), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n391), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NOR4_X1   g0207(.A1(new_n370), .A2(new_n395), .A3(new_n403), .A4(new_n407), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n271), .A2(G77), .B1(G20), .B2(new_n321), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n202), .B2(new_n382), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n277), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT12), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n288), .A2(new_n413), .A3(new_n321), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT12), .B1(new_n284), .B2(G68), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n412), .A2(KEYINPUT11), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT74), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT11), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n321), .B1(new_n249), .B2(G20), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n411), .A2(new_n418), .B1(new_n389), .B2(new_n419), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n416), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n417), .B1(new_n416), .B2(new_n420), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n333), .A2(new_n241), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n225), .A2(G1698), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n424), .B(new_n425), .C1(new_n313), .C2(new_n314), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G97), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n247), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT13), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n253), .A2(G238), .B1(new_n255), .B2(new_n256), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n246), .B1(new_n426), .B2(new_n427), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n246), .A2(G238), .A3(new_n344), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n343), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT13), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n432), .A2(KEYINPUT72), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT72), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n429), .A2(new_n431), .A3(new_n438), .A4(new_n430), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(G169), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT14), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT14), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n437), .A2(new_n442), .A3(G169), .A4(new_n439), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n432), .A2(G179), .A3(new_n436), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT73), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT73), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n432), .A2(new_n436), .A3(new_n446), .A4(G179), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n441), .A2(new_n443), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n423), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n437), .A2(G200), .A3(new_n439), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n432), .A2(G190), .A3(new_n436), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n451), .A2(new_n420), .A3(new_n416), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n454), .A2(KEYINPUT75), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(KEYINPUT75), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n307), .A2(new_n408), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT6), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT78), .ZN(new_n459));
  INV_X1    g0259(.A(G97), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(new_n371), .ZN(new_n461));
  NOR2_X1   g0261(.A1(G97), .A2(G107), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g0263(.A(G97), .B(G107), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT78), .ZN(new_n465));
  MUX2_X1   g0265(.A(new_n465), .B(G97), .S(KEYINPUT6), .Z(new_n466));
  OAI211_X1 g0266(.A(new_n463), .B(G20), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n262), .A2(G77), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n371), .B1(new_n357), .B2(new_n358), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n275), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n249), .A2(G33), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n363), .A2(G97), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n288), .A2(new_n460), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(G244), .B(new_n241), .C1(new_n313), .C2(new_n314), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT4), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n240), .A2(KEYINPUT4), .A3(G244), .A4(new_n241), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n240), .A2(G250), .A3(G1698), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n478), .A2(new_n479), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n247), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n251), .A2(G1), .ZN(new_n484));
  AND2_X1   g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  NOR2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(G257), .A3(new_n246), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT5), .B(G41), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n255), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n483), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(KEYINPUT79), .A3(G200), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT79), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n491), .B1(new_n482), .B2(new_n247), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(new_n295), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(G190), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n475), .A2(new_n494), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n493), .A2(new_n397), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n496), .A2(new_n260), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n281), .A2(new_n371), .A3(new_n283), .ZN(new_n505));
  XOR2_X1   g0305(.A(new_n505), .B(KEYINPUT25), .Z(new_n506));
  NAND4_X1  g0306(.A1(new_n279), .A2(G107), .A3(new_n284), .A4(new_n472), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n316), .B(G87), .C1(new_n313), .C2(new_n314), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT22), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT22), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n240), .A2(new_n511), .A3(new_n316), .A4(G87), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(KEYINPUT86), .B(KEYINPUT23), .C1(new_n316), .C2(G107), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n316), .A2(G33), .A3(G116), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n371), .A2(G20), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n514), .B(new_n515), .C1(KEYINPUT23), .C2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT86), .B1(new_n516), .B2(KEYINPUT23), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT24), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n513), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(new_n513), .B2(new_n519), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n275), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n508), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(G257), .B(G1698), .C1(new_n313), .C2(new_n314), .ZN(new_n525));
  OAI211_X1 g0325(.A(G250), .B(new_n241), .C1(new_n313), .C2(new_n314), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G294), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n247), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n487), .A2(G264), .A3(new_n246), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n490), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G169), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n489), .A2(new_n484), .B1(new_n219), .B2(new_n245), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT87), .B1(new_n533), .B2(G264), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n487), .A2(KEYINPUT87), .A3(G264), .A4(new_n246), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n529), .B(new_n490), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n532), .B1(new_n260), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n524), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT87), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n530), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(new_n535), .B1(new_n247), .B2(new_n528), .ZN(new_n542));
  AOI21_X1  g0342(.A(G200), .B1(new_n542), .B2(new_n490), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n531), .A2(G190), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n508), .B(new_n523), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n249), .A2(G45), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n546), .A2(G250), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n246), .A2(new_n547), .B1(new_n255), .B2(new_n484), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(G244), .B(G1698), .C1(new_n313), .C2(new_n314), .ZN(new_n550));
  OAI211_X1 g0350(.A(G238), .B(new_n241), .C1(new_n313), .C2(new_n314), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G116), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT80), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n246), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT80), .A4(new_n552), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n549), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G190), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n240), .A2(new_n316), .A3(G68), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n272), .A2(new_n460), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n560), .B2(KEYINPUT19), .ZN(new_n561));
  NAND3_X1  g0361(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT81), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n562), .A2(new_n563), .A3(new_n316), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n563), .B1(new_n562), .B2(new_n316), .ZN(new_n565));
  NOR3_X1   g0365(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n566));
  NOR3_X1   g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n275), .B1(new_n561), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n279), .A2(G87), .A3(new_n284), .A4(new_n472), .ZN(new_n569));
  INV_X1    g0369(.A(new_n380), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n288), .A2(new_n570), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n558), .B(new_n572), .C1(new_n295), .C2(new_n557), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n557), .A2(new_n260), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n279), .A2(new_n284), .A3(new_n380), .A4(new_n472), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n568), .A2(new_n575), .A3(new_n571), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n574), .B(new_n576), .C1(G169), .C2(new_n557), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n545), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n504), .A2(new_n539), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n490), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n487), .A2(G270), .A3(new_n246), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT82), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n487), .A2(KEYINPUT82), .A3(G270), .A4(new_n246), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n580), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(G257), .B(new_n241), .C1(new_n313), .C2(new_n314), .ZN(new_n586));
  OAI211_X1 g0386(.A(G264), .B(G1698), .C1(new_n313), .C2(new_n314), .ZN(new_n587));
  INV_X1    g0387(.A(G303), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n240), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT83), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n589), .A2(new_n590), .A3(new_n247), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n590), .B1(new_n589), .B2(new_n247), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n585), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G116), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n281), .A2(new_n594), .A3(new_n283), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n595), .B(KEYINPUT84), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n480), .B(new_n316), .C1(G33), .C2(new_n460), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(G20), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n275), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT20), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n597), .A2(new_n275), .A3(KEYINPUT20), .A4(new_n598), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n594), .B1(new_n249), .B2(G33), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n601), .A2(new_n602), .B1(new_n389), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n397), .B1(new_n596), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n593), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT21), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT85), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n585), .B(G179), .C1(new_n591), .C2(new_n592), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n596), .A2(new_n604), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n608), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT85), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n593), .A2(new_n605), .A3(new_n615), .A4(KEYINPUT21), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n593), .A2(G200), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n589), .A2(new_n247), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT83), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n589), .A2(new_n590), .A3(new_n247), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n621), .A2(G190), .A3(new_n585), .ZN(new_n622));
  INV_X1    g0422(.A(new_n612), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n617), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n614), .A2(new_n616), .A3(new_n624), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n457), .A2(new_n579), .A3(new_n625), .ZN(G372));
  INV_X1    g0426(.A(new_n457), .ZN(new_n627));
  INV_X1    g0427(.A(new_n577), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n499), .A2(new_n503), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n545), .A2(new_n573), .A3(new_n577), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n612), .A2(new_n611), .B1(new_n606), .B2(new_n607), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(new_n539), .A3(new_n616), .A4(new_n608), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n628), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n573), .A2(new_n577), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n503), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(KEYINPUT26), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n635), .B2(new_n503), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n627), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n304), .A2(new_n306), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n396), .A2(new_n398), .A3(new_n401), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n401), .B1(new_n396), .B2(new_n398), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n423), .A2(new_n449), .B1(new_n407), .B2(new_n453), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(new_n370), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n293), .B1(new_n644), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n643), .A2(new_n650), .ZN(G369));
  NAND4_X1  g0451(.A1(new_n608), .A2(new_n609), .A3(new_n616), .A4(new_n613), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n249), .A2(new_n316), .A3(G13), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  OAI21_X1  g0454(.A(G213), .B1(new_n653), .B2(KEYINPUT27), .ZN(new_n655));
  OR3_X1    g0455(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT88), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT88), .B1(new_n654), .B2(new_n655), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(new_n623), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n652), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n625), .B2(new_n662), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n539), .A2(new_n661), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT89), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n524), .A2(new_n660), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n669), .A2(new_n539), .A3(new_n545), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n652), .A2(new_n661), .ZN(new_n673));
  INV_X1    g0473(.A(new_n539), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n671), .A2(new_n673), .B1(new_n674), .B2(new_n661), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n675), .ZN(G399));
  NAND2_X1  g0476(.A1(new_n566), .A2(new_n594), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n207), .A2(new_n250), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G1), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n221), .B2(new_n679), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n642), .A2(new_n661), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(KEYINPUT29), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT29), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n642), .B2(new_n661), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G330), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n614), .A2(new_n616), .A3(new_n624), .A4(new_n661), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n579), .ZN(new_n690));
  XOR2_X1   g0490(.A(KEYINPUT90), .B(KEYINPUT31), .Z(new_n691));
  NAND2_X1  g0491(.A1(new_n553), .A2(new_n554), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(new_n247), .A3(new_n556), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n548), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n593), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n493), .A2(new_n260), .A3(new_n537), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n496), .A2(new_n542), .A3(new_n693), .A4(new_n548), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(new_n610), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n697), .B1(KEYINPUT30), .B2(new_n699), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n557), .A2(new_n542), .A3(new_n496), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(new_n611), .A3(KEYINPUT91), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT91), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n698), .B2(new_n610), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  AOI211_X1 g0506(.A(new_n661), .B(new_n691), .C1(new_n700), .C2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n690), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n557), .B1(new_n621), .B2(new_n585), .ZN(new_n709));
  AOI21_X1  g0509(.A(G179), .B1(new_n542), .B2(new_n490), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n709), .A2(KEYINPUT92), .A3(new_n710), .A4(new_n493), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT92), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n695), .B2(new_n696), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n701), .A2(new_n611), .A3(KEYINPUT30), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n661), .B1(new_n716), .B2(new_n706), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(KEYINPUT31), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n688), .B1(new_n708), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n687), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n682), .B1(new_n723), .B2(G1), .ZN(G364));
  OR2_X1    g0524(.A1(new_n664), .A2(G330), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n316), .A2(G13), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n249), .B1(new_n726), .B2(G45), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n679), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n725), .A2(new_n665), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n728), .B(KEYINPUT93), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n240), .A2(new_n207), .ZN(new_n731));
  INV_X1    g0531(.A(G355), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n731), .A2(new_n732), .B1(G116), .B2(new_n207), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n235), .A2(new_n251), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n315), .A2(new_n207), .ZN(new_n735));
  INV_X1    g0535(.A(new_n221), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(new_n251), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n733), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n274), .B1(G20), .B2(new_n397), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n730), .B1(new_n738), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n316), .A2(G190), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G179), .A2(G200), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n748), .A2(KEYINPUT94), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(KEYINPUT94), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G329), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n316), .A2(new_n351), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n260), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G322), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n746), .A2(new_n755), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n756), .A2(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n754), .A2(new_n260), .A3(G200), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n240), .B(new_n760), .C1(G303), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n316), .A2(new_n260), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(G190), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(G326), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n316), .B1(new_n747), .B2(G190), .ZN(new_n767));
  INV_X1    g0567(.A(G294), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n765), .A2(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n764), .A2(new_n351), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT33), .B(G317), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n746), .A2(new_n260), .A3(G200), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT95), .Z(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G283), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n753), .A2(new_n763), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n752), .A2(G159), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT32), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n767), .A2(new_n460), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n321), .B2(new_n770), .ZN(new_n782));
  INV_X1    g0582(.A(new_n765), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(G50), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n775), .A2(G107), .ZN(new_n785));
  INV_X1    g0585(.A(new_n756), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n315), .B1(new_n786), .B2(G58), .ZN(new_n787));
  INV_X1    g0587(.A(new_n758), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n762), .A2(G87), .B1(new_n788), .B2(new_n379), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n784), .A2(new_n785), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n777), .B1(new_n779), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n745), .B1(new_n791), .B2(new_n742), .ZN(new_n792));
  INV_X1    g0592(.A(new_n741), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n664), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n729), .A2(new_n794), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT96), .Z(G396));
  NOR2_X1   g0596(.A1(new_n406), .A2(new_n660), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n392), .A2(new_n394), .B1(new_n391), .B2(new_n660), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n799), .B2(new_n407), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n683), .B(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n802), .A2(new_n720), .B1(new_n679), .B2(new_n727), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(KEYINPUT98), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n802), .A2(new_n720), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n803), .B2(KEYINPUT98), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n800), .A2(new_n739), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n742), .A2(new_n739), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT97), .Z(new_n811));
  OAI21_X1  g0611(.A(new_n730), .B1(new_n811), .B2(G77), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G143), .A2(new_n786), .B1(new_n788), .B2(G159), .ZN(new_n813));
  INV_X1    g0613(.A(G137), .ZN(new_n814));
  INV_X1    g0614(.A(G150), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n813), .B1(new_n814), .B2(new_n765), .C1(new_n815), .C2(new_n770), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n775), .A2(G68), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n752), .A2(G132), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n240), .B1(new_n761), .B2(new_n202), .ZN(new_n821));
  INV_X1    g0621(.A(new_n767), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(G58), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n816), .A2(new_n817), .ZN(new_n825));
  INV_X1    g0625(.A(G283), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n781), .B1(new_n765), .B2(new_n588), .C1(new_n826), .C2(new_n770), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n761), .A2(new_n371), .B1(new_n756), .B2(new_n768), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n240), .B(new_n828), .C1(G116), .C2(new_n788), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n775), .A2(G87), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n829), .B(new_n830), .C1(new_n759), .C2(new_n751), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n824), .A2(new_n825), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n812), .B1(new_n832), .B2(new_n742), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n809), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n808), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G384));
  OAI21_X1  g0636(.A(new_n463), .B1(new_n464), .B2(new_n466), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT35), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n594), .B(new_n220), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT99), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n839), .A2(new_n840), .B1(new_n838), .B2(new_n837), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n840), .B2(new_n839), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT36), .ZN(new_n843));
  OR3_X1    g0643(.A1(new_n210), .A2(new_n221), .A3(new_n322), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n321), .A2(G50), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT100), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n249), .B(G13), .C1(new_n844), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n453), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n449), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n423), .A2(new_n660), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AND4_X1   g0653(.A1(KEYINPUT101), .A2(new_n450), .A3(new_n851), .A4(new_n453), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n849), .B1(new_n423), .B2(new_n449), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT101), .B1(new_n855), .B2(new_n851), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n853), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT103), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n660), .A2(KEYINPUT31), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n858), .B(new_n859), .C1(new_n860), .C2(new_n715), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n697), .A2(KEYINPUT92), .B1(new_n699), .B2(KEYINPUT30), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(new_n706), .A3(new_n713), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n858), .B1(new_n864), .B2(new_n859), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n691), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n717), .A2(new_n867), .B1(new_n689), .B2(new_n579), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n801), .B(new_n857), .C1(new_n866), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT104), .ZN(new_n870));
  INV_X1    g0670(.A(new_n624), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n652), .A2(new_n871), .A3(new_n660), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n629), .A2(new_n630), .A3(new_n674), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n660), .B1(new_n860), .B2(new_n715), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n691), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n874), .B(new_n876), .C1(new_n862), .C2(new_n865), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT104), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n877), .A2(new_n878), .A3(new_n801), .A4(new_n857), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT40), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  INV_X1    g0681(.A(new_n658), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n396), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n399), .A2(new_n883), .A3(new_n367), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n884), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n356), .A2(new_n369), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n883), .B1(new_n647), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n881), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n360), .A2(new_n330), .A3(new_n277), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n364), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n882), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n370), .B2(new_n403), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n891), .A2(new_n398), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(new_n892), .A3(new_n367), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n399), .A2(new_n883), .A3(new_n885), .A4(new_n367), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n880), .B1(new_n889), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n870), .A2(new_n879), .A3(new_n901), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n331), .A2(new_n353), .B1(new_n891), .B2(new_n398), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n885), .B1(new_n903), .B2(new_n892), .ZN(new_n904));
  AND4_X1   g0704(.A1(new_n885), .A2(new_n399), .A3(new_n883), .A4(new_n367), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n892), .B1(new_n647), .B2(new_n887), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n881), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n900), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n877), .A2(new_n909), .A3(new_n801), .A4(new_n857), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n880), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n902), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n627), .A2(new_n877), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(G330), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n912), .B2(new_n913), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT101), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n454), .B2(new_n852), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n855), .A2(KEYINPUT101), .A3(new_n851), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n918), .A2(new_n919), .B1(new_n852), .B2(new_n850), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n642), .A2(new_n661), .A3(new_n801), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(new_n921), .B2(new_n798), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n922), .A2(new_n909), .B1(new_n403), .B2(new_n658), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n909), .A2(KEYINPUT39), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n889), .A2(new_n925), .A3(new_n900), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(KEYINPUT102), .A3(new_n926), .ZN(new_n927));
  AOI211_X1 g0727(.A(KEYINPUT102), .B(new_n925), .C1(new_n908), .C2(new_n900), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n450), .A2(new_n660), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n923), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n627), .B1(new_n684), .B2(new_n686), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n650), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n933), .B(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n916), .A2(new_n937), .B1(new_n249), .B2(new_n726), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n916), .A2(new_n937), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n848), .B1(new_n938), .B2(new_n939), .ZN(G367));
  OAI21_X1  g0740(.A(new_n504), .B1(new_n475), .B2(new_n661), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n637), .A2(new_n660), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n675), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT44), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n675), .A2(new_n943), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT45), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n946), .B(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(KEYINPUT106), .A3(new_n672), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n671), .B(new_n673), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(new_n666), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n723), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n949), .A2(KEYINPUT106), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n945), .A2(new_n672), .A3(new_n948), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n672), .B1(new_n945), .B2(new_n948), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n722), .B1(new_n955), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n679), .B(KEYINPUT41), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n727), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n672), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n941), .A2(new_n539), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n660), .B1(new_n965), .B2(new_n503), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n671), .A2(new_n673), .A3(new_n943), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT42), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n661), .A2(new_n572), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n628), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n635), .B2(new_n972), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT105), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n971), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AND4_X1   g0780(.A1(new_n964), .A2(new_n977), .A3(new_n943), .A4(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n977), .A2(new_n980), .B1(new_n964), .B2(new_n943), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n963), .A2(new_n983), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n743), .B1(new_n207), .B2(new_n570), .C1(new_n231), .C2(new_n735), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n730), .ZN(new_n986));
  XOR2_X1   g0786(.A(KEYINPUT108), .B(G137), .Z(new_n987));
  NOR2_X1   g0787(.A1(new_n751), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n774), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n379), .A2(new_n989), .B1(new_n786), .B2(G150), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n267), .B2(new_n761), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n240), .B1(new_n758), .B2(new_n202), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G159), .B2(new_n771), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n767), .A2(new_n321), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G143), .B2(new_n783), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n992), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n765), .A2(new_n759), .B1(new_n767), .B2(new_n371), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n756), .A2(new_n588), .B1(new_n758), .B2(new_n826), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n315), .B1(new_n774), .B2(new_n460), .ZN(new_n1000));
  NOR3_X1   g0800(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(G317), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n762), .A2(G116), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT46), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n1003), .A2(new_n1004), .B1(new_n771), .B2(G294), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n1004), .B2(new_n1003), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT107), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1001), .B1(new_n1002), .B2(new_n751), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n997), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT47), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n986), .B1(new_n1011), .B2(new_n742), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n974), .A2(new_n793), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n984), .A2(new_n1014), .ZN(G387));
  INV_X1    g0815(.A(new_n727), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n668), .A2(new_n670), .A3(new_n741), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n678), .A2(new_n731), .B1(G107), .B2(new_n207), .ZN(new_n1018));
  AOI211_X1 g0818(.A(G45), .B(new_n677), .C1(G68), .C2(G77), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1020), .A2(KEYINPUT109), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(KEYINPUT109), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n264), .A2(G50), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT50), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n735), .B1(new_n228), .B2(G45), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1018), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n730), .B1(new_n1027), .B2(new_n744), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n752), .A2(G150), .B1(G97), .B2(new_n775), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n269), .B2(new_n770), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n240), .B1(new_n758), .B2(new_n321), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n761), .A2(new_n210), .B1(new_n756), .B2(new_n202), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n822), .A2(new_n380), .ZN(new_n1033));
  INV_X1    g0833(.A(G159), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n1034), .B2(new_n765), .ZN(new_n1035));
  NOR4_X1   g0835(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .A4(new_n1035), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT110), .Z(new_n1037));
  OAI22_X1  g0837(.A1(new_n770), .A2(new_n759), .B1(new_n765), .B2(new_n757), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1038), .A2(KEYINPUT111), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(KEYINPUT111), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G317), .A2(new_n786), .B1(new_n788), .B2(G303), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT48), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n761), .A2(new_n768), .B1(new_n767), .B2(new_n826), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1046));
  AOI21_X1  g0846(.A(KEYINPUT49), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1044), .A2(KEYINPUT49), .A3(new_n1046), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n240), .B1(new_n989), .B2(G116), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n766), .C2(new_n751), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1037), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1028), .B1(new_n1051), .B2(new_n742), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n952), .A2(new_n1016), .B1(new_n1017), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n679), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n953), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n723), .A2(new_n952), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(G393));
  NAND2_X1  g0857(.A1(new_n955), .A2(new_n960), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n959), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n957), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1058), .B(new_n1054), .C1(new_n1061), .C2(new_n954), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n943), .A2(new_n793), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n752), .A2(G322), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n315), .B1(new_n758), .B2(new_n768), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G283), .B2(new_n762), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n771), .A2(G303), .B1(new_n822), .B2(G116), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1064), .A2(new_n785), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n765), .A2(new_n1002), .B1(new_n756), .B2(new_n759), .ZN(new_n1069));
  XOR2_X1   g0869(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n1070));
  XNOR2_X1  g0870(.A(new_n1069), .B(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n752), .A2(G143), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n240), .B1(new_n758), .B2(new_n264), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G68), .B2(new_n762), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n822), .A2(G77), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G50), .B2(new_n771), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1072), .A2(new_n830), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n765), .A2(new_n815), .B1(new_n756), .B2(new_n1034), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT51), .Z(new_n1079));
  OAI22_X1  g0879(.A1(new_n1068), .A2(new_n1071), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n742), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n743), .B1(new_n460), .B2(new_n207), .C1(new_n238), .C2(new_n735), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1081), .A2(new_n730), .A3(new_n1082), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1062), .B1(new_n727), .B2(new_n1060), .C1(new_n1063), .C2(new_n1083), .ZN(G390));
  OAI21_X1  g0884(.A(new_n859), .B1(new_n860), .B2(new_n715), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(KEYINPUT103), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n861), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n875), .A2(new_n691), .B1(new_n872), .B2(new_n873), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n800), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1089), .A2(G330), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n857), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n660), .B(new_n800), .C1(new_n634), .C2(new_n641), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n857), .B1(new_n1092), .B2(new_n797), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n927), .A2(new_n929), .B1(new_n1093), .B2(new_n932), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n889), .A2(new_n900), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1093), .A2(new_n932), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1091), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n720), .A2(new_n801), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1098), .A2(new_n920), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1093), .A2(new_n932), .A3(new_n1095), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT102), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n909), .B2(KEYINPUT39), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n928), .B1(new_n1102), .B2(new_n926), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n922), .A2(new_n931), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1099), .B(new_n1100), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1097), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n1016), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n930), .A2(new_n739), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n761), .A2(new_n815), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT53), .ZN(new_n1110));
  INV_X1    g0910(.A(G128), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n1109), .A2(new_n1110), .B1(new_n1111), .B2(new_n765), .ZN(new_n1112));
  INV_X1    g0912(.A(G125), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n751), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n1034), .B2(new_n767), .ZN(new_n1116));
  INV_X1    g0916(.A(G132), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n240), .B1(new_n756), .B2(new_n1117), .C1(new_n202), .C2(new_n774), .ZN(new_n1118));
  OR4_X1    g0918(.A1(new_n1112), .A2(new_n1114), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT54), .B(G143), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n770), .A2(new_n987), .B1(new_n758), .B2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT113), .Z(new_n1122));
  AOI21_X1  g0922(.A(new_n1075), .B1(G283), .B2(new_n783), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n371), .B2(new_n770), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n752), .A2(G294), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n756), .A2(new_n594), .B1(new_n758), .B2(new_n460), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n240), .B(new_n1126), .C1(G87), .C2(new_n762), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1127), .A3(new_n819), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n1119), .A2(new_n1122), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n742), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n811), .A2(new_n308), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1108), .A2(new_n730), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1107), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(KEYINPUT114), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT114), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1107), .A2(new_n1135), .A3(new_n1132), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n627), .A2(G330), .A3(new_n877), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n934), .A2(new_n650), .A3(new_n1138), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1092), .A2(new_n797), .A3(new_n857), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1140), .A2(new_n922), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n1098), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1090), .B1(new_n1140), .B2(new_n922), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1139), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1106), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1145), .A2(new_n679), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1106), .A2(new_n1144), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1137), .A2(new_n1148), .ZN(G378));
  INV_X1    g0949(.A(KEYINPUT119), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n688), .B1(new_n910), .B2(new_n880), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n292), .A2(new_n882), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT55), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n307), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n307), .A2(new_n1155), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1153), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1158), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n1152), .A3(new_n1156), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n902), .A2(new_n1151), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1162), .B1(new_n902), .B2(new_n1151), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1163), .A2(new_n1164), .A3(new_n933), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n403), .A2(new_n658), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n909), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1166), .B1(new_n1093), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n1103), .B2(new_n931), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1162), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n879), .A2(new_n901), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n878), .B1(new_n1089), .B2(new_n857), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n911), .A2(G330), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1170), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n902), .A2(new_n1151), .A3(new_n1162), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1169), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(KEYINPUT57), .B1(new_n1165), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1139), .B1(new_n1106), .B2(new_n1144), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1150), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1139), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1147), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n933), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1175), .A2(new_n1169), .A3(new_n1176), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1182), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1180), .A2(new_n1054), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT118), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n1165), .B2(new_n1177), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1183), .A2(KEYINPUT118), .A3(new_n1184), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT57), .B1(new_n1191), .B2(new_n1182), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1187), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1170), .A2(new_n739), .ZN(new_n1194));
  AOI21_X1  g0994(.A(G50), .B1(new_n270), .B2(new_n250), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n240), .B2(G41), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT115), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G58), .A2(new_n989), .B1(new_n786), .B2(G107), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(new_n570), .B2(new_n758), .C1(new_n751), .C2(new_n826), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n250), .B(new_n315), .C1(new_n761), .C2(new_n210), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n770), .A2(new_n460), .B1(new_n765), .B2(new_n594), .ZN(new_n1201));
  NOR4_X1   g1001(.A1(new_n1199), .A2(new_n995), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1197), .B1(new_n1202), .B2(KEYINPUT58), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n770), .A2(new_n1117), .B1(new_n767), .B2(new_n815), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n788), .A2(G137), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n1111), .B2(new_n756), .C1(new_n761), .C2(new_n1120), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(G125), .C2(new_n783), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n752), .A2(G124), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G33), .B(G41), .C1(new_n989), .C2(G159), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT59), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1210), .B(new_n1211), .C1(new_n1207), .C2(new_n1212), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1203), .B1(KEYINPUT58), .B2(new_n1202), .C1(new_n1209), .C2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n742), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT116), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n728), .B(new_n1216), .C1(new_n202), .C2(new_n810), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1194), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1191), .B2(new_n1016), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1193), .A2(new_n1220), .ZN(G375));
  NAND2_X1  g1021(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n920), .A2(new_n739), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n730), .B1(new_n811), .B2(G68), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n752), .A2(G303), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n775), .A2(G77), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n240), .B1(new_n788), .B2(G107), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n762), .A2(G97), .B1(new_n786), .B2(G283), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1033), .B1(new_n765), .B2(new_n768), .C1(new_n594), .C2(new_n770), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n762), .A2(G159), .B1(new_n788), .B2(G150), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n756), .B2(new_n987), .C1(new_n751), .C2(new_n1111), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n783), .A2(G132), .B1(new_n822), .B2(G50), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n315), .B1(new_n989), .B2(G58), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1233), .B(new_n1234), .C1(new_n770), .C2(new_n1120), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n1229), .A2(new_n1230), .B1(new_n1232), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1224), .B1(new_n1236), .B2(new_n742), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1222), .A2(new_n1016), .B1(new_n1223), .B2(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1144), .A2(new_n962), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1222), .A2(new_n1181), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(G381));
  OR4_X1    g1041(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1242), .A2(G387), .A3(G381), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1134), .A2(new_n1136), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1244));
  INV_X1    g1044(.A(G375), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(G407));
  NAND2_X1  g1046(.A1(new_n659), .A2(G213), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT120), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1245), .A2(new_n1244), .A3(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(G407), .A2(new_n1249), .A3(G213), .ZN(G409));
  INV_X1    g1050(.A(KEYINPUT127), .ZN(new_n1251));
  OAI211_X1 g1051(.A(G378), .B(new_n1220), .C1(new_n1187), .C2(new_n1192), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n727), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(KEYINPUT121), .A3(new_n1218), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT121), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1253), .B2(new_n1219), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n962), .B(new_n1179), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1244), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1248), .B1(new_n1252), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1222), .A2(new_n1181), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1240), .B1(KEYINPUT60), .B2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1240), .A2(KEYINPUT60), .A3(new_n1262), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1054), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G384), .B(new_n1238), .C1(new_n1263), .C2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1238), .B1(new_n1265), .B2(new_n1263), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n835), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1261), .A2(KEYINPUT62), .A3(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1247), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n1273), .B(new_n1269), .C1(new_n1252), .C2(new_n1260), .ZN(new_n1274));
  OAI21_X1  g1074(.A(KEYINPUT126), .B1(new_n1274), .B2(KEYINPUT62), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1252), .A2(new_n1260), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1247), .A3(new_n1270), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT62), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1272), .B1(new_n1275), .B2(new_n1280), .ZN(new_n1281));
  XOR2_X1   g1081(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1269), .A2(G2897), .A3(new_n1248), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1273), .A2(G2897), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1266), .A2(new_n1268), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(KEYINPUT122), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT122), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1284), .A2(new_n1289), .A3(new_n1286), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1283), .B1(new_n1291), .B2(new_n1261), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1251), .B1(new_n1281), .B2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1273), .B1(new_n1252), .B2(new_n1260), .ZN(new_n1294));
  AOI211_X1 g1094(.A(KEYINPUT126), .B(KEYINPUT62), .C1(new_n1294), .C2(new_n1270), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1278), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1271), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1290), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1289), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1261), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1282), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1297), .A2(KEYINPUT127), .A3(new_n1302), .ZN(new_n1303));
  XOR2_X1   g1103(.A(G393), .B(G396), .Z(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  AOI22_X1  g1105(.A1(new_n963), .A2(new_n983), .B1(new_n1013), .B2(new_n1012), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT123), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1305), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(G387), .A2(new_n1304), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1308), .A2(new_n1309), .A3(G390), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G390), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1293), .A2(new_n1303), .A3(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT124), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  OAI211_X1 g1117(.A(KEYINPUT124), .B(new_n1314), .C1(new_n1310), .C2(new_n1311), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  OR2_X1    g1119(.A1(new_n1274), .A2(KEYINPUT63), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1261), .A2(KEYINPUT63), .A3(new_n1270), .ZN(new_n1321));
  OR2_X1    g1121(.A1(new_n1291), .A2(new_n1294), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .A4(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1313), .A2(new_n1323), .ZN(G405));
  NAND2_X1  g1124(.A1(G375), .A2(new_n1244), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1252), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1326), .B(new_n1270), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1327), .B(new_n1312), .ZN(G402));
endmodule


