//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n210), .B(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n206), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n208), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n217), .B1(KEYINPUT1), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XOR2_X1   g0039(.A(G58), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n206), .A2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G159), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AND2_X1   g0049(.A1(G58), .A2(G68), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G58), .A2(G68), .ZN(new_n251));
  OAI21_X1  g0051(.A(G20), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT71), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT71), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n254), .B(G20), .C1(new_n250), .C2(new_n251), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n249), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n246), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(new_n206), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT7), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT7), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n258), .A2(new_n262), .A3(new_n206), .A4(new_n259), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(G68), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n256), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT16), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n213), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n256), .A2(KEYINPUT16), .A3(new_n264), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G200), .ZN(new_n272));
  INV_X1    g0072(.A(G226), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G1698), .ZN(new_n274));
  AND2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n274), .B1(G223), .B2(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G87), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G1), .A3(G13), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n282), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n284), .B1(new_n288), .B2(G232), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n272), .B1(new_n281), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n286), .B1(new_n277), .B2(new_n278), .ZN(new_n291));
  INV_X1    g0091(.A(new_n282), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G274), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(new_n287), .B2(new_n220), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  NOR3_X1   g0095(.A1(new_n291), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  OR2_X1    g0097(.A1(KEYINPUT8), .A2(G58), .ZN(new_n298));
  NAND2_X1  g0098(.A1(KEYINPUT8), .A2(G58), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(new_n213), .A3(new_n268), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n205), .A2(G20), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n298), .A2(new_n303), .A3(new_n299), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n300), .A2(new_n301), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT72), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n271), .A2(new_n297), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT17), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n269), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(new_n265), .B2(new_n266), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n307), .B1(new_n313), .B2(new_n270), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n291), .A2(new_n294), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n291), .A2(new_n294), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT18), .B1(new_n314), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT18), .ZN(new_n322));
  INV_X1    g0122(.A(new_n319), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n316), .B2(new_n315), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n256), .A2(KEYINPUT16), .A3(new_n264), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT16), .B1(new_n256), .B2(new_n264), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n325), .A2(new_n326), .A3(new_n312), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n322), .B(new_n324), .C1(new_n327), .C2(new_n307), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n314), .A2(KEYINPUT17), .A3(new_n297), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n311), .A2(new_n321), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT15), .B(G87), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n206), .A2(G33), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n331), .A2(new_n332), .B1(new_n206), .B2(new_n202), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n298), .A2(new_n299), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n247), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n269), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n301), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n202), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n269), .B1(new_n205), .B2(G20), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G77), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n336), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G244), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n293), .B1(new_n287), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n258), .A2(new_n259), .ZN(new_n344));
  INV_X1    g0144(.A(G1698), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(G232), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(G238), .A3(G1698), .ZN(new_n347));
  INV_X1    g0147(.A(G107), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n346), .B(new_n347), .C1(new_n348), .C2(new_n344), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n343), .B1(new_n349), .B2(new_n280), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n341), .B1(new_n350), .B2(G169), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT67), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n341), .B(KEYINPUT67), .C1(new_n350), .C2(G169), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n350), .A2(new_n318), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n350), .A2(G190), .ZN(new_n357));
  INV_X1    g0157(.A(new_n341), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n357), .B(new_n358), .C1(new_n272), .C2(new_n350), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n330), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n293), .B1(new_n287), .B2(new_n273), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n344), .A2(G222), .A3(new_n345), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n344), .A2(G223), .A3(G1698), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n363), .B(new_n364), .C1(new_n202), .C2(new_n344), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n365), .A2(KEYINPUT66), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n286), .B1(new_n365), .B2(KEYINPUT66), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n362), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G190), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n334), .A2(new_n332), .ZN(new_n370));
  INV_X1    g0170(.A(G150), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n201), .A2(new_n206), .B1(new_n247), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n269), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n339), .A2(G50), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n373), .B(new_n374), .C1(G50), .C2(new_n301), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT9), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n369), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n368), .A2(new_n272), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT10), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n378), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT10), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n380), .A2(new_n381), .A3(new_n369), .A4(new_n376), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n368), .A2(new_n318), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n375), .B1(new_n368), .B2(G169), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n361), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n339), .A2(G68), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT12), .ZN(new_n390));
  INV_X1    g0190(.A(G68), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n337), .B2(new_n391), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n301), .A2(KEYINPUT12), .A3(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n389), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n332), .A2(new_n202), .B1(new_n206), .B2(G68), .ZN(new_n395));
  INV_X1    g0195(.A(G50), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n247), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n269), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT11), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n398), .A2(new_n399), .ZN(new_n401));
  OR3_X1    g0201(.A1(new_n394), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(G232), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n403));
  OAI211_X1 g0203(.A(G226), .B(new_n345), .C1(new_n275), .C2(new_n276), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G97), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n280), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n284), .B1(new_n288), .B2(G238), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(KEYINPUT13), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT13), .B1(new_n407), .B2(new_n408), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n402), .B1(new_n412), .B2(G200), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n407), .A2(new_n408), .B1(KEYINPUT68), .B2(KEYINPUT13), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT68), .A4(KEYINPUT13), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G190), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n416), .ZN(new_n420));
  OAI21_X1  g0220(.A(G179), .B1(new_n420), .B2(new_n414), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT70), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n417), .A2(KEYINPUT70), .A3(G179), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT69), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT14), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n412), .A2(G169), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n407), .A2(new_n408), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT13), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(G169), .A3(new_n409), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n427), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n419), .B1(new_n436), .B2(new_n402), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n388), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G45), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(G1), .ZN(new_n441));
  AND2_X1   g0241(.A1(KEYINPUT5), .A2(G41), .ZN(new_n442));
  NOR2_X1   g0242(.A1(KEYINPUT5), .A2(G41), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(G270), .A3(new_n286), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT5), .B(G41), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n446), .A2(G274), .A3(new_n286), .A4(new_n441), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(G264), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n449));
  OAI211_X1 g0249(.A(G257), .B(new_n345), .C1(new_n275), .C2(new_n276), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n258), .A2(G303), .A3(new_n259), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n280), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n316), .B1(new_n448), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n455), .B(new_n206), .C1(G33), .C2(new_n221), .ZN(new_n456));
  INV_X1    g0256(.A(G116), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G20), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n456), .A2(KEYINPUT20), .A3(new_n269), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT74), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n268), .A2(new_n213), .B1(G20), .B2(new_n457), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n462), .A2(KEYINPUT74), .A3(new_n456), .A4(KEYINPUT20), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n456), .A2(new_n269), .A3(new_n458), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT20), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n301), .A2(new_n457), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n205), .A2(G33), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n301), .A2(new_n469), .A3(new_n213), .A4(new_n268), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n471), .B2(new_n457), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n454), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT21), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n467), .A2(new_n472), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n448), .A2(G190), .A3(new_n453), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n445), .A2(new_n447), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n280), .B2(new_n452), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n477), .B(new_n478), .C1(new_n272), .C2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n454), .A2(new_n473), .A3(KEYINPUT21), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n473), .A2(new_n480), .A3(G179), .ZN(new_n483));
  AND4_X1   g0283(.A1(new_n476), .A2(new_n481), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  NOR3_X1   g0284(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n485));
  INV_X1    g0285(.A(new_n405), .ZN(new_n486));
  AND2_X1   g0286(.A1(KEYINPUT73), .A2(KEYINPUT19), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT73), .A2(KEYINPUT19), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n485), .B1(new_n489), .B2(new_n206), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n206), .B(G68), .C1(new_n275), .C2(new_n276), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n206), .A2(G33), .A3(G97), .ZN(new_n492));
  OR2_X1    g0292(.A1(KEYINPUT73), .A2(KEYINPUT19), .ZN(new_n493));
  NAND2_X1  g0293(.A1(KEYINPUT73), .A2(KEYINPUT19), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n269), .B1(new_n490), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n471), .A2(G87), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n331), .A2(new_n337), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(G244), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n501));
  OAI211_X1 g0301(.A(G238), .B(new_n345), .C1(new_n275), .C2(new_n276), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G116), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n504), .A2(new_n280), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n441), .A2(G274), .ZN(new_n506));
  OAI21_X1  g0306(.A(G250), .B1(new_n440), .B2(G1), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n506), .B1(new_n280), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(G200), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n508), .B1(new_n504), .B2(new_n280), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G190), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n500), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n497), .B(new_n499), .C1(new_n331), .C2(new_n470), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n510), .A2(new_n316), .ZN(new_n514));
  AOI211_X1 g0314(.A(new_n318), .B(new_n508), .C1(new_n504), .C2(new_n280), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n206), .B(G87), .C1(new_n275), .C2(new_n276), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT22), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT22), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n344), .A2(new_n520), .A3(new_n206), .A4(G87), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT24), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n503), .A2(G20), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT23), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n206), .B2(G107), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n348), .A2(KEYINPUT23), .A3(G20), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n522), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n523), .B1(new_n522), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n269), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n337), .A2(KEYINPUT25), .A3(new_n348), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT25), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n301), .B2(G107), .ZN(new_n534));
  AOI22_X1  g0334(.A1(G107), .A2(new_n471), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(G250), .B(new_n345), .C1(new_n275), .C2(new_n276), .ZN(new_n537));
  OAI211_X1 g0337(.A(G257), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n538));
  AND2_X1   g0338(.A1(KEYINPUT75), .A2(G294), .ZN(new_n539));
  NOR2_X1   g0339(.A1(KEYINPUT75), .A2(G294), .ZN(new_n540));
  OAI21_X1  g0340(.A(G33), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n537), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n280), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n280), .B1(new_n441), .B2(new_n446), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G264), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n545), .A3(new_n447), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n316), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n542), .A2(new_n280), .B1(new_n544), .B2(G264), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n548), .A2(new_n318), .A3(new_n447), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n536), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n517), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n546), .A2(G190), .ZN(new_n553));
  AOI21_X1  g0353(.A(G200), .B1(new_n548), .B2(new_n447), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n531), .B(new_n535), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(G244), .B(new_n345), .C1(new_n275), .C2(new_n276), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT4), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n344), .A2(KEYINPUT4), .A3(G244), .A4(new_n345), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n344), .A2(G250), .A3(G1698), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n455), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n280), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n444), .A2(new_n286), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n447), .B1(new_n563), .B2(new_n222), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n316), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n564), .B1(new_n561), .B2(new_n280), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n318), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n247), .A2(new_n202), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT6), .ZN(new_n571));
  AND2_X1   g0371(.A1(G97), .A2(G107), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G97), .A2(G107), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n348), .A2(KEYINPUT6), .A3(G97), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n570), .B1(new_n576), .B2(G20), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n261), .A2(G107), .A3(new_n263), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n269), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n301), .A2(G97), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n471), .B2(G97), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n567), .A2(new_n569), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n568), .A2(G190), .ZN(new_n585));
  INV_X1    g0385(.A(new_n582), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(new_n579), .B2(new_n269), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n585), .B(new_n587), .C1(new_n272), .C2(new_n568), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n555), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n552), .A2(new_n589), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n439), .A2(new_n484), .A3(new_n590), .ZN(G372));
  INV_X1    g0391(.A(new_n383), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n311), .A2(new_n329), .ZN(new_n593));
  INV_X1    g0393(.A(new_n402), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n425), .B2(new_n435), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n356), .B1(new_n413), .B2(new_n418), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n593), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n321), .A2(new_n328), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n592), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(KEYINPUT79), .B1(new_n600), .B2(new_n386), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT79), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n423), .A2(new_n424), .B1(new_n429), .B2(new_n434), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n594), .A2(new_n603), .B1(new_n419), .B2(new_n356), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n598), .B1(new_n604), .B2(new_n593), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n602), .B(new_n387), .C1(new_n605), .C2(new_n592), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n500), .A2(new_n509), .A3(new_n511), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT76), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n514), .B2(new_n515), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n510), .A2(G179), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n611), .B(KEYINPUT76), .C1(new_n316), .C2(new_n510), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n608), .B1(new_n613), .B2(new_n513), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT26), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT78), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n584), .A2(new_n616), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n566), .A2(new_n316), .B1(new_n580), .B2(new_n582), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(KEYINPUT78), .A3(new_n569), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n614), .A2(new_n615), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n513), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n610), .B2(new_n612), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n618), .A2(new_n569), .A3(new_n512), .A4(new_n516), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n622), .B1(new_n623), .B2(KEYINPUT26), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n584), .A2(new_n588), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(new_n555), .A3(new_n614), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n547), .A2(new_n549), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n531), .B2(new_n535), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT77), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n482), .A2(new_n483), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT21), .B1(new_n454), .B2(new_n473), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n476), .A2(KEYINPUT77), .A3(new_n482), .A4(new_n483), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n628), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n620), .B(new_n624), .C1(new_n626), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n439), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n607), .A2(new_n636), .ZN(G369));
  NAND3_X1  g0437(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(new_n640), .A3(G213), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G343), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n473), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n484), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n632), .A2(new_n633), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n646), .B1(new_n647), .B2(new_n645), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G330), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n555), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n536), .B2(new_n644), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(new_n628), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n628), .A2(new_n643), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n476), .A2(new_n482), .A3(new_n483), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n652), .A2(new_n658), .A3(new_n551), .A4(new_n643), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n654), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n657), .A2(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n209), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n485), .A2(new_n457), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G1), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n215), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  INV_X1    g0468(.A(G330), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n555), .A2(new_n584), .A3(new_n588), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n512), .A2(new_n516), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n628), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n670), .A2(new_n672), .A3(new_n484), .A4(new_n643), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT82), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT82), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n590), .A2(new_n675), .A3(new_n484), .A4(new_n643), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n548), .A2(new_n510), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT80), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT81), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT30), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n448), .A2(G179), .A3(new_n453), .A4(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT80), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n548), .A2(new_n510), .A3(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n679), .A2(new_n684), .A3(new_n568), .A4(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n680), .A2(new_n681), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n566), .A2(new_n683), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(new_n688), .A3(new_n686), .A4(new_n679), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n480), .A2(G179), .A3(new_n510), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n566), .A3(new_n546), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n690), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n644), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT31), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT31), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n698), .A3(new_n644), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n669), .B1(new_n677), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n670), .B(new_n614), .C1(new_n658), .C2(new_n628), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n617), .A2(new_n619), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n613), .A2(new_n513), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n512), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT26), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n623), .A2(KEYINPUT26), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n622), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n703), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n702), .B1(new_n710), .B2(new_n643), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n635), .A2(new_n702), .A3(new_n643), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n701), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n668), .B1(new_n713), .B2(G1), .ZN(G364));
  INV_X1    g0514(.A(G13), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n715), .A2(new_n440), .A3(G20), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n716), .A2(KEYINPUT83), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(KEYINPUT83), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G1), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n663), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n650), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(G330), .B2(new_n648), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n209), .A2(new_n344), .ZN(new_n723));
  INV_X1    g0523(.A(G355), .ZN(new_n724));
  OAI22_X1  g0524(.A1(new_n723), .A2(new_n724), .B1(G116), .B2(new_n209), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n241), .A2(G45), .ZN(new_n726));
  AOI211_X1 g0526(.A(new_n344), .B(new_n662), .C1(new_n440), .C2(new_n216), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n715), .A2(new_n246), .A3(KEYINPUT84), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT84), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(G13), .B2(G33), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n213), .B1(G20), .B2(new_n316), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n720), .B1(new_n728), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(G20), .A2(G179), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT85), .Z(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(G190), .A3(new_n272), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n740), .A2(new_n295), .A3(G200), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  XNOR2_X1  g0544(.A(KEYINPUT33), .B(G317), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G322), .A2(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT89), .Z(new_n747));
  NOR2_X1   g0547(.A1(new_n206), .A2(G179), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(new_n295), .A3(G200), .ZN(new_n749));
  INV_X1    g0549(.A(G283), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(new_n295), .A3(new_n272), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n344), .B1(new_n753), .B2(G329), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n539), .A2(new_n540), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n295), .A2(G179), .A3(G200), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n206), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n754), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n740), .A2(new_n295), .A3(new_n272), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n751), .B(new_n758), .C1(G311), .C2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n748), .A2(G190), .A3(G200), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT88), .Z(new_n763));
  NAND3_X1  g0563(.A1(new_n740), .A2(G190), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n763), .A2(G303), .B1(new_n765), .B2(G326), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n747), .A2(new_n761), .A3(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n757), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G97), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(new_n743), .B2(new_n391), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT87), .Z(new_n771));
  NOR2_X1   g0571(.A1(new_n752), .A2(new_n248), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(KEYINPUT32), .ZN(new_n774));
  INV_X1    g0574(.A(G87), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n774), .B1(new_n775), .B2(new_n762), .C1(new_n348), .C2(new_n749), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n344), .B1(new_n773), .B2(KEYINPUT32), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n396), .A2(new_n764), .B1(new_n759), .B2(new_n202), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n741), .B(KEYINPUT86), .Z(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n219), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n767), .B1(new_n771), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n738), .B1(new_n782), .B2(new_n735), .ZN(new_n783));
  INV_X1    g0583(.A(new_n734), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n783), .B1(new_n648), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n722), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(G396));
  NAND2_X1  g0587(.A1(new_n635), .A2(new_n643), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n358), .A2(new_n643), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n353), .A2(new_n354), .A3(new_n355), .A4(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(new_n360), .B2(new_n789), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n626), .A2(new_n634), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n620), .A2(new_n624), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n643), .B(new_n791), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n701), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n719), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(new_n664), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n701), .A2(new_n793), .A3(new_n796), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n720), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n732), .A2(new_n735), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(new_n202), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n344), .B1(new_n763), .B2(G107), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT90), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n749), .A2(new_n775), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n769), .B1(new_n808), .B2(new_n752), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n807), .B(new_n809), .C1(G116), .C2(new_n760), .ZN(new_n810));
  INV_X1    g0610(.A(G294), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n750), .A2(new_n743), .B1(new_n741), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G303), .B2(new_n765), .ZN(new_n813));
  AND3_X1   g0613(.A1(new_n806), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G150), .A2(new_n744), .B1(new_n760), .B2(G159), .ZN(new_n815));
  INV_X1    g0615(.A(G137), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n816), .B2(new_n764), .ZN(new_n817));
  INV_X1    g0617(.A(new_n780), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(G143), .B2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT34), .Z(new_n820));
  NOR2_X1   g0620(.A1(new_n275), .A2(new_n276), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n753), .B2(G132), .ZN(new_n822));
  INV_X1    g0622(.A(new_n749), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G68), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n822), .B(new_n824), .C1(new_n219), .C2(new_n757), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G50), .B2(new_n763), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n814), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n735), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n804), .B1(new_n733), .B2(new_n791), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT91), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n801), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G384));
  NAND2_X1  g0632(.A1(new_n214), .A2(G116), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n576), .B2(KEYINPUT35), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(KEYINPUT35), .B2(new_n576), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT36), .ZN(new_n836));
  OAI21_X1  g0636(.A(G77), .B1(new_n219), .B2(new_n391), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n837), .A2(new_n215), .B1(G50), .B2(new_n391), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(G1), .A3(new_n715), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT92), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT37), .ZN(new_n842));
  INV_X1    g0642(.A(new_n305), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n271), .A2(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n844), .A2(new_n642), .B1(new_n314), .B2(new_n297), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n324), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n324), .B1(new_n327), .B2(new_n307), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n642), .B1(new_n327), .B2(new_n307), .ZN(new_n849));
  AND4_X1   g0649(.A1(new_n842), .A2(new_n848), .A3(new_n849), .A4(new_n309), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT93), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n305), .B1(new_n313), .B2(new_n270), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n309), .B1(new_n641), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n320), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT37), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT93), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n848), .A2(new_n849), .A3(new_n842), .A4(new_n309), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n852), .A2(new_n641), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n330), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n851), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n851), .A2(KEYINPUT38), .A3(new_n858), .A4(new_n860), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(KEYINPUT39), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n848), .A2(new_n849), .A3(new_n309), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n857), .ZN(new_n868));
  INV_X1    g0668(.A(new_n849), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n330), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n862), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT39), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n865), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n595), .A2(new_n643), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n599), .A2(new_n642), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n863), .A2(new_n864), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n402), .A2(new_n644), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n603), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n437), .B2(new_n881), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n356), .A2(new_n644), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n883), .B1(new_n796), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n879), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT94), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n876), .A2(new_n878), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n439), .B1(new_n711), .B2(new_n712), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n607), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n891), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n677), .A2(new_n700), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT40), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n863), .A2(new_n896), .A3(new_n864), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n674), .A2(new_n676), .B1(new_n697), .B2(new_n699), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n413), .A2(new_n418), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n899), .B(new_n881), .C1(new_n603), .C2(new_n594), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n436), .A2(new_n402), .A3(new_n644), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n791), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT95), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n904), .A2(new_n896), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n898), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n897), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT95), .B1(new_n898), .B2(new_n903), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n896), .B1(new_n908), .B2(new_n873), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n439), .B(new_n895), .C1(new_n907), .C2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n792), .B1(new_n900), .B2(new_n901), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n904), .B1(new_n895), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n873), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT40), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n897), .A2(new_n906), .ZN(new_n915));
  INV_X1    g0715(.A(new_n439), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n914), .B(new_n915), .C1(new_n916), .C2(new_n898), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n910), .A2(new_n917), .A3(G330), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n894), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(G1), .B1(new_n715), .B2(G20), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n894), .A2(new_n918), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n841), .B1(new_n921), .B2(new_n922), .ZN(G367));
  OAI21_X1  g0723(.A(new_n625), .B1(new_n587), .B2(new_n643), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n618), .A2(new_n569), .A3(new_n644), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT98), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n657), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n500), .A2(new_n643), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n706), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(KEYINPUT96), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n930), .A2(KEYINPUT96), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n931), .B(new_n932), .C1(new_n622), .C2(new_n929), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT97), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n933), .B(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT43), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n927), .A2(new_n551), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n644), .B1(new_n939), .B2(new_n584), .ZN(new_n940));
  INV_X1    g0740(.A(new_n926), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n941), .A2(new_n659), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT42), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n935), .A2(KEYINPUT43), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n938), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n944), .A2(new_n936), .A3(KEYINPUT99), .A4(new_n937), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT99), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n938), .B2(new_n945), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n928), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n951), .A2(new_n947), .A3(new_n928), .A4(new_n948), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(KEYINPUT100), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT100), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n949), .A2(new_n955), .A3(new_n928), .A4(new_n951), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n952), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT45), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n660), .A2(new_n926), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT101), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n959), .A2(KEYINPUT101), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n962), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(KEYINPUT45), .A3(new_n960), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n660), .A2(new_n926), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT44), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n963), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n657), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n658), .A2(new_n643), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n653), .B2(new_n655), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n659), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(KEYINPUT102), .B2(new_n649), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n649), .B(KEYINPUT102), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n974), .B1(new_n975), .B2(new_n973), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n713), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n963), .A2(new_n965), .A3(new_n657), .A4(new_n967), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n970), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n980), .A2(new_n713), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n663), .B(KEYINPUT41), .Z(new_n982));
  OAI21_X1  g0782(.A(new_n798), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n957), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n662), .A2(new_n344), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n985), .A2(new_n236), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n736), .B1(new_n209), .B2(new_n331), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n750), .A2(new_n759), .B1(new_n743), .B2(new_n755), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n344), .B1(new_n753), .B2(G317), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n221), .B2(new_n749), .C1(new_n348), .C2(new_n757), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n988), .B(new_n990), .C1(G311), .C2(new_n765), .ZN(new_n991));
  INV_X1    g0791(.A(G303), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT46), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n763), .B2(G116), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n762), .A2(KEYINPUT46), .A3(new_n457), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n991), .B1(new_n992), .B2(new_n780), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n752), .A2(new_n816), .B1(new_n762), .B2(new_n219), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n741), .A2(new_n371), .B1(new_n997), .B2(KEYINPUT103), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G143), .B2(new_n765), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n768), .A2(G68), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n1000), .B(new_n344), .C1(new_n202), .C2(new_n749), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G159), .B2(new_n744), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n760), .A2(G50), .B1(new_n997), .B2(KEYINPUT103), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n999), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n996), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT47), .Z(new_n1006));
  OAI221_X1 g0806(.A(new_n720), .B1(new_n986), .B2(new_n987), .C1(new_n1006), .C2(new_n828), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT104), .Z(new_n1008));
  NAND2_X1  g0808(.A1(new_n936), .A2(new_n734), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n984), .A2(new_n1010), .ZN(G387));
  OR3_X1    g0811(.A1(new_n976), .A2(new_n713), .A3(KEYINPUT108), .ZN(new_n1012));
  OAI21_X1  g0812(.A(KEYINPUT108), .B1(new_n976), .B2(new_n713), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1012), .A2(new_n663), .A3(new_n977), .A4(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n440), .B1(new_n391), .B2(new_n202), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT105), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1015), .B1(new_n665), .B2(new_n1016), .ZN(new_n1017));
  AND3_X1   g0817(.A1(new_n300), .A2(KEYINPUT50), .A3(new_n396), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT50), .B1(new_n300), .B2(new_n396), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1017), .B1(new_n1016), .B2(new_n665), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n985), .B(new_n1020), .C1(new_n233), .C2(new_n440), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(G107), .B2(new_n209), .C1(new_n665), .C2(new_n723), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n802), .B1(new_n1022), .B2(new_n736), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n656), .B2(new_n784), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n344), .B1(new_n752), .B2(new_n371), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n762), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(G77), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n331), .B2(new_n757), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1025), .B(new_n1028), .C1(G97), .C2(new_n823), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n248), .A2(new_n764), .B1(new_n743), .B2(new_n334), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G68), .B2(new_n760), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1029), .B(new_n1031), .C1(new_n396), .C2(new_n741), .ZN(new_n1032));
  XOR2_X1   g0832(.A(KEYINPUT106), .B(G322), .Z(new_n1033));
  NAND2_X1  g0833(.A1(new_n765), .A2(new_n1033), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n992), .B2(new_n759), .C1(new_n808), .C2(new_n743), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n818), .B2(G317), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1036), .A2(KEYINPUT48), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(KEYINPUT48), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n757), .A2(new_n750), .B1(new_n762), .B2(new_n755), .ZN(new_n1039));
  OR3_X1    g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  XOR2_X1   g0840(.A(KEYINPUT107), .B(KEYINPUT49), .Z(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n344), .B1(new_n753), .B2(G326), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(new_n457), .C2(new_n749), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1032), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1024), .B1(new_n1046), .B2(new_n735), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n976), .B2(new_n719), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1014), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(KEYINPUT109), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT109), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1014), .A2(new_n1051), .A3(new_n1048), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(G393));
  INV_X1    g0853(.A(KEYINPUT110), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n970), .A2(new_n1054), .A3(new_n979), .ZN(new_n1055));
  OR3_X1    g0855(.A1(new_n968), .A2(new_n1054), .A3(new_n969), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n663), .B(new_n980), .C1(new_n1057), .C2(new_n978), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n927), .A2(new_n734), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT111), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n985), .A2(new_n244), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n736), .B1(new_n221), .B2(new_n209), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n749), .A2(new_n348), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n344), .B(new_n1063), .C1(new_n753), .C2(new_n1033), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n750), .B2(new_n762), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G294), .B2(new_n760), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT113), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n744), .A2(G303), .B1(G116), .B2(new_n768), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G311), .A2(new_n742), .B1(new_n765), .B2(G317), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1071), .B(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n371), .A2(new_n764), .B1(new_n741), .B2(new_n248), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT51), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n821), .B(new_n807), .C1(G143), .C2(new_n753), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n768), .A2(G77), .B1(new_n1026), .B2(G68), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(new_n334), .C2(new_n759), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G50), .B2(new_n744), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1070), .A2(new_n1073), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n720), .B1(new_n1061), .B2(new_n1062), .C1(new_n1080), .C2(new_n828), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1060), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n1057), .B2(new_n719), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1058), .A2(new_n1083), .ZN(G390));
  AOI22_X1  g0884(.A1(new_n763), .A2(G87), .B1(new_n765), .B2(G283), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n348), .B2(new_n743), .C1(new_n457), .C2(new_n741), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n821), .B1(new_n752), .B2(new_n811), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G68), .B2(new_n823), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n202), .B2(new_n757), .C1(new_n221), .C2(new_n759), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G132), .A2(new_n742), .B1(new_n744), .B2(G137), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n762), .A2(new_n371), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT53), .ZN(new_n1092));
  INV_X1    g0892(.A(G128), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1090), .B(new_n1092), .C1(new_n1093), .C2(new_n764), .ZN(new_n1094));
  XOR2_X1   g0894(.A(KEYINPUT54), .B(G143), .Z(new_n1095));
  NAND2_X1  g0895(.A1(new_n760), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n768), .A2(G159), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n823), .A2(G50), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n821), .B1(new_n753), .B2(G125), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1086), .A2(new_n1089), .B1(new_n1094), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n735), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n802), .B1(new_n334), .B2(new_n803), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n865), .A2(new_n875), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n732), .ZN(new_n1106));
  NOR4_X1   g0906(.A1(new_n898), .A2(new_n669), .A3(new_n883), .A4(new_n792), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n796), .A2(new_n885), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n902), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n875), .A2(new_n865), .B1(new_n1109), .B2(new_n877), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n873), .A2(new_n877), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n710), .A2(new_n643), .A3(new_n791), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n902), .A2(KEYINPUT114), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT114), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n900), .A2(new_n901), .A3(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1112), .A2(new_n885), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1107), .B1(new_n1110), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1109), .A2(new_n877), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1105), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n895), .A2(G330), .A3(new_n791), .A4(new_n902), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1118), .A2(new_n1123), .A3(new_n719), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(KEYINPUT116), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT116), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1118), .A2(new_n1123), .A3(new_n1126), .A4(new_n719), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1106), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n701), .A2(new_n439), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n607), .A2(new_n892), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n902), .B1(new_n701), .B2(new_n791), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1108), .B1(new_n1131), .B2(new_n1107), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1112), .A2(new_n885), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n898), .A2(new_n669), .A3(new_n792), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1121), .B(new_n1133), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1130), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1137), .A2(new_n1118), .A3(new_n1123), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT115), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n1139), .A3(new_n663), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1118), .A2(new_n1123), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1137), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1139), .B1(new_n1138), .B2(new_n663), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1128), .B1(new_n1144), .B2(new_n1145), .ZN(G378));
  INV_X1    g0946(.A(new_n1130), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1138), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(G330), .B1(new_n907), .B2(new_n909), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n889), .A2(new_n1149), .A3(new_n890), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n669), .B1(new_n914), .B2(new_n915), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n879), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n855), .A2(new_n857), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1153), .A2(KEYINPUT93), .B1(new_n330), .B2(new_n859), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT38), .B1(new_n1154), .B2(new_n858), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n864), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n888), .B(new_n1152), .C1(new_n1157), .C2(new_n1109), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n865), .A2(new_n875), .A3(new_n878), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n887), .A2(new_n888), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1151), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n375), .A2(new_n642), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n592), .A2(new_n386), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1163), .B1(new_n383), .B2(new_n387), .ZN(new_n1166));
  OR3_X1    g0966(.A1(new_n1165), .A2(KEYINPUT119), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(KEYINPUT119), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g0969(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1167), .A2(new_n1170), .A3(new_n1168), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1150), .A2(new_n1162), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1150), .B2(new_n1162), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1148), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT57), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1148), .B(KEYINPUT57), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n663), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1150), .A2(new_n1162), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n1174), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1150), .A2(new_n1162), .A3(new_n1175), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n798), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1174), .A2(new_n733), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n802), .B1(new_n396), .B2(new_n803), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n768), .A2(G150), .B1(new_n1026), .B2(new_n1095), .ZN(new_n1189));
  INV_X1    g0989(.A(G132), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1189), .B1(new_n1190), .B2(new_n743), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n1093), .A2(new_n741), .B1(new_n759), .B2(new_n816), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(G125), .C2(new_n765), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1196));
  AOI211_X1 g0996(.A(G33), .B(G41), .C1(new_n753), .C2(G124), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n248), .B2(new_n749), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT118), .Z(new_n1199));
  NAND3_X1  g0999(.A1(new_n1195), .A2(new_n1196), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1000), .B1(new_n764), .B2(new_n457), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT117), .Z(new_n1202));
  NOR2_X1   g1002(.A1(new_n743), .A2(new_n221), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n749), .A2(new_n219), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n753), .A2(G283), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n344), .A2(G41), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1205), .A2(new_n1027), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n348), .A2(new_n741), .B1(new_n759), .B2(new_n331), .ZN(new_n1209));
  NOR4_X1   g1009(.A1(new_n1202), .A2(new_n1203), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1210), .A2(KEYINPUT58), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(KEYINPUT58), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n396), .B1(new_n275), .B2(G41), .ZN(new_n1213));
  AND4_X1   g1013(.A1(new_n1200), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1188), .B1(new_n1214), .B2(new_n828), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1187), .A2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1186), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1182), .A2(new_n1217), .ZN(G375));
  AND2_X1   g1018(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1130), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n982), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1220), .A2(new_n1221), .A3(new_n1142), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n821), .B(new_n1204), .C1(G128), .C2(new_n753), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n763), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1223), .B1(new_n396), .B2(new_n757), .C1(new_n1224), .C2(new_n248), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n744), .A2(new_n1095), .B1(new_n765), .B2(G132), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n371), .B2(new_n759), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1225), .B(new_n1227), .C1(G137), .C2(new_n818), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n821), .B1(new_n749), .B2(new_n202), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT120), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n331), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n768), .A2(new_n1231), .B1(new_n753), .B2(G303), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1230), .B(new_n1232), .C1(new_n457), .C2(new_n743), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1224), .A2(new_n221), .B1(new_n811), .B2(new_n764), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n348), .A2(new_n759), .B1(new_n741), .B2(new_n750), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n735), .B1(new_n1228), .B2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n802), .B1(new_n391), .B2(new_n803), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1237), .B(new_n1238), .C1(new_n1135), .C2(new_n733), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n1219), .B2(new_n798), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1222), .A2(new_n1241), .ZN(G381));
  INV_X1    g1042(.A(G378), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1182), .A2(new_n1243), .A3(new_n1217), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n957), .A2(new_n983), .B1(new_n1009), .B2(new_n1008), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(G390), .A2(G384), .A3(G381), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1050), .A2(new_n786), .A3(new_n1052), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1249), .ZN(G407));
  OAI211_X1 g1050(.A(G407), .B(G213), .C1(G343), .C2(new_n1244), .ZN(G409));
  AOI21_X1  g1051(.A(new_n786), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1058), .B(new_n1083), .C1(new_n1249), .C2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1252), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(G390), .A3(new_n1248), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(G387), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1246), .A2(new_n1255), .A3(new_n1253), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(G375), .A2(G378), .ZN(new_n1261));
  INV_X1    g1061(.A(G343), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(G213), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT121), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1186), .B2(new_n1216), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n719), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1216), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(KEYINPUT121), .A3(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1148), .B(new_n1221), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1265), .A2(new_n1243), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1261), .A2(KEYINPUT124), .A3(new_n1263), .A4(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT124), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1270), .A2(new_n1263), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1243), .B1(new_n1182), .B2(new_n1217), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1272), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1219), .A2(KEYINPUT60), .A3(new_n1130), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT123), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1276), .B(new_n1277), .ZN(new_n1278));
  XOR2_X1   g1078(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n1279));
  NAND2_X1  g1079(.A1(new_n1220), .A2(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1137), .A2(new_n664), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AOI211_X1 g1082(.A(new_n831), .B(new_n1240), .C1(new_n1278), .C2(new_n1282), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1280), .B(new_n1281), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G384), .B1(new_n1286), .B2(new_n1241), .ZN(new_n1287));
  INV_X1    g1087(.A(G2897), .ZN(new_n1288));
  OAI22_X1  g1088(.A1(new_n1283), .A2(new_n1287), .B1(new_n1288), .B2(new_n1263), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1276), .B(KEYINPUT123), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1241), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n831), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1286), .A2(G384), .A3(new_n1241), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1263), .A2(new_n1288), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1289), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1271), .A2(new_n1275), .A3(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1283), .A2(new_n1287), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1261), .A2(new_n1263), .A3(new_n1299), .A4(new_n1270), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT63), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1273), .A2(new_n1274), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(KEYINPUT63), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1260), .A2(new_n1298), .A3(new_n1302), .A4(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1297), .B1(new_n1274), .B2(new_n1273), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1259), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT125), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1311), .B1(new_n1304), .B2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1300), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1308), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1306), .B1(new_n1315), .B2(new_n1317), .ZN(G405));
  INV_X1    g1118(.A(KEYINPUT126), .ZN(new_n1319));
  OAI21_X1  g1119(.A(KEYINPUT127), .B1(new_n1303), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT127), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1299), .A2(KEYINPUT126), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1323), .A2(new_n1244), .A3(new_n1261), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1320), .B(new_n1322), .C1(new_n1245), .C2(new_n1274), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1316), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1317), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(G402));
endmodule


