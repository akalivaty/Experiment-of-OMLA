//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT70), .A2(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT70), .A2(G953), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G227), .ZN(new_n192));
  XOR2_X1   g006(.A(G110), .B(G140), .Z(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G134), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n199), .B1(G134), .B2(new_n196), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  NOR3_X1   g015(.A1(new_n201), .A2(KEYINPUT11), .A3(G137), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n198), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G131), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT11), .B1(new_n201), .B2(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n199), .A2(new_n196), .A3(G134), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n197), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n212), .A2(new_n214), .A3(new_n215), .A4(G128), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT82), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n213), .A2(G146), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n218), .B1(new_n219), .B2(new_n215), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n212), .A2(KEYINPUT82), .A3(KEYINPUT1), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(G128), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n212), .A2(new_n214), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n217), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT80), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(KEYINPUT80), .ZN(new_n227));
  INV_X1    g041(.A(G107), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G104), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n226), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G101), .ZN(new_n231));
  INV_X1    g045(.A(G104), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G107), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT80), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(KEYINPUT3), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n232), .A2(G107), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n230), .A2(new_n231), .A3(new_n233), .A4(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n229), .A2(new_n233), .A3(KEYINPUT81), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n239), .B(G101), .C1(KEYINPUT81), .C2(new_n229), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n224), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT64), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n243), .B1(new_n211), .B2(G143), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n213), .A2(KEYINPUT64), .A3(G146), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n219), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G128), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n247), .B1(new_n212), .B2(KEYINPUT1), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n216), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n238), .B2(new_n240), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n210), .B1(new_n242), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT12), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI211_X1 g067(.A(KEYINPUT12), .B(new_n210), .C1(new_n242), .C2(new_n250), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n234), .A2(KEYINPUT3), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n235), .B1(new_n236), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n233), .B1(new_n226), .B2(new_n229), .ZN(new_n258));
  OAI21_X1  g072(.A(G101), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT4), .A3(new_n238), .ZN(new_n260));
  AND2_X1   g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n212), .A2(new_n214), .A3(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n262), .B1(new_n246), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT69), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n268), .B(new_n262), .C1(new_n246), .C2(new_n265), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n270), .B(G101), .C1(new_n257), .C2(new_n258), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n260), .A2(new_n267), .A3(new_n269), .A4(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n241), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(KEYINPUT10), .A3(new_n249), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(new_n224), .B2(new_n241), .ZN(new_n276));
  INV_X1    g090(.A(new_n210), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n272), .A2(new_n274), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT84), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n278), .A2(new_n279), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n255), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT85), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT85), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n284), .B(new_n255), .C1(new_n280), .C2(new_n281), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n195), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G469), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n272), .A2(new_n274), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n288), .A2(KEYINPUT84), .A3(new_n277), .A4(new_n276), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n278), .A2(new_n279), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n194), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n272), .A2(new_n274), .A3(new_n276), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n210), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n286), .A2(new_n287), .A3(new_n295), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n195), .B(new_n255), .C1(new_n280), .C2(new_n281), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n289), .A2(new_n290), .B1(new_n210), .B2(new_n292), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n298), .B2(new_n195), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n287), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n287), .A2(new_n300), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n188), .B1(new_n296), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT93), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT13), .B1(new_n247), .B2(G143), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(new_n201), .ZN(new_n308));
  XNOR2_X1  g122(.A(G128), .B(G143), .ZN(new_n309));
  XOR2_X1   g123(.A(new_n308), .B(new_n309), .Z(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G122), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G116), .ZN(new_n313));
  INV_X1    g127(.A(G116), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G122), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT91), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT91), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(G107), .ZN(new_n319));
  INV_X1    g133(.A(new_n318), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n228), .B1(new_n320), .B2(new_n316), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT92), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n322), .B1(new_n319), .B2(new_n321), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n311), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n309), .B(new_n201), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n314), .A2(KEYINPUT14), .A3(G122), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n313), .A2(new_n315), .ZN(new_n329));
  OAI211_X1 g143(.A(G107), .B(new_n328), .C1(new_n329), .C2(KEYINPUT14), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n321), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT75), .B(G217), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n332), .A2(new_n187), .A3(G953), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n326), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n333), .ZN(new_n335));
  AOI21_X1  g149(.A(G107), .B1(new_n317), .B2(new_n318), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n320), .A2(new_n228), .A3(new_n316), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT92), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n310), .B1(new_n338), .B2(new_n323), .ZN(new_n339));
  INV_X1    g153(.A(new_n331), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n335), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI211_X1 g155(.A(new_n306), .B(G902), .C1(new_n334), .C2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G478), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(KEYINPUT15), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n334), .A2(new_n341), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n300), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n306), .ZN(new_n349));
  AOI21_X1  g163(.A(G902), .B1(new_n334), .B2(new_n341), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT93), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n346), .B1(new_n352), .B2(new_n345), .ZN(new_n353));
  INV_X1    g167(.A(G952), .ZN(new_n354));
  AOI211_X1 g168(.A(G953), .B(new_n354), .C1(G234), .C2(G237), .ZN(new_n355));
  AOI211_X1 g169(.A(new_n300), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT21), .B(G898), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G113), .B(G122), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(new_n232), .ZN(new_n361));
  INV_X1    g175(.A(G125), .ZN(new_n362));
  NOR3_X1   g176(.A1(new_n362), .A2(KEYINPUT16), .A3(G140), .ZN(new_n363));
  XNOR2_X1  g177(.A(G125), .B(G140), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n363), .B1(new_n364), .B2(KEYINPUT16), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G146), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  XOR2_X1   g181(.A(G125), .B(G140), .Z(new_n368));
  INV_X1    g182(.A(KEYINPUT19), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n364), .A2(KEYINPUT19), .ZN(new_n371));
  AOI21_X1  g185(.A(G146), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G237), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n191), .A2(G143), .A3(G214), .A4(new_n374), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n189), .A2(G214), .A3(new_n374), .A4(new_n190), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n213), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n208), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n208), .B1(new_n375), .B2(new_n377), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n373), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(KEYINPUT18), .A2(G131), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(new_n375), .B2(new_n377), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n368), .A2(G146), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n364), .A2(new_n211), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n375), .A2(new_n377), .A3(new_n382), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n384), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n361), .B1(new_n381), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n387), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(new_n383), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n366), .A2(KEYINPUT76), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n365), .A2(G146), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT76), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n365), .A2(new_n395), .A3(G146), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT17), .ZN(new_n398));
  AOI211_X1 g212(.A(new_n398), .B(new_n208), .C1(new_n375), .C2(new_n377), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n380), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n398), .A3(new_n378), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n392), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n390), .B1(new_n403), .B2(new_n361), .ZN(new_n404));
  NOR2_X1   g218(.A1(G475), .A2(G902), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT20), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n402), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n380), .A2(KEYINPUT17), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n409), .A2(new_n393), .A3(new_n394), .A4(new_n396), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n361), .B(new_n389), .C1(new_n408), .C2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n390), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT20), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(new_n405), .ZN(new_n415));
  INV_X1    g229(.A(new_n411), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n403), .A2(new_n361), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n300), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n407), .A2(new_n415), .B1(new_n418), .B2(G475), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n353), .A2(new_n359), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n305), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(G210), .B1(G237), .B2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n362), .B(new_n216), .C1(new_n246), .C2(new_n248), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n212), .A2(new_n214), .A3(new_n261), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n213), .A2(KEYINPUT64), .A3(G146), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT64), .B1(new_n213), .B2(G146), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n212), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n425), .B1(new_n428), .B2(new_n264), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n424), .B1(new_n429), .B2(new_n362), .ZN(new_n430));
  INV_X1    g244(.A(G953), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G224), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT7), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT87), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n430), .A2(new_n436), .A3(new_n433), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  XOR2_X1   g252(.A(KEYINPUT86), .B(KEYINPUT8), .Z(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G122), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G113), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n314), .A2(G119), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT5), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT67), .ZN(new_n446));
  INV_X1    g260(.A(G119), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n446), .B1(new_n447), .B2(G116), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n314), .A2(KEYINPUT67), .A3(G119), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(G116), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n445), .B1(new_n452), .B2(new_n444), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n442), .A2(KEYINPUT2), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT2), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G113), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n443), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT68), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n457), .A2(new_n458), .A3(new_n450), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n458), .B1(new_n457), .B2(new_n450), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n453), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(new_n241), .ZN(new_n462));
  INV_X1    g276(.A(new_n450), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n455), .A2(G113), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n442), .A2(KEYINPUT2), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n451), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT68), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n457), .A2(new_n458), .A3(new_n450), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n469), .A2(new_n453), .B1(new_n238), .B2(new_n240), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n441), .B1(new_n462), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n273), .A2(new_n469), .A3(new_n453), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n464), .A2(new_n465), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n467), .A2(new_n468), .B1(new_n452), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n260), .A2(new_n271), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n472), .B(new_n440), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n430), .A2(new_n433), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n438), .A2(new_n471), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(KEYINPUT88), .A3(new_n300), .ZN(new_n479));
  OAI22_X1  g293(.A1(new_n475), .A2(new_n474), .B1(new_n461), .B2(new_n241), .ZN(new_n480));
  INV_X1    g294(.A(new_n440), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(KEYINPUT6), .A3(new_n476), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT6), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n480), .A2(new_n484), .A3(new_n481), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n430), .B(new_n432), .Z(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n479), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT88), .B1(new_n478), .B2(new_n300), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n423), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT89), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n478), .A2(new_n300), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT88), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n495), .A2(new_n422), .A3(new_n487), .A4(new_n479), .ZN(new_n496));
  OAI211_X1 g310(.A(KEYINPUT89), .B(new_n423), .C1(new_n488), .C2(new_n489), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n492), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n499));
  OAI21_X1  g313(.A(G214), .B1(G237), .B2(G902), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n498), .B2(new_n500), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n421), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n267), .A2(new_n210), .A3(new_n269), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n196), .B2(G134), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT65), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n201), .B2(G137), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n201), .A2(KEYINPUT66), .A3(G137), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n196), .A2(KEYINPUT65), .A3(G134), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n506), .A2(new_n508), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(G131), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n249), .A2(new_n209), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n504), .A2(new_n474), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n504), .A2(new_n513), .ZN(new_n517));
  INV_X1    g331(.A(new_n474), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n514), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n516), .B1(new_n520), .B2(KEYINPUT28), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n191), .A2(G210), .A3(new_n374), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT27), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT26), .B(G101), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT29), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(G902), .B1(new_n521), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n512), .A2(new_n209), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n530), .A2(new_n249), .B1(new_n210), .B2(new_n429), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT71), .B1(new_n531), .B2(new_n474), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n210), .A2(new_n429), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n513), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT71), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(new_n518), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(new_n514), .A3(new_n536), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n537), .A2(KEYINPUT72), .A3(KEYINPUT28), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT72), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n539), .B1(new_n514), .B2(new_n515), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n537), .B2(KEYINPUT28), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n538), .A2(new_n541), .A3(new_n526), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT30), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n534), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n504), .A2(KEYINPUT30), .A3(new_n513), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n518), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n514), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n526), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n527), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n529), .B1(new_n542), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G472), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT32), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n526), .B1(new_n538), .B2(new_n541), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n546), .A2(new_n525), .A3(new_n514), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT31), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n546), .A2(KEYINPUT31), .A3(new_n525), .A4(new_n514), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(G472), .A2(G902), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT73), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n552), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  AOI211_X1 g377(.A(KEYINPUT32), .B(new_n561), .C1(new_n553), .C2(new_n558), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n551), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT74), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT23), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n447), .B2(G128), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n247), .A2(KEYINPUT23), .A3(G119), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n568), .B(new_n569), .C1(G119), .C2(new_n247), .ZN(new_n570));
  XNOR2_X1  g384(.A(G119), .B(G128), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT24), .B(G110), .Z(new_n572));
  AOI22_X1  g386(.A1(new_n570), .A2(G110), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n397), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT22), .B(G137), .ZN(new_n575));
  AND2_X1   g389(.A1(G221), .A2(G234), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n189), .A2(new_n190), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(KEYINPUT77), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(KEYINPUT77), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n575), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n580), .ZN(new_n582));
  INV_X1    g396(.A(new_n575), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n582), .A2(new_n578), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n366), .A2(new_n386), .ZN(new_n586));
  OAI22_X1  g400(.A1(new_n570), .A2(G110), .B1(new_n571), .B2(new_n572), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n574), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n583), .B1(new_n582), .B2(new_n578), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n579), .A2(new_n580), .A3(new_n575), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n590), .A2(new_n591), .A3(KEYINPUT78), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT78), .B1(new_n590), .B2(new_n591), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n397), .A2(new_n573), .B1(new_n587), .B2(new_n586), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n589), .B(new_n300), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT25), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n574), .A2(new_n588), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n592), .B2(new_n593), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n600), .A2(KEYINPUT25), .A3(new_n300), .A4(new_n589), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n332), .B1(G234), .B2(new_n300), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(G902), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n604), .B(KEYINPUT79), .Z(new_n605));
  AND2_X1   g419(.A1(new_n600), .A2(new_n589), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n602), .A2(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT74), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n551), .B(new_n608), .C1(new_n563), .C2(new_n564), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n566), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n503), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(new_n231), .ZN(G3));
  NAND2_X1  g426(.A1(new_n559), .A2(new_n562), .ZN(new_n613));
  INV_X1    g427(.A(G472), .ZN(new_n614));
  AOI21_X1  g428(.A(G902), .B1(new_n553), .B2(new_n558), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n613), .B(new_n607), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n305), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT94), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n490), .A2(KEYINPUT95), .A3(new_n496), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT95), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n620), .B(new_n423), .C1(new_n488), .C2(new_n489), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n619), .A2(new_n500), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n347), .A2(KEYINPUT33), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n334), .A2(new_n341), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n624), .A2(G478), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n343), .A2(new_n300), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n350), .B2(new_n343), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n419), .A2(new_n358), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n618), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NOR2_X1   g450(.A1(new_n350), .A2(KEYINPUT93), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n345), .B1(new_n637), .B2(new_n342), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n351), .A2(new_n344), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n640), .A2(new_n359), .A3(new_n419), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n622), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n618), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT35), .B(G107), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  OR2_X1    g459(.A1(new_n615), .A2(new_n614), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n602), .A2(new_n603), .ZN(new_n647));
  INV_X1    g461(.A(new_n594), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n599), .B1(new_n648), .B2(KEYINPUT36), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT36), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n594), .A2(new_n650), .A3(new_n595), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n605), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n646), .A2(new_n613), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n421), .B(new_n656), .C1(new_n501), .C2(new_n502), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n355), .B1(new_n356), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n640), .A2(new_n654), .A3(new_n419), .A4(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n305), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n664), .A2(new_n566), .A3(new_n609), .A4(new_n623), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  INV_X1    g480(.A(new_n305), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n661), .B(KEYINPUT39), .Z(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n669), .A2(KEYINPUT40), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(KEYINPUT40), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n498), .B(KEYINPUT38), .ZN(new_n672));
  INV_X1    g486(.A(new_n520), .ZN(new_n673));
  AOI21_X1  g487(.A(G902), .B1(new_n673), .B2(new_n526), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n547), .A2(new_n525), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI22_X1  g490(.A1(new_n563), .A2(new_n564), .B1(new_n614), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n654), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n407), .A2(new_n415), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n418), .A2(G475), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n638), .A2(new_n639), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AND4_X1   g495(.A1(new_n500), .A2(new_n677), .A3(new_n678), .A4(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n670), .A2(new_n671), .A3(new_n672), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  NOR3_X1   g498(.A1(new_n419), .A2(new_n630), .A3(new_n661), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n654), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n305), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n687), .A2(new_n566), .A3(new_n609), .A4(new_n623), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  OAI21_X1  g503(.A(new_n293), .B1(new_n280), .B2(new_n281), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n194), .A2(new_n690), .B1(new_n291), .B2(new_n255), .ZN(new_n691));
  OAI21_X1  g505(.A(G469), .B1(new_n691), .B2(G902), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n188), .A3(new_n301), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n566), .A2(new_n607), .A3(new_n609), .A4(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n632), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT41), .B(G113), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  INV_X1    g512(.A(new_n642), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n314), .ZN(G18));
  NOR2_X1   g515(.A1(new_n622), .A2(new_n693), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n420), .A2(new_n678), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n566), .A2(new_n702), .A3(new_n703), .A4(new_n609), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  NAND4_X1  g519(.A1(new_n619), .A2(new_n681), .A3(new_n500), .A4(new_n621), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n692), .A2(new_n359), .A3(new_n188), .A4(new_n301), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n556), .A2(new_n557), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n521), .A2(new_n525), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n562), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n607), .B(new_n710), .C1(new_n615), .C2(new_n614), .ZN(new_n711));
  NOR4_X1   g525(.A1(new_n706), .A2(new_n707), .A3(new_n711), .A4(KEYINPUT96), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT96), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n707), .A2(new_n711), .ZN(new_n714));
  AND4_X1   g528(.A1(new_n500), .A2(new_n619), .A3(new_n681), .A4(new_n621), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT97), .B(G122), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G24));
  OAI211_X1 g533(.A(new_n654), .B(new_n710), .C1(new_n615), .C2(new_n614), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT98), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n685), .B(new_n702), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  NAND4_X1  g539(.A1(new_n492), .A2(new_n500), .A3(new_n496), .A4(new_n497), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT100), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n496), .A2(new_n500), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT100), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n492), .A3(new_n729), .A4(new_n497), .ZN(new_n730));
  INV_X1    g544(.A(new_n188), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n283), .A2(new_n285), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n194), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(G469), .A3(new_n294), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n302), .B(KEYINPUT99), .Z(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n690), .A2(new_n194), .ZN(new_n737));
  AOI21_X1  g551(.A(G902), .B1(new_n737), .B2(new_n297), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n736), .B1(new_n738), .B2(new_n287), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n731), .B1(new_n734), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n727), .A2(new_n730), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT101), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT101), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n727), .A2(new_n743), .A3(new_n740), .A4(new_n730), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n610), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n685), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n742), .A2(new_n744), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n565), .A2(new_n607), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n750), .A2(KEYINPUT42), .A3(new_n685), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n746), .A2(new_n747), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n208), .ZN(G33));
  AND3_X1   g567(.A1(new_n566), .A2(new_n607), .A3(new_n609), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n640), .A2(new_n419), .A3(new_n662), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n748), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  NAND3_X1  g572(.A1(new_n419), .A2(new_n627), .A3(new_n629), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT43), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n646), .A2(new_n613), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n654), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n727), .A2(new_n730), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n733), .A2(KEYINPUT45), .A3(new_n294), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n769), .B1(new_n286), .B2(new_n295), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(G469), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT46), .B1(new_n771), .B2(new_n735), .ZN(new_n772));
  INV_X1    g586(.A(new_n301), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n735), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n731), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n763), .A2(new_n764), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n767), .A2(new_n668), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(KEYINPUT103), .B(G137), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G39));
  OR2_X1    g594(.A1(new_n776), .A2(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n776), .A2(KEYINPUT47), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n566), .A2(new_n609), .ZN(new_n784));
  INV_X1    g598(.A(new_n607), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n766), .A3(new_n785), .A4(new_n685), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT104), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT104), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n783), .A2(new_n790), .A3(new_n787), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  NAND2_X1  g607(.A1(new_n692), .A2(new_n301), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT105), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT49), .Z(new_n796));
  INV_X1    g610(.A(new_n672), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n607), .A2(new_n500), .A3(new_n188), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n677), .A2(new_n759), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n761), .A2(new_n355), .ZN(new_n801));
  INV_X1    g615(.A(new_n711), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n766), .ZN(new_n805));
  INV_X1    g619(.A(new_n783), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n795), .A2(new_n188), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n672), .A2(new_n500), .A3(new_n693), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n804), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT50), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n766), .A2(new_n694), .ZN(new_n812));
  INV_X1    g626(.A(new_n355), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n677), .A2(new_n785), .A3(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n419), .A3(new_n630), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n812), .B(new_n801), .C1(new_n722), .C2(new_n723), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n808), .A2(new_n811), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n812), .A2(new_n750), .A3(new_n801), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT48), .ZN(new_n821));
  INV_X1    g635(.A(new_n702), .ZN(new_n822));
  OAI211_X1 g636(.A(G952), .B(new_n431), .C1(new_n803), .C2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n419), .A2(new_n630), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n823), .B1(new_n815), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT115), .B1(new_n821), .B2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n821), .A2(KEYINPUT115), .A3(new_n825), .ZN(new_n827));
  OAI22_X1  g641(.A1(new_n819), .A2(KEYINPUT51), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n810), .B(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT113), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(new_n831), .A3(new_n817), .A4(new_n816), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n832), .A2(KEYINPUT51), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n834));
  INV_X1    g648(.A(new_n808), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT113), .B1(new_n811), .B2(new_n818), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n833), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n832), .A3(KEYINPUT51), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT114), .B1(new_n838), .B2(new_n808), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n828), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n665), .A2(new_n724), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n654), .A2(new_n661), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n740), .A2(KEYINPUT109), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n301), .A2(new_n735), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n188), .B(new_n842), .C1(new_n296), .C2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT109), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n843), .A2(new_n847), .A3(new_n677), .A4(new_n715), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n841), .A2(KEYINPUT52), .A3(new_n688), .A4(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(KEYINPUT110), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n848), .A2(new_n665), .A3(new_n688), .A4(new_n724), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n850), .B1(new_n854), .B2(KEYINPUT110), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n419), .A2(new_n353), .A3(new_n654), .A4(new_n662), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n667), .A2(new_n727), .A3(new_n730), .A4(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n784), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n745), .B2(new_n756), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT108), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n685), .B1(new_n722), .B2(new_n723), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n861), .B1(new_n748), .B2(new_n863), .ZN(new_n864));
  AOI211_X1 g678(.A(KEYINPUT108), .B(new_n862), .C1(new_n742), .C2(new_n744), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n752), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n754), .A2(new_n633), .A3(new_n694), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n754), .A2(new_n642), .A3(new_n694), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n868), .A2(new_n869), .A3(new_n717), .A4(new_n704), .ZN(new_n870));
  INV_X1    g684(.A(new_n617), .ZN(new_n871));
  INV_X1    g685(.A(new_n641), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(new_n501), .B2(new_n502), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT107), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT107), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n875), .B(new_n872), .C1(new_n501), .C2(new_n502), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n871), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n824), .A2(KEYINPUT106), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT106), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n879), .B1(new_n419), .B2(new_n630), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(new_n358), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n882), .B(new_n617), .C1(new_n501), .C2(new_n502), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n883), .B(new_n657), .C1(new_n610), .C2(new_n503), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n870), .A2(new_n877), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n855), .A2(new_n856), .A3(new_n867), .A4(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n866), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n746), .A2(new_n747), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n748), .A2(new_n751), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n849), .A2(new_n853), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n887), .A2(new_n885), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT53), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n886), .A2(new_n893), .A3(KEYINPUT54), .ZN(new_n894));
  XNOR2_X1  g708(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n704), .B1(new_n712), .B2(new_n716), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n696), .A2(new_n897), .A3(new_n700), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n874), .A2(new_n876), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n617), .ZN(new_n900));
  INV_X1    g714(.A(new_n884), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n898), .A2(KEYINPUT53), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n902), .A2(new_n866), .A3(new_n752), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n896), .B1(new_n903), .B2(new_n855), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n892), .A2(new_n856), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n894), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT112), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT112), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n894), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n840), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT116), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n354), .A2(new_n431), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n911), .A2(KEYINPUT116), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n800), .B1(new_n914), .B2(new_n915), .ZN(G75));
  INV_X1    g730(.A(KEYINPUT56), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n903), .A2(new_n855), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n905), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(G902), .ZN(new_n920));
  INV_X1    g734(.A(G210), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n483), .A2(new_n485), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(new_n486), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT55), .Z(new_n925));
  XNOR2_X1  g739(.A(new_n922), .B(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n191), .A2(G952), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT117), .Z(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n926), .A2(new_n929), .ZN(G51));
  AOI22_X1  g744(.A1(new_n856), .A2(new_n892), .B1(new_n903), .B2(new_n855), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT119), .B1(new_n931), .B2(new_n895), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n919), .A2(new_n933), .A3(new_n896), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT118), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n904), .A2(new_n935), .A3(new_n905), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n935), .B1(new_n904), .B2(new_n905), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n932), .B(new_n934), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n735), .B(KEYINPUT57), .Z(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT120), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n938), .A2(KEYINPUT120), .A3(new_n939), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n299), .A3(new_n943), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n920), .A2(new_n771), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n927), .B1(new_n944), .B2(new_n945), .ZN(G54));
  AND4_X1   g760(.A1(KEYINPUT58), .A2(new_n919), .A3(G475), .A4(G902), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n947), .A2(new_n413), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n947), .A2(new_n413), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n948), .A2(new_n949), .A3(new_n927), .ZN(G60));
  AND2_X1   g764(.A1(new_n624), .A2(new_n626), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n908), .A2(new_n910), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n628), .B(KEYINPUT59), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n951), .A2(new_n953), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n929), .B1(new_n938), .B2(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n954), .A2(new_n956), .ZN(G63));
  INV_X1    g771(.A(KEYINPUT60), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n958), .A2(G217), .A3(G902), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(G217), .B2(G902), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n931), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n652), .ZN(new_n962));
  NOR2_X1   g776(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n929), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n962), .B(new_n964), .C1(new_n606), .C2(new_n961), .ZN(new_n965));
  NAND2_X1  g779(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(G66));
  INV_X1    g781(.A(G224), .ZN(new_n968));
  OAI21_X1  g782(.A(G953), .B1(new_n357), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n191), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n969), .B1(new_n885), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n923), .B1(G898), .B2(new_n191), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT122), .Z(new_n973));
  XNOR2_X1  g787(.A(new_n971), .B(new_n973), .ZN(G69));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n776), .A2(new_n668), .A3(new_n715), .A4(new_n750), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n841), .A2(new_n688), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n778), .A2(new_n757), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n978), .A2(new_n752), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n792), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n792), .A2(new_n982), .A3(new_n979), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n981), .A2(new_n191), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n544), .A2(new_n545), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n370), .A2(new_n371), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n985), .B(new_n986), .Z(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n660), .B2(new_n191), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n975), .B1(new_n984), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n977), .A2(new_n683), .ZN(new_n993));
  OR3_X1    g807(.A1(new_n993), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n994));
  OAI21_X1  g808(.A(KEYINPUT124), .B1(new_n993), .B2(KEYINPUT62), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n640), .A2(new_n419), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n669), .B1(new_n997), .B2(new_n881), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n998), .A2(new_n754), .A3(new_n766), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n778), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(KEYINPUT62), .B2(new_n993), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n996), .A2(new_n792), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n191), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n987), .B(KEYINPUT123), .Z(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  AOI22_X1  g820(.A1(new_n1006), .A2(KEYINPUT125), .B1(new_n984), .B2(new_n989), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT125), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1003), .A2(new_n1008), .A3(new_n1005), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n992), .B(new_n1010), .ZN(G72));
  NAND3_X1  g825(.A1(new_n981), .A2(new_n885), .A3(new_n983), .ZN(new_n1012));
  NAND2_X1  g826(.A1(G472), .A2(G902), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT63), .Z(new_n1014));
  AOI211_X1 g828(.A(new_n525), .B(new_n547), .C1(new_n1012), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n885), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n1002), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n675), .B1(new_n1017), .B2(new_n1014), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n548), .A2(new_n554), .ZN(new_n1019));
  AND4_X1   g833(.A1(new_n893), .A2(new_n886), .A3(new_n1014), .A4(new_n1019), .ZN(new_n1020));
  NOR4_X1   g834(.A1(new_n1015), .A2(new_n1018), .A3(new_n927), .A4(new_n1020), .ZN(G57));
endmodule


