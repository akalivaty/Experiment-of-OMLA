//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G43gat), .ZN(new_n203));
  INV_X1    g002(.A(G43gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G50gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT15), .ZN(new_n206));
  NAND2_X1  g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT82), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(new_n202), .B2(G43gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(new_n203), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n205), .A2(new_n210), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(KEYINPUT83), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(KEYINPUT83), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n208), .B(new_n214), .C1(new_n219), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n218), .A2(new_n221), .B1(G29gat), .B2(G36gat), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n224), .A2(new_n206), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G8gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(G15gat), .B(G22gat), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n228), .A2(G1gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT16), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n228), .B1(new_n230), .B2(G1gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n227), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n227), .A3(new_n231), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n226), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G229gat), .A2(G233gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT18), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT85), .B1(new_n234), .B2(new_n232), .ZN(new_n240));
  INV_X1    g039(.A(new_n232), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT85), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n242), .A3(new_n233), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT17), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n240), .B(new_n243), .C1(new_n244), .C2(new_n226), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT84), .B(KEYINPUT17), .Z(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n226), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n235), .B(new_n239), .C1(new_n245), .C2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT86), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n223), .A2(new_n225), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n234), .A2(new_n232), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(new_n235), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n236), .B(KEYINPUT13), .Z(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n253), .A2(KEYINPUT17), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n259), .A2(new_n248), .A3(new_n243), .A4(new_n240), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n260), .A2(KEYINPUT86), .A3(new_n235), .A4(new_n239), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n252), .A2(new_n258), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT87), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n260), .A2(new_n235), .A3(new_n236), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n238), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n252), .A2(KEYINPUT87), .A3(new_n258), .A4(new_n261), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G113gat), .B(G141gat), .ZN(new_n269));
  INV_X1    g068(.A(G197gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT11), .B(G169gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n273), .B(KEYINPUT12), .Z(new_n274));
  INV_X1    g073(.A(KEYINPUT88), .ZN(new_n275));
  INV_X1    g074(.A(new_n274), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n266), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n275), .B1(new_n277), .B2(new_n262), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n261), .A2(new_n258), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n274), .B1(new_n265), .B2(new_n238), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT88), .A4(new_n252), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n268), .A2(new_n274), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g081(.A1(G232gat), .A2(G233gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(KEYINPUT41), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT92), .ZN(new_n285));
  NAND2_X1  g084(.A1(G85gat), .A2(G92gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT7), .ZN(new_n287));
  NAND2_X1  g086(.A1(G99gat), .A2(G106gat), .ZN(new_n288));
  INV_X1    g087(.A(G85gat), .ZN(new_n289));
  INV_X1    g088(.A(G92gat), .ZN(new_n290));
  AOI22_X1  g089(.A1(KEYINPUT8), .A2(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G99gat), .B(G106gat), .Z(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n293), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(new_n287), .A3(new_n291), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n226), .A2(new_n297), .B1(KEYINPUT41), .B2(new_n283), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n296), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(new_n226), .B2(new_n244), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n249), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT93), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G190gat), .B(G218gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(new_n301), .B2(new_n302), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n285), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n301), .A2(new_n302), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n303), .B1(new_n308), .B2(new_n305), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n284), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n303), .A3(new_n305), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n304), .A2(new_n306), .ZN(new_n312));
  INV_X1    g111(.A(new_n284), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n285), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G134gat), .B(G162gat), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n310), .A2(new_n316), .A3(new_n314), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G57gat), .B(G64gat), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n321), .A2(KEYINPUT90), .ZN(new_n322));
  NAND2_X1  g121(.A1(G71gat), .A2(G78gat), .ZN(new_n323));
  INV_X1    g122(.A(G71gat), .ZN(new_n324));
  INV_X1    g123(.A(G78gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT9), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n321), .A2(KEYINPUT90), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(G71gat), .B(G78gat), .Z(new_n329));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n329), .B1(new_n330), .B2(new_n321), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT89), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G57gat), .B(G64gat), .Z(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT9), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT89), .B1(new_n335), .B2(new_n329), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n328), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT21), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G231gat), .A2(G233gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(G127gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(G183gat), .B(G211gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n254), .B1(new_n337), .B2(new_n338), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(KEYINPUT91), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n347));
  INV_X1    g146(.A(G155gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n346), .B(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n344), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT10), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n332), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n335), .A2(KEYINPUT89), .A3(new_n329), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n353), .A2(new_n354), .B1(new_n322), .B2(new_n327), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n296), .A2(KEYINPUT94), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n299), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n299), .B1(new_n355), .B2(new_n356), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n352), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n337), .A2(new_n299), .A3(new_n352), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(KEYINPUT95), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT95), .ZN(new_n364));
  INV_X1    g163(.A(new_n356), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n297), .B1(new_n337), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT10), .B1(new_n366), .B2(new_n357), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n364), .B1(new_n367), .B2(new_n361), .ZN(new_n368));
  NAND2_X1  g167(.A1(G230gat), .A2(G233gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n363), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n358), .A2(new_n359), .A3(new_n369), .ZN(new_n371));
  XOR2_X1   g170(.A(G120gat), .B(G148gat), .Z(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT96), .ZN(new_n373));
  XOR2_X1   g172(.A(G176gat), .B(G204gat), .Z(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n371), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n367), .A2(new_n361), .ZN(new_n380));
  INV_X1    g179(.A(new_n369), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n382), .A2(KEYINPUT97), .A3(new_n376), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT97), .B1(new_n382), .B2(new_n376), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n378), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n320), .A2(new_n351), .A3(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT23), .ZN(new_n389));
  NAND2_X1  g188(.A1(G169gat), .A2(G176gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT23), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(G169gat), .B2(G176gat), .ZN(new_n392));
  OR2_X1    g191(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n389), .A2(new_n390), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G183gat), .A2(G190gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT24), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n397), .B(new_n398), .C1(G183gat), .C2(G190gat), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n394), .B(new_n399), .C1(new_n400), .C2(KEYINPUT64), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT26), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n390), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(new_n388), .ZN(new_n404));
  INV_X1    g203(.A(G169gat), .ZN(new_n405));
  INV_X1    g204(.A(G176gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT26), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n395), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT27), .B(G183gat), .ZN(new_n410));
  INV_X1    g209(.A(G190gat), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT28), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G183gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT27), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT27), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G183gat), .ZN(new_n416));
  AND4_X1   g215(.A1(KEYINPUT28), .A2(new_n414), .A3(new_n416), .A4(new_n411), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n409), .B1(new_n412), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT25), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n395), .A2(KEYINPUT65), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT65), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n422), .A2(G183gat), .A3(G190gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n423), .A3(new_n396), .ZN(new_n424));
  AND3_X1   g223(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n413), .A2(new_n411), .A3(KEYINPUT66), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT66), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(G183gat), .B2(G190gat), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n425), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n420), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n401), .B(new_n418), .C1(new_n419), .C2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT29), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(G226gat), .A2(G233gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n429), .A2(new_n424), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n400), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n414), .A2(new_n416), .A3(new_n411), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT28), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n410), .A2(KEYINPUT28), .A3(new_n411), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n437), .A2(KEYINPUT25), .B1(new_n442), .B2(new_n409), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n434), .B1(new_n443), .B2(new_n401), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  XOR2_X1   g244(.A(G211gat), .B(G218gat), .Z(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(G211gat), .A2(G218gat), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT22), .ZN(new_n449));
  OR2_X1    g248(.A1(G197gat), .A2(G204gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(G197gat), .A2(G204gat), .ZN(new_n451));
  AOI221_X4 g250(.A(KEYINPUT70), .B1(new_n448), .B2(new_n449), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT70), .ZN(new_n453));
  XNOR2_X1  g252(.A(G197gat), .B(G204gat), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n447), .B1(new_n452), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n454), .A2(new_n453), .A3(new_n456), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n446), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n435), .A2(new_n445), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n461), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n431), .A2(new_n432), .B1(G226gat), .B2(G233gat), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(new_n444), .ZN(new_n465));
  XNOR2_X1  g264(.A(G8gat), .B(G36gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT71), .ZN(new_n467));
  XNOR2_X1  g266(.A(G64gat), .B(G92gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n467), .B(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n462), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT30), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n469), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n461), .B1(new_n435), .B2(new_n445), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n464), .A2(new_n444), .A3(new_n463), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n462), .A2(new_n465), .A3(KEYINPUT30), .A4(new_n469), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n473), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(G1gat), .B(G29gat), .Z(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G57gat), .B(G85gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  XOR2_X1   g284(.A(KEYINPUT76), .B(KEYINPUT5), .Z(new_n486));
  AND2_X1   g285(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n487));
  NOR2_X1   g286(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n488));
  OAI21_X1  g287(.A(G127gat), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G113gat), .ZN(new_n490));
  INV_X1    g289(.A(G120gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT1), .ZN(new_n493));
  NAND2_X1  g292(.A1(G113gat), .A2(G120gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OR2_X1    g294(.A1(G127gat), .A2(G134gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n489), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT1), .B1(new_n490), .B2(new_n491), .ZN(new_n498));
  XNOR2_X1  g297(.A(G127gat), .B(G134gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT68), .B(G113gat), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n498), .B(new_n499), .C1(new_n500), .C2(new_n491), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT75), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT73), .ZN(new_n505));
  AND2_X1   g304(.A1(G141gat), .A2(G148gat), .ZN(new_n506));
  NOR2_X1   g305(.A1(G141gat), .A2(G148gat), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G141gat), .ZN(new_n509));
  INV_X1    g308(.A(G148gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G141gat), .A2(G148gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(KEYINPUT73), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT2), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n508), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G155gat), .B(G162gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n506), .A2(new_n507), .ZN(new_n519));
  NAND2_X1  g318(.A1(G155gat), .A2(G162gat), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n520), .A2(KEYINPUT74), .A3(KEYINPUT2), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT74), .B1(new_n520), .B2(KEYINPUT2), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n516), .B(new_n519), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n497), .A2(new_n501), .A3(KEYINPUT75), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n504), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n502), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(new_n518), .A3(new_n523), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G225gat), .A2(G233gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n486), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT4), .B1(new_n524), .B2(new_n502), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT4), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n527), .A2(new_n534), .A3(new_n518), .A4(new_n523), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n524), .A2(KEYINPUT3), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT3), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n518), .A2(new_n538), .A3(new_n523), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n537), .A2(new_n504), .A3(new_n525), .A4(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(new_n540), .A3(new_n530), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n532), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT78), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n533), .A2(new_n535), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n528), .A2(KEYINPUT78), .A3(KEYINPUT4), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n540), .A2(new_n530), .A3(new_n486), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n485), .B1(new_n542), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT6), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n541), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n551), .B(new_n484), .C1(new_n546), .C2(new_n547), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(KEYINPUT6), .B(new_n485), .C1(new_n542), .C2(new_n548), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(KEYINPUT80), .B(KEYINPUT35), .Z(new_n556));
  NAND3_X1  g355(.A1(new_n479), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT34), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n431), .A2(new_n527), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n437), .A2(KEYINPUT25), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n560), .A2(new_n502), .A3(new_n401), .A4(new_n418), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G227gat), .A2(G233gat), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n558), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n563), .ZN(new_n565));
  AOI211_X1 g364(.A(KEYINPUT34), .B(new_n565), .C1(new_n559), .C2(new_n561), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n559), .A2(new_n565), .A3(new_n561), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT33), .ZN(new_n569));
  XNOR2_X1  g368(.A(G15gat), .B(G43gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(G71gat), .B(G99gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n568), .B(KEYINPUT32), .C1(new_n569), .C2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n572), .B1(new_n568), .B2(KEYINPUT32), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n568), .A2(KEYINPUT69), .A3(new_n569), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT69), .B1(new_n568), .B2(new_n569), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n567), .B(new_n573), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n568), .A2(new_n569), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT69), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n575), .A3(new_n574), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n567), .B1(new_n583), .B2(new_n573), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G228gat), .A2(G233gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G78gat), .B(G106gat), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n518), .A2(new_n523), .ZN(new_n589));
  AND2_X1   g388(.A1(G197gat), .A2(G204gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(G197gat), .A2(G204gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT70), .B1(new_n592), .B2(new_n455), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n446), .B1(new_n593), .B2(new_n459), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n452), .A2(new_n447), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n432), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n589), .B1(new_n596), .B2(new_n538), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n461), .B1(new_n432), .B2(new_n539), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n588), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT31), .B(G50gat), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT29), .B1(new_n458), .B2(new_n460), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n524), .B1(new_n601), .B2(KEYINPUT3), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n539), .A2(new_n432), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(new_n463), .ZN(new_n604));
  INV_X1    g403(.A(new_n588), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n599), .A2(new_n600), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n600), .B1(new_n599), .B2(new_n606), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n587), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT79), .B(G22gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n600), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n597), .A2(new_n598), .A3(new_n588), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n605), .B1(new_n602), .B2(new_n604), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n599), .A2(new_n606), .A3(new_n600), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(new_n586), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n609), .A2(new_n610), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n610), .B1(new_n609), .B2(new_n616), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n585), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n557), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n610), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n607), .A2(new_n608), .A3(new_n587), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n586), .B1(new_n614), .B2(new_n615), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n617), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n472), .B1(new_n553), .B2(new_n554), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT72), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n477), .A2(new_n629), .A3(new_n478), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n477), .B2(new_n478), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n627), .A2(new_n628), .A3(new_n585), .A4(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT81), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n633), .A2(new_n634), .A3(KEYINPUT35), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n634), .B1(new_n633), .B2(KEYINPUT35), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n622), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n544), .A2(new_n540), .A3(new_n545), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n531), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n639), .A2(KEYINPUT39), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n639), .B(KEYINPUT39), .C1(new_n531), .C2(new_n529), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n641), .A3(new_n484), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n473), .A2(new_n477), .A3(new_n478), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n644), .A2(new_n549), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n475), .A2(new_n476), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT37), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n648), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT37), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n474), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT38), .ZN(new_n654));
  INV_X1    g453(.A(new_n555), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n470), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n627), .B(new_n647), .C1(new_n654), .C2(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n585), .A2(KEYINPUT36), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n585), .A2(KEYINPUT36), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n627), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n555), .A2(new_n632), .A3(new_n473), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n657), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  AOI211_X1 g463(.A(new_n282), .B(new_n387), .C1(new_n637), .C2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n655), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g466(.A(KEYINPUT16), .B(G8gat), .Z(new_n668));
  AND3_X1   g467(.A1(new_n665), .A2(new_n645), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n227), .B1(new_n665), .B2(new_n645), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT42), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n671), .B1(KEYINPUT42), .B2(new_n669), .ZN(G1325gat));
  INV_X1    g471(.A(G15gat), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n665), .A2(new_n673), .A3(new_n585), .ZN(new_n674));
  INV_X1    g473(.A(new_n660), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n665), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n674), .B1(new_n676), .B2(new_n673), .ZN(G1326gat));
  NAND2_X1  g476(.A1(new_n665), .A2(new_n661), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT43), .B(G22gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  NOR3_X1   g479(.A1(new_n351), .A2(new_n282), .A3(new_n385), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT98), .Z(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT35), .B1(new_n620), .B2(new_n662), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT81), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n633), .A2(new_n634), .A3(KEYINPUT35), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT99), .B1(new_n687), .B2(new_n622), .ZN(new_n688));
  OAI211_X1 g487(.A(KEYINPUT99), .B(new_n622), .C1(new_n635), .C2(new_n636), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n664), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n318), .A2(new_n319), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n320), .B1(new_n637), .B2(new_n664), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n692), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n683), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(G29gat), .B1(new_n699), .B2(new_n555), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n695), .A2(new_n681), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n216), .A3(new_n655), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(G1328gat));
  AOI21_X1  g503(.A(new_n217), .B1(new_n698), .B2(new_n645), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n695), .A2(new_n681), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n645), .A2(new_n217), .ZN(new_n707));
  OR3_X1    g506(.A1(new_n706), .A2(KEYINPUT46), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT46), .B1(new_n706), .B2(new_n707), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OR3_X1    g509(.A1(new_n705), .A2(KEYINPUT100), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT100), .B1(new_n705), .B2(new_n710), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(G1329gat));
  INV_X1    g512(.A(new_n585), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n204), .B1(new_n706), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n675), .A2(G43gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(new_n699), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g517(.A(KEYINPUT48), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n693), .A2(new_n692), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT99), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n637), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n689), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n720), .B1(new_n723), .B2(new_n664), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n661), .B(new_n682), .C1(new_n724), .C2(new_n696), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G50gat), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n627), .A2(G50gat), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n706), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n719), .B1(new_n726), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT101), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n701), .A2(new_n732), .A3(new_n727), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT101), .B1(new_n706), .B2(new_n728), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(new_n719), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n735), .B1(G50gat), .B2(new_n725), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT102), .B1(new_n731), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT48), .B1(new_n729), .B2(new_n732), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n726), .A2(new_n734), .A3(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT102), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n729), .B1(new_n725), .B2(G50gat), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n739), .B(new_n740), .C1(new_n719), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n737), .A2(new_n742), .ZN(G1331gat));
  INV_X1    g542(.A(new_n664), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n722), .B2(new_n689), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n320), .A2(new_n282), .A3(new_n351), .A4(new_n385), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n655), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g548(.A1(new_n745), .A2(new_n479), .A3(new_n746), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  AND2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n750), .B2(new_n751), .ZN(G1333gat));
  AOI21_X1  g553(.A(new_n324), .B1(new_n747), .B2(new_n675), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n714), .A2(G71gat), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n747), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g557(.A1(new_n747), .A2(new_n661), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G78gat), .ZN(G1335gat));
  INV_X1    g559(.A(new_n351), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(new_n282), .A3(new_n693), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n691), .A2(KEYINPUT51), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n745), .B2(new_n762), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n386), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n767), .A2(new_n289), .A3(new_n655), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n761), .A2(new_n282), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n386), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n694), .B2(new_n697), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n772), .A2(new_n655), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n768), .B1(new_n773), .B2(new_n289), .ZN(G1336gat));
  OAI211_X1 g573(.A(new_n645), .B(new_n770), .C1(new_n724), .C2(new_n696), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n775), .A2(KEYINPUT103), .A3(G92gat), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT103), .B1(new_n775), .B2(G92gat), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n385), .A2(new_n290), .A3(new_n645), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT104), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n764), .B2(new_n766), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n776), .A2(new_n777), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n764), .A2(new_n766), .ZN(new_n783));
  INV_X1    g582(.A(new_n779), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT52), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n775), .A2(G92gat), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n785), .A2(KEYINPUT105), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT105), .B1(new_n785), .B2(new_n786), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n781), .A2(new_n782), .B1(new_n787), .B2(new_n788), .ZN(G1337gat));
  INV_X1    g588(.A(G99gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n675), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n791), .B2(KEYINPUT106), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(KEYINPUT106), .B2(new_n791), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n767), .A2(new_n790), .A3(new_n585), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(G1338gat));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n627), .A2(G106gat), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n783), .A2(new_n385), .A3(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n661), .B(new_n770), .C1(new_n724), .C2(new_n696), .ZN(new_n799));
  XOR2_X1   g598(.A(KEYINPUT107), .B(G106gat), .Z(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g600(.A(KEYINPUT108), .B(KEYINPUT53), .ZN(new_n802));
  AND4_X1   g601(.A1(new_n796), .A2(new_n798), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n767), .A2(new_n797), .B1(new_n799), .B2(new_n800), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n796), .B1(new_n804), .B2(new_n802), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n798), .A2(new_n801), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT53), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n803), .B1(new_n805), .B2(new_n807), .ZN(G1339gat));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n278), .A2(new_n281), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n236), .B1(new_n260), .B2(new_n235), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI22_X1  g613(.A1(new_n811), .A2(KEYINPUT111), .B1(new_n256), .B2(new_n257), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n273), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n385), .A2(new_n810), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n380), .B2(new_n381), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n370), .A2(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n818), .B(new_n369), .C1(new_n367), .C2(new_n361), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n821), .A2(KEYINPUT110), .A3(new_n376), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT110), .B1(new_n821), .B2(new_n376), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n820), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n820), .B(KEYINPUT55), .C1(new_n822), .C2(new_n823), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n378), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n817), .B1(new_n828), .B2(new_n282), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n320), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n810), .A2(new_n816), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n318), .B2(new_n319), .ZN(new_n832));
  INV_X1    g631(.A(new_n828), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n351), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n320), .A2(new_n351), .A3(new_n386), .A4(new_n282), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n809), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n829), .A2(new_n320), .B1(new_n832), .B2(new_n833), .ZN(new_n839));
  OAI211_X1 g638(.A(KEYINPUT112), .B(new_n836), .C1(new_n839), .C2(new_n351), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n620), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n645), .A2(new_n555), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G113gat), .B1(new_n843), .B2(new_n282), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n841), .A2(new_n845), .A3(new_n842), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n845), .B1(new_n841), .B2(new_n842), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n282), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n500), .ZN(new_n851));
  XOR2_X1   g650(.A(new_n851), .B(KEYINPUT114), .Z(new_n852));
  OAI21_X1  g651(.A(new_n844), .B1(new_n849), .B2(new_n852), .ZN(G1340gat));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n385), .A2(new_n491), .ZN(new_n855));
  INV_X1    g654(.A(new_n848), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n846), .ZN(new_n857));
  OAI21_X1  g656(.A(G120gat), .B1(new_n843), .B2(new_n386), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n854), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  OAI211_X1 g659(.A(KEYINPUT115), .B(new_n858), .C1(new_n849), .C2(new_n855), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1341gat));
  NOR2_X1   g661(.A1(new_n843), .A2(new_n761), .ZN(new_n863));
  XNOR2_X1  g662(.A(KEYINPUT116), .B(G127gat), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n863), .B(new_n864), .ZN(G1342gat));
  NOR2_X1   g664(.A1(new_n320), .A2(new_n645), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n555), .A2(new_n488), .A3(new_n487), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n841), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n868), .B(KEYINPUT56), .Z(new_n869));
  OAI21_X1  g668(.A(G134gat), .B1(new_n843), .B2(new_n320), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1343gat));
  NAND2_X1  g670(.A1(new_n838), .A2(new_n840), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n873), .A3(new_n661), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n660), .A2(new_n842), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n836), .B1(new_n839), .B2(new_n351), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n661), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n877), .B2(KEYINPUT57), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G141gat), .B1(new_n879), .B2(new_n282), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n555), .B1(new_n838), .B2(new_n840), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(KEYINPUT118), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n675), .A2(new_n627), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n881), .B2(KEYINPUT118), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n282), .A2(G141gat), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n882), .A2(new_n885), .A3(new_n479), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n880), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n890), .A3(KEYINPUT58), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT58), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n880), .B(new_n887), .C1(new_n889), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(G1344gat));
  NAND2_X1  g693(.A1(new_n882), .A2(new_n885), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n645), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n510), .A3(new_n385), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n879), .A2(new_n386), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(KEYINPUT59), .A3(new_n510), .ZN(new_n899));
  XOR2_X1   g698(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n900));
  NOR2_X1   g699(.A1(new_n875), .A2(new_n386), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n873), .B(new_n627), .C1(new_n838), .C2(new_n840), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n877), .A2(new_n873), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n901), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n900), .B1(new_n905), .B2(G148gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n897), .B1(new_n899), .B2(new_n906), .ZN(G1345gat));
  NAND3_X1  g706(.A1(new_n896), .A2(new_n348), .A3(new_n351), .ZN(new_n908));
  OAI21_X1  g707(.A(G155gat), .B1(new_n879), .B2(new_n761), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1346gat));
  OAI21_X1  g709(.A(G162gat), .B1(new_n879), .B2(new_n320), .ZN(new_n911));
  INV_X1    g710(.A(G162gat), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n866), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n911), .B1(new_n895), .B2(new_n913), .ZN(G1347gat));
  NOR2_X1   g713(.A1(new_n655), .A2(new_n479), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n841), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n916), .A2(new_n282), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(new_n405), .ZN(G1348gat));
  OAI21_X1  g717(.A(new_n385), .B1(KEYINPUT120), .B2(G176gat), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(KEYINPUT120), .A2(G176gat), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n920), .B(new_n921), .ZN(G1349gat));
  OR3_X1    g721(.A1(new_n916), .A2(new_n410), .A3(new_n761), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n413), .B1(new_n916), .B2(new_n761), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n924), .B1(new_n923), .B2(new_n925), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(G1350gat));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n916), .A2(new_n320), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n929), .B(new_n930), .C1(new_n931), .C2(new_n411), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n411), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n411), .B1(KEYINPUT121), .B2(KEYINPUT61), .ZN(new_n934));
  OAI221_X1 g733(.A(new_n934), .B1(KEYINPUT121), .B2(KEYINPUT61), .C1(new_n916), .C2(new_n320), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(G1351gat));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n937), .B1(new_n902), .B2(new_n904), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n660), .A2(new_n915), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT125), .Z(new_n940));
  NAND3_X1  g739(.A1(new_n872), .A2(KEYINPUT57), .A3(new_n661), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n941), .A2(KEYINPUT124), .A3(new_n903), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n938), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n943), .A2(new_n270), .A3(new_n282), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n660), .A2(new_n661), .A3(new_n645), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n947), .A2(new_n948), .A3(new_n655), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n872), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n950), .B(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(G197gat), .B1(new_n952), .B2(new_n850), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n944), .A2(new_n953), .ZN(G1352gat));
  OAI21_X1  g753(.A(G204gat), .B1(new_n943), .B2(new_n386), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n950), .A2(G204gat), .A3(new_n386), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT62), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1353gat));
  INV_X1    g757(.A(G211gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n952), .A2(new_n959), .A3(new_n351), .ZN(new_n960));
  NOR2_X1   g759(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n940), .A2(new_n351), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n962), .B1(new_n941), .B2(new_n903), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n961), .B1(new_n963), .B2(new_n959), .ZN(new_n964));
  NAND2_X1  g763(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n963), .A2(new_n959), .A3(new_n961), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n960), .B1(new_n966), .B2(new_n967), .ZN(G1354gat));
  AOI21_X1  g767(.A(G218gat), .B1(new_n952), .B2(new_n693), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n693), .A2(G218gat), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n970), .B1(new_n943), .B2(KEYINPUT127), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n938), .A2(new_n972), .A3(new_n942), .A4(new_n940), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n969), .B1(new_n971), .B2(new_n973), .ZN(G1355gat));
endmodule


