//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n844, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202));
  INV_X1    g001(.A(G228gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT72), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n211));
  INV_X1    g010(.A(G197gat), .ZN(new_n212));
  INV_X1    g011(.A(G204gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G197gat), .A2(G204gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n211), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n210), .B(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n207), .B1(new_n217), .B2(KEYINPUT29), .ZN(new_n218));
  XOR2_X1   g017(.A(G155gat), .B(G162gat), .Z(new_n219));
  XNOR2_X1  g018(.A(G141gat), .B(G148gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(KEYINPUT2), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G155gat), .ZN(new_n222));
  INV_X1    g021(.A(G162gat), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT2), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n219), .B1(KEYINPUT77), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(KEYINPUT77), .B2(new_n224), .ZN(new_n226));
  INV_X1    g025(.A(G148gat), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n227), .A2(G141gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT76), .B(G141gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(G148gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n221), .B1(new_n226), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n206), .B1(new_n218), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT81), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n207), .B(new_n221), .C1(new_n226), .C2(new_n230), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n217), .B1(new_n235), .B2(KEYINPUT29), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n232), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n233), .B1(new_n232), .B2(new_n236), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT80), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n236), .A2(new_n240), .B1(new_n231), .B2(new_n218), .ZN(new_n241));
  INV_X1    g040(.A(new_n217), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT29), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n242), .B1(new_n234), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT80), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n205), .B1(new_n241), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(G22gat), .B1(new_n239), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n245), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n218), .A2(new_n231), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(new_n244), .B2(KEYINPUT80), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n206), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G22gat), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n251), .B(new_n252), .C1(new_n238), .C2(new_n237), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n202), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G78gat), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n255), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT31), .B(G50gat), .ZN(new_n258));
  INV_X1    g057(.A(G106gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n256), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n260), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n254), .A2(new_n255), .ZN(new_n263));
  AOI211_X1 g062(.A(new_n202), .B(G78gat), .C1(new_n247), .C2(new_n253), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT24), .ZN(new_n267));
  XOR2_X1   g066(.A(KEYINPUT66), .B(G190gat), .Z(new_n268));
  OAI21_X1  g067(.A(new_n267), .B1(G183gat), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G169gat), .ZN(new_n270));
  INV_X1    g069(.A(G176gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n271), .A3(KEYINPUT23), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT23), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(G169gat), .B2(G176gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n269), .A2(KEYINPUT25), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n276), .B(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n267), .B1(G183gat), .B2(G190gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT64), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n267), .B(KEYINPUT64), .C1(G183gat), .C2(G190gat), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n280), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n278), .B1(new_n285), .B2(KEYINPUT25), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT27), .B(G183gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(new_n268), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(KEYINPUT28), .ZN(new_n290));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT26), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n275), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(new_n293), .A3(new_n266), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n286), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G226gat), .A2(G233gat), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n242), .B(new_n297), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n295), .A2(new_n301), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n303), .B1(new_n300), .B2(new_n296), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n302), .B1(new_n304), .B2(new_n242), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT37), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n217), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n242), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT37), .ZN(new_n311));
  XNOR2_X1  g110(.A(G8gat), .B(G36gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(G64gat), .B(G92gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n314), .B(KEYINPUT73), .Z(new_n315));
  INV_X1    g114(.A(KEYINPUT38), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n307), .A2(new_n311), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT6), .ZN(new_n319));
  OR2_X1    g118(.A1(new_n226), .A2(new_n230), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT4), .ZN(new_n321));
  XOR2_X1   g120(.A(G127gat), .B(G134gat), .Z(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G113gat), .ZN(new_n324));
  INV_X1    g123(.A(G120gat), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT1), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT68), .B(G120gat), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n323), .B(new_n326), .C1(new_n324), .C2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n324), .B2(new_n325), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n322), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n320), .A2(new_n321), .A3(new_n221), .A4(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT4), .B1(new_n231), .B2(new_n331), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G225gat), .A2(G233gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(KEYINPUT78), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n231), .A2(KEYINPUT3), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(new_n331), .A3(new_n234), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT5), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n231), .B(new_n331), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n337), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n342), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G1gat), .B(G29gat), .ZN(new_n348));
  INV_X1    g147(.A(G85gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT0), .B(G57gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  OR4_X1    g152(.A1(new_n319), .A2(new_n344), .A3(new_n347), .A4(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n314), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n305), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n341), .A2(new_n346), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n352), .B(new_n343), .C1(new_n357), .C2(new_n342), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n353), .B1(new_n344), .B2(new_n347), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n359), .A3(new_n319), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n354), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n318), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n307), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n314), .B1(new_n305), .B2(new_n306), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT38), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n261), .A2(new_n265), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT83), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n335), .A2(new_n340), .ZN(new_n368));
  OR3_X1    g167(.A1(new_n368), .A2(KEYINPUT39), .A3(new_n338), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT40), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n352), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n368), .A2(new_n338), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT39), .B1(new_n345), .B2(new_n337), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n369), .B(new_n372), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n370), .A2(new_n371), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  OR2_X1    g177(.A1(new_n373), .A2(new_n374), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n379), .A2(new_n376), .A3(new_n369), .A4(new_n372), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n378), .A2(new_n358), .A3(new_n380), .ZN(new_n381));
  OR2_X1    g180(.A1(KEYINPUT75), .A2(KEYINPUT30), .ZN(new_n382));
  NAND2_X1  g181(.A1(KEYINPUT75), .A2(KEYINPUT30), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n305), .A2(new_n355), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n383), .B1(new_n305), .B2(new_n355), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n382), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n300), .A2(new_n296), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n217), .B1(new_n387), .B2(new_n303), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT74), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n302), .A4(new_n315), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n302), .B(new_n315), .C1(new_n304), .C2(new_n242), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT74), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n367), .B(new_n381), .C1(new_n386), .C2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n390), .A2(new_n392), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n396), .B(new_n382), .C1(new_n385), .C2(new_n384), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n367), .B1(new_n397), .B2(new_n381), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n366), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT84), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n366), .B(KEYINPUT84), .C1(new_n395), .C2(new_n398), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n300), .A2(new_n332), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n331), .B(new_n294), .C1(new_n298), .C2(new_n299), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AND2_X1   g205(.A1(G227gat), .A2(G233gat), .ZN(new_n407));
  AND2_X1   g206(.A1(KEYINPUT71), .A2(KEYINPUT34), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412));
  XOR2_X1   g211(.A(G71gat), .B(G99gat), .Z(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT70), .ZN(new_n414));
  XNOR2_X1  g213(.A(G15gat), .B(G43gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n411), .B(KEYINPUT32), .C1(new_n412), .C2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(KEYINPUT71), .A2(KEYINPUT34), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n416), .B1(new_n411), .B2(KEYINPUT32), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n411), .A2(KEYINPUT69), .A3(new_n412), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT69), .B1(new_n411), .B2(new_n412), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n417), .B(new_n419), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n411), .A2(new_n412), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT69), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(new_n421), .A3(new_n420), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n419), .B1(new_n429), .B2(new_n417), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n410), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n417), .B1(new_n422), .B2(new_n423), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n418), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(new_n409), .A3(new_n424), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT36), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n261), .A2(new_n265), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n354), .A2(new_n360), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n397), .A2(new_n439), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n431), .A2(KEYINPUT36), .A3(new_n434), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n436), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT35), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n431), .A2(new_n434), .B1(new_n261), .B2(new_n265), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(new_n440), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n434), .ZN(new_n447));
  AND4_X1   g246(.A1(new_n444), .A2(new_n447), .A3(new_n440), .A4(new_n437), .ZN(new_n448));
  OAI22_X1  g247(.A1(new_n403), .A2(new_n443), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT98), .ZN(new_n450));
  XNOR2_X1  g249(.A(G15gat), .B(G22gat), .ZN(new_n451));
  OR2_X1    g250(.A1(new_n451), .A2(G1gat), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT16), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n451), .B1(new_n453), .B2(G1gat), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G8gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n451), .A2(G1gat), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n456), .B1(new_n457), .B2(KEYINPUT88), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n455), .B(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(G57gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(G64gat), .ZN(new_n461));
  INV_X1    g260(.A(G64gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(G57gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(G71gat), .A2(G78gat), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT9), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT90), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(G71gat), .A3(G78gat), .ZN(new_n470));
  NOR2_X1   g269(.A1(G71gat), .A2(G78gat), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(KEYINPUT90), .B2(new_n465), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n468), .A2(KEYINPUT91), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT91), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n461), .A2(new_n463), .B1(new_n466), .B2(new_n465), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n465), .A2(KEYINPUT90), .ZN(new_n476));
  INV_X1    g275(.A(G71gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n255), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n470), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n474), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(new_n465), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n482), .A2(new_n464), .A3(new_n467), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT21), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n459), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n452), .A2(new_n454), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(new_n458), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n481), .A2(KEYINPUT92), .A3(new_n484), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT92), .B1(new_n481), .B2(new_n484), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n488), .B1(new_n491), .B2(KEYINPUT21), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n486), .B1(new_n492), .B2(new_n485), .ZN(new_n493));
  NAND2_X1  g292(.A1(G231gat), .A2(G233gat), .ZN(new_n494));
  INV_X1    g293(.A(G183gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G211gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n493), .B(new_n498), .Z(new_n499));
  XNOR2_X1  g298(.A(G127gat), .B(G155gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n499), .B(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G190gat), .B(G218gat), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT87), .ZN(new_n507));
  INV_X1    g306(.A(G29gat), .ZN(new_n508));
  INV_X1    g307(.A(G36gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT86), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT14), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n511), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(G29gat), .A2(G36gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT14), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n515), .A2(KEYINPUT86), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G43gat), .B(G50gat), .Z(new_n520));
  INV_X1    g319(.A(KEYINPUT15), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n508), .A2(new_n509), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(new_n520), .B2(new_n521), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n519), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n522), .B1(new_n519), .B2(new_n524), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n507), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n516), .B1(new_n515), .B2(KEYINPUT86), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(new_n511), .B2(new_n510), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n524), .B1(new_n529), .B2(new_n517), .ZN(new_n530));
  INV_X1    g329(.A(new_n522), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n519), .A2(new_n522), .A3(new_n524), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(KEYINPUT87), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n527), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G85gat), .A2(G92gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n536), .B(new_n537), .Z(new_n538));
  NOR2_X1   g337(.A1(G85gat), .A2(G92gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT8), .ZN(new_n540));
  NAND2_X1  g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n540), .B1(new_n541), .B2(KEYINPUT95), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT95), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n543), .A2(G99gat), .A3(G106gat), .ZN(new_n544));
  AOI211_X1 g343(.A(KEYINPUT96), .B(new_n539), .C1(new_n542), .C2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT96), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(KEYINPUT95), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n547), .A2(new_n544), .A3(KEYINPUT8), .ZN(new_n548));
  INV_X1    g347(.A(new_n539), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n538), .B1(new_n545), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G99gat), .B(G106gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n552), .B(new_n538), .C1(new_n545), .C2(new_n550), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n535), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT41), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT17), .B1(new_n527), .B2(new_n534), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n532), .A2(KEYINPUT17), .A3(new_n533), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n506), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n567));
  NOR3_X1   g366(.A1(new_n525), .A2(new_n526), .A3(new_n507), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT87), .B1(new_n532), .B2(new_n533), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(new_n563), .A3(new_n556), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n571), .A2(new_n558), .A3(new_n560), .A4(new_n505), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n566), .A2(new_n572), .A3(KEYINPUT93), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT97), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n559), .A2(KEYINPUT41), .ZN(new_n576));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n566), .A2(new_n572), .A3(KEYINPUT97), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n575), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n573), .A2(new_n574), .A3(new_n578), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n450), .B1(new_n504), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n583), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(KEYINPUT98), .A3(new_n503), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT99), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n481), .B(new_n484), .C1(new_n588), .C2(new_n552), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n548), .A2(new_n549), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT96), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n548), .A2(new_n546), .A3(new_n549), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n552), .B1(new_n593), .B2(new_n538), .ZN(new_n594));
  INV_X1    g393(.A(new_n555), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n589), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n552), .A2(new_n588), .ZN(new_n597));
  AOI211_X1 g396(.A(new_n597), .B(new_n483), .C1(new_n473), .C2(new_n480), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(new_n554), .A3(new_n555), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n601), .B(KEYINPUT101), .Z(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G120gat), .B(G148gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(G176gat), .B(G204gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT102), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT10), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n596), .A2(new_n609), .A3(new_n599), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT100), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n596), .A2(KEYINPUT100), .A3(new_n599), .A4(new_n609), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT10), .B1(new_n489), .B2(new_n490), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(new_n556), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n602), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n608), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n616), .B1(new_n612), .B2(new_n613), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n621), .A2(KEYINPUT102), .A3(new_n602), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n603), .B(new_n607), .C1(new_n620), .C2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n602), .B(KEYINPUT103), .Z(new_n624));
  OR2_X1    g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n603), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n606), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n587), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n488), .B1(new_n568), .B2(new_n569), .ZN(new_n631));
  NAND2_X1  g430(.A1(G229gat), .A2(G233gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n459), .A2(new_n563), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n631), .B(new_n632), .C1(new_n562), .C2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT18), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n459), .A2(new_n563), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n570), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n638), .A2(KEYINPUT18), .A3(new_n632), .A4(new_n631), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n632), .B(KEYINPUT13), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n631), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n535), .A2(new_n488), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n636), .A2(new_n639), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n646));
  XNOR2_X1  g445(.A(G113gat), .B(G141gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(G169gat), .B(G197gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT12), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n645), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n636), .A2(new_n639), .A3(new_n644), .ZN(new_n653));
  INV_X1    g452(.A(new_n651), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(KEYINPUT89), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n630), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n449), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n439), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  INV_X1    g462(.A(new_n397), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT42), .B1(new_n665), .B2(new_n456), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT104), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(new_n456), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  MUX2_X1   g468(.A(KEYINPUT42), .B(new_n666), .S(new_n669), .Z(G1325gat));
  INV_X1    g469(.A(G15gat), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n431), .A2(KEYINPUT36), .A3(new_n434), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n435), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n660), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n661), .A2(new_n447), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n674), .B1(new_n671), .B2(new_n675), .ZN(G1326gat));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n437), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  NAND2_X1  g478(.A1(new_n449), .A2(new_n583), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n673), .A2(new_n401), .A3(new_n441), .A4(new_n402), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n447), .A2(new_n440), .A3(new_n437), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT35), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n445), .A2(new_n444), .A3(new_n440), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n585), .B1(new_n683), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT44), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n628), .A2(KEYINPUT105), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n628), .A2(KEYINPUT105), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n656), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n682), .A2(new_n504), .A3(new_n689), .A4(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G29gat), .B1(new_n696), .B2(new_n438), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n658), .A2(new_n503), .A3(new_n628), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n688), .A2(new_n508), .A3(new_n439), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT45), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT106), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n697), .A2(new_n703), .A3(new_n700), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(G1328gat));
  OAI21_X1  g504(.A(G36gat), .B1(new_n696), .B2(new_n664), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n688), .A2(new_n509), .A3(new_n397), .A4(new_n698), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT46), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n708), .A2(KEYINPUT107), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(KEYINPUT107), .ZN(new_n710));
  OAI221_X1 g509(.A(new_n706), .B1(KEYINPUT46), .B2(new_n707), .C1(new_n709), .C2(new_n710), .ZN(G1329gat));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(KEYINPUT108), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n688), .A2(new_n698), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n447), .ZN(new_n715));
  INV_X1    g514(.A(G43gat), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n713), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n504), .B1(new_n688), .B2(KEYINPUT44), .ZN(new_n718));
  AOI211_X1 g517(.A(new_n681), .B(new_n585), .C1(new_n683), .C2(new_n687), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n673), .A2(new_n716), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n695), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n712), .A2(KEYINPUT108), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n717), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n723), .B1(new_n717), .B2(new_n722), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(G1330gat));
  OAI21_X1  g525(.A(G50gat), .B1(new_n696), .B2(new_n437), .ZN(new_n727));
  INV_X1    g526(.A(G50gat), .ZN(new_n728));
  INV_X1    g527(.A(new_n437), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT48), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n727), .A2(KEYINPUT48), .A3(new_n730), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(G1331gat));
  AND3_X1   g534(.A1(new_n587), .A2(new_n694), .A3(new_n693), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n449), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n438), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(new_n460), .ZN(G1332gat));
  NOR2_X1   g538(.A1(new_n737), .A2(new_n664), .ZN(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  AND2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n740), .B2(new_n741), .ZN(G1333gat));
  OR3_X1    g543(.A1(new_n737), .A2(new_n477), .A3(new_n673), .ZN(new_n745));
  INV_X1    g544(.A(new_n447), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n477), .B1(new_n737), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g548(.A1(new_n737), .A2(new_n437), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(new_n255), .ZN(G1335gat));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n449), .A2(KEYINPUT109), .A3(new_n583), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n503), .A2(new_n656), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n688), .A2(KEYINPUT109), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n754), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n758), .B1(new_n688), .B2(KEYINPUT109), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n680), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n759), .A2(new_n761), .A3(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n763), .A2(new_n349), .A3(new_n439), .A4(new_n628), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n629), .A2(new_n656), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n682), .A2(new_n504), .A3(new_n689), .A4(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766), .B2(new_n438), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(G1336gat));
  INV_X1    g567(.A(G92gat), .ZN(new_n769));
  INV_X1    g568(.A(new_n765), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n718), .A2(new_n719), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n769), .B1(new_n771), .B2(new_n397), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n692), .A2(new_n664), .A3(G92gat), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n757), .B2(new_n762), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT52), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n755), .A2(new_n756), .A3(new_n752), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT51), .B1(new_n759), .B2(new_n761), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n773), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  OAI21_X1  g579(.A(G92gat), .B1(new_n766), .B2(new_n664), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n776), .A2(new_n782), .ZN(G1337gat));
  NOR2_X1   g582(.A1(new_n746), .A2(G99gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n763), .A2(new_n628), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(G99gat), .B1(new_n766), .B2(new_n673), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(G1338gat));
  AOI21_X1  g586(.A(new_n259), .B1(new_n771), .B2(new_n729), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n437), .A2(new_n692), .A3(G106gat), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n757), .B2(new_n762), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT53), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n789), .B1(new_n777), .B2(new_n778), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794));
  OAI21_X1  g593(.A(G106gat), .B1(new_n766), .B2(new_n437), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n796), .ZN(G1339gat));
  NAND2_X1  g596(.A1(new_n447), .A2(new_n437), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n614), .A2(new_n617), .A3(new_n624), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT54), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT102), .B1(new_n621), .B2(new_n602), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n618), .A2(new_n608), .A3(new_n619), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n606), .B1(new_n625), .B2(KEYINPUT54), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n799), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(new_n621), .B2(new_n624), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n620), .B2(new_n622), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n621), .A2(new_n624), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n607), .B1(new_n810), .B2(new_n807), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n809), .A2(KEYINPUT55), .A3(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n806), .A2(new_n812), .A3(new_n656), .A4(new_n623), .ZN(new_n813));
  INV_X1    g612(.A(new_n632), .ZN(new_n814));
  INV_X1    g613(.A(new_n638), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n642), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT110), .ZN(new_n817));
  OR3_X1    g616(.A1(new_n642), .A2(new_n643), .A3(new_n641), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT110), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n819), .B(new_n814), .C1(new_n815), .C2(new_n642), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n821), .A2(new_n650), .B1(new_n651), .B2(new_n645), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n628), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n583), .B1(new_n813), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n806), .A2(new_n623), .A3(new_n812), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n583), .A2(new_n822), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OR3_X1    g626(.A1(new_n824), .A2(new_n827), .A3(KEYINPUT111), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT111), .B1(new_n824), .B2(new_n827), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n504), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n587), .A2(new_n694), .A3(new_n629), .ZN(new_n831));
  AOI211_X1 g630(.A(new_n438), .B(new_n798), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n664), .ZN(new_n833));
  OAI21_X1  g632(.A(G113gat), .B1(new_n833), .B2(new_n658), .ZN(new_n834));
  XOR2_X1   g633(.A(new_n834), .B(KEYINPUT112), .Z(new_n835));
  INV_X1    g634(.A(new_n833), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(new_n324), .A3(new_n656), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(G1340gat));
  OAI21_X1  g637(.A(G120gat), .B1(new_n833), .B2(new_n692), .ZN(new_n839));
  XOR2_X1   g638(.A(new_n839), .B(KEYINPUT113), .Z(new_n840));
  NAND2_X1  g639(.A1(new_n628), .A2(new_n327), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT114), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n840), .B1(new_n833), .B2(new_n842), .ZN(G1341gat));
  NAND2_X1  g642(.A1(new_n836), .A2(new_n503), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g644(.A1(new_n397), .A2(new_n585), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n846), .B(KEYINPUT115), .Z(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(G134gat), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT56), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n849), .A2(KEYINPUT56), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n832), .A2(new_n848), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n832), .A2(new_n848), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(G134gat), .B1(new_n833), .B2(new_n585), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n855), .A2(KEYINPUT116), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(KEYINPUT116), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n860), .B(new_n854), .C1(new_n856), .C2(new_n857), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(G1343gat));
  NOR4_X1   g661(.A1(new_n672), .A2(new_n435), .A3(new_n438), .A4(new_n397), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n657), .A2(new_n623), .A3(new_n812), .A4(new_n806), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n583), .B1(new_n864), .B2(new_n823), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n504), .B1(new_n865), .B2(new_n827), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n831), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(KEYINPUT57), .A3(new_n729), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n829), .A2(new_n504), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n824), .A2(new_n827), .A3(KEYINPUT111), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n831), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT57), .B1(new_n871), .B2(new_n729), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n868), .B1(new_n872), .B2(KEYINPUT119), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n437), .B1(new_n830), .B2(new_n831), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT57), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n656), .B(new_n863), .C1(new_n873), .C2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n229), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(KEYINPUT120), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n658), .A2(G141gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n874), .A2(new_n863), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT120), .B1(new_n877), .B2(new_n878), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT58), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n874), .A2(new_n439), .A3(new_n673), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n885), .B(KEYINPUT121), .Z(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n664), .A3(new_n880), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n863), .B1(new_n873), .B2(new_n876), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n878), .B1(new_n888), .B2(new_n658), .ZN(new_n889));
  XOR2_X1   g688(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n890));
  NAND3_X1  g689(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n884), .A2(new_n891), .ZN(G1344gat));
  NAND4_X1  g691(.A1(new_n886), .A2(new_n227), .A3(new_n664), .A4(new_n628), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n888), .A2(new_n629), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(KEYINPUT59), .A3(new_n227), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n871), .A2(new_n729), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT57), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n866), .B1(new_n630), .B2(new_n657), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n900), .A3(new_n729), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n628), .A3(new_n863), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n896), .B1(new_n903), .B2(G148gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n893), .B1(new_n895), .B2(new_n904), .ZN(G1345gat));
  NOR3_X1   g704(.A1(new_n888), .A2(new_n222), .A3(new_n504), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n886), .A2(new_n664), .A3(new_n503), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(new_n222), .ZN(G1346gat));
  INV_X1    g707(.A(new_n847), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n886), .A2(new_n223), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G162gat), .B1(new_n888), .B2(new_n585), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1347gat));
  AOI21_X1  g711(.A(new_n439), .B1(new_n830), .B2(new_n831), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n798), .A2(new_n664), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G169gat), .B1(new_n915), .B2(new_n658), .ZN(new_n916));
  XOR2_X1   g715(.A(new_n914), .B(KEYINPUT123), .Z(new_n917));
  AND3_X1   g716(.A1(new_n917), .A2(KEYINPUT124), .A3(new_n913), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT124), .B1(new_n917), .B2(new_n913), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n656), .A2(new_n270), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(G1348gat));
  NOR3_X1   g721(.A1(new_n915), .A2(new_n271), .A3(new_n692), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n628), .B1(new_n918), .B2(new_n919), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n924), .B2(new_n271), .ZN(G1349gat));
  NAND4_X1  g724(.A1(new_n917), .A2(new_n287), .A3(new_n503), .A4(new_n913), .ZN(new_n926));
  OAI21_X1  g725(.A(G183gat), .B1(new_n915), .B2(new_n504), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT60), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n928), .B(new_n930), .ZN(G1350gat));
  OR2_X1    g730(.A1(new_n585), .A2(new_n268), .ZN(new_n932));
  OAI21_X1  g731(.A(G190gat), .B1(new_n915), .B2(new_n585), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n933), .A2(KEYINPUT61), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n933), .A2(KEYINPUT61), .ZN(new_n935));
  OAI22_X1  g734(.A1(new_n920), .A2(new_n932), .B1(new_n934), .B2(new_n935), .ZN(G1351gat));
  NAND3_X1  g735(.A1(new_n673), .A2(new_n438), .A3(new_n397), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT126), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n902), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(G197gat), .B1(new_n939), .B2(new_n658), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n897), .A2(new_n937), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n941), .A2(new_n212), .A3(new_n656), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(G1352gat));
  NAND3_X1  g742(.A1(new_n941), .A2(new_n213), .A3(new_n628), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n944), .B(KEYINPUT62), .Z(new_n945));
  OAI21_X1  g744(.A(G204gat), .B1(new_n939), .B2(new_n692), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1353gat));
  NOR2_X1   g746(.A1(new_n937), .A2(new_n504), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n497), .A3(new_n874), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n898), .A2(new_n901), .A3(new_n948), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n950), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT63), .B1(new_n950), .B2(G211gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n953), .B(new_n954), .ZN(G1354gat));
  NAND2_X1  g754(.A1(new_n583), .A2(G218gat), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n897), .A2(new_n585), .A3(new_n937), .ZN(new_n957));
  OAI22_X1  g756(.A1(new_n939), .A2(new_n956), .B1(new_n957), .B2(G218gat), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(G1355gat));
endmodule


