//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1243,
    new_n1244, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1304, new_n1305;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n213), .A2(G20), .A3(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT64), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n208), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n211), .B(new_n216), .C1(new_n223), .C2(KEYINPUT1), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G87), .B(G97), .Z(new_n234));
  XOR2_X1   g0034(.A(G107), .B(G116), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  INV_X1    g0040(.A(G33), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(KEYINPUT3), .ZN(new_n242));
  INV_X1    g0042(.A(KEYINPUT3), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G33), .ZN(new_n244));
  INV_X1    g0044(.A(G1698), .ZN(new_n245));
  NAND4_X1  g0045(.A1(new_n242), .A2(new_n244), .A3(G226), .A4(new_n245), .ZN(new_n246));
  NAND4_X1  g0046(.A1(new_n242), .A2(new_n244), .A3(G232), .A4(G1698), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G97), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n255));
  AND3_X1   g0055(.A1(new_n251), .A2(KEYINPUT65), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT65), .B1(new_n251), .B2(new_n255), .ZN(new_n257));
  OAI21_X1  g0057(.A(G238), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(new_n251), .A3(G274), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n253), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT13), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT13), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n253), .A2(new_n258), .A3(new_n265), .A4(new_n262), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(KEYINPUT66), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT66), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n263), .A2(new_n268), .A3(KEYINPUT13), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(G169), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT69), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n267), .A2(KEYINPUT69), .A3(G169), .A4(new_n269), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(KEYINPUT14), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT70), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n272), .A2(KEYINPUT70), .A3(KEYINPUT14), .A4(new_n273), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n264), .B(KEYINPUT67), .ZN(new_n278));
  XOR2_X1   g0078(.A(new_n266), .B(KEYINPUT68), .Z(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(new_n279), .A3(G179), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT14), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n267), .A2(new_n281), .A3(G169), .A4(new_n269), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n276), .A2(new_n277), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G13), .ZN(new_n285));
  INV_X1    g0085(.A(G20), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n285), .A2(new_n286), .A3(G1), .ZN(new_n287));
  INV_X1    g0087(.A(G68), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT12), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n291), .A2(G50), .B1(G20), .B2(new_n288), .ZN(new_n292));
  INV_X1    g0092(.A(G77), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n286), .A2(G33), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n214), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(KEYINPUT11), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n287), .A2(new_n297), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n254), .A2(G20), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(G68), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n290), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT11), .B1(new_n295), .B2(new_n297), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n284), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n278), .A2(new_n279), .A3(G190), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n267), .A2(G200), .A3(new_n269), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n299), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT8), .B(G58), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n300), .ZN(new_n314));
  INV_X1    g0114(.A(new_n287), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n311), .A2(new_n314), .B1(new_n315), .B2(new_n313), .ZN(new_n316));
  INV_X1    g0116(.A(G58), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(new_n288), .ZN(new_n318));
  OAI21_X1  g0118(.A(G20), .B1(new_n318), .B2(new_n201), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n291), .A2(G159), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n319), .A2(KEYINPUT73), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT73), .B1(new_n319), .B2(new_n320), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n243), .A2(G33), .ZN(new_n324));
  AND2_X1   g0124(.A1(KEYINPUT71), .A2(KEYINPUT3), .ZN(new_n325));
  NOR2_X1   g0125(.A1(KEYINPUT71), .A2(KEYINPUT3), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n324), .B1(new_n327), .B2(G33), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT7), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(G20), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT72), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n325), .A2(new_n326), .A3(new_n241), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(new_n334), .B2(new_n324), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT71), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n243), .ZN(new_n337));
  NAND2_X1  g0137(.A1(KEYINPUT71), .A2(KEYINPUT3), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(G33), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(KEYINPUT72), .A3(new_n242), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n335), .A2(new_n286), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n332), .B1(new_n341), .B2(new_n329), .ZN(new_n342));
  OAI211_X1 g0142(.A(KEYINPUT16), .B(new_n323), .C1(new_n342), .C2(new_n288), .ZN(new_n343));
  INV_X1    g0143(.A(new_n297), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n241), .B1(new_n325), .B2(new_n326), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n331), .B1(new_n345), .B2(new_n244), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n242), .A2(new_n244), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT7), .B1(new_n347), .B2(new_n286), .ZN(new_n348));
  OAI21_X1  g0148(.A(G68), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n323), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT16), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n344), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n316), .B1(new_n343), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n251), .A2(G232), .A3(new_n255), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n262), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G33), .A2(G87), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  MUX2_X1   g0157(.A(G223), .B(G226), .S(G1698), .Z(new_n358));
  AOI21_X1  g0158(.A(new_n357), .B1(new_n328), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n355), .B1(new_n359), .B2(new_n251), .ZN(new_n360));
  INV_X1    g0160(.A(G169), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT74), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n262), .A2(new_n354), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n363), .B1(new_n262), .B2(new_n354), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n359), .B2(new_n251), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n362), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT18), .B1(new_n353), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n343), .A2(new_n352), .ZN(new_n372));
  INV_X1    g0172(.A(new_n316), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT18), .ZN(new_n375));
  INV_X1    g0175(.A(new_n370), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n358), .A2(new_n339), .A3(new_n242), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n356), .ZN(new_n380));
  AOI21_X1  g0180(.A(G190), .B1(new_n380), .B2(new_n252), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n360), .A2(new_n378), .B1(new_n381), .B2(new_n366), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(KEYINPUT75), .A2(KEYINPUT17), .ZN(new_n384));
  AND4_X1   g0184(.A1(new_n372), .A2(new_n383), .A3(new_n373), .A4(new_n384), .ZN(new_n385));
  XOR2_X1   g0185(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n353), .B2(new_n383), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n371), .B(new_n377), .C1(new_n385), .C2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n241), .A2(KEYINPUT3), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n324), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G1698), .ZN(new_n391));
  INV_X1    g0191(.A(G223), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n391), .A2(new_n392), .B1(new_n293), .B2(new_n390), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n390), .A2(G222), .A3(new_n245), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n252), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n256), .A2(new_n257), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G226), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n262), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G200), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n291), .A2(G150), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(new_n312), .B2(new_n294), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(G20), .B2(new_n203), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n344), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT9), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n300), .A2(G50), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n311), .A2(new_n405), .B1(G50), .B2(new_n315), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n403), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n395), .A2(G190), .A3(new_n262), .A4(new_n397), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n404), .B1(new_n403), .B2(new_n406), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n399), .A2(new_n408), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n411), .B(KEYINPUT10), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n403), .A2(new_n406), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n398), .B2(new_n361), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(G179), .B2(new_n398), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n313), .A2(new_n291), .B1(G20), .B2(G77), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT15), .B(G87), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n417), .A2(new_n294), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n344), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n299), .A2(G77), .A3(new_n300), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(G77), .B2(new_n315), .ZN(new_n421));
  OR2_X1    g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n390), .A2(G232), .A3(new_n245), .ZN(new_n423));
  INV_X1    g0223(.A(G107), .ZN(new_n424));
  INV_X1    g0224(.A(G238), .ZN(new_n425));
  OAI221_X1 g0225(.A(new_n423), .B1(new_n424), .B2(new_n390), .C1(new_n391), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n252), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n396), .A2(G244), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n262), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n422), .B1(new_n430), .B2(G190), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(G200), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n422), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n361), .B2(new_n429), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n430), .A2(new_n368), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n412), .A2(new_n415), .A3(new_n433), .A4(new_n437), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n310), .A2(new_n388), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n329), .B1(new_n390), .B2(G20), .ZN(new_n441));
  AOI21_X1  g0241(.A(G33), .B1(new_n337), .B2(new_n338), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n330), .B1(new_n442), .B2(new_n389), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n424), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n291), .A2(G77), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT76), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(KEYINPUT6), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT6), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(KEYINPUT76), .ZN(new_n449));
  INV_X1    g0249(.A(G97), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n447), .A2(new_n449), .B1(new_n450), .B2(G107), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(KEYINPUT76), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n446), .A2(KEYINPUT6), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G97), .A2(G107), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n206), .A2(new_n452), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n445), .B1(new_n456), .B2(new_n286), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n297), .B1(new_n444), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT77), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n315), .A2(G97), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n254), .A2(G33), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n299), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n460), .B1(new_n463), .B2(G97), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n458), .A2(new_n459), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n459), .B1(new_n458), .B2(new_n464), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G274), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n468), .B1(new_n215), .B2(new_n250), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n254), .B(G45), .C1(new_n259), .C2(KEYINPUT5), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT79), .B1(new_n472), .B2(G41), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT79), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(new_n259), .A3(KEYINPUT5), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n469), .A2(new_n471), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G257), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n472), .A2(G41), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n251), .B1(new_n470), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n476), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n390), .A2(G250), .A3(G1698), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT4), .ZN(new_n482));
  INV_X1    g0282(.A(G244), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n390), .A2(new_n245), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n481), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n339), .A2(G244), .A3(new_n245), .A4(new_n242), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT78), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n488), .A2(new_n489), .A3(new_n482), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(new_n488), .B2(new_n482), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n480), .B1(new_n492), .B2(new_n252), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G190), .ZN(new_n494));
  OAI21_X1  g0294(.A(G200), .B1(new_n493), .B2(KEYINPUT80), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT80), .ZN(new_n496));
  AOI211_X1 g0296(.A(new_n496), .B(new_n480), .C1(new_n492), .C2(new_n252), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n467), .B(new_n494), .C1(new_n495), .C2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n480), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n481), .A2(new_n485), .A3(new_n486), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n488), .A2(new_n482), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT78), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n488), .A2(new_n489), .A3(new_n482), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n499), .B1(new_n504), .B2(new_n251), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G169), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n493), .A2(G179), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n458), .A2(new_n464), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(G87), .ZN(new_n511));
  OR4_X1    g0311(.A1(KEYINPUT22), .A2(new_n347), .A3(G20), .A4(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n339), .A2(new_n286), .A3(G87), .A4(new_n242), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n513), .A2(KEYINPUT84), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT22), .B1(new_n513), .B2(KEYINPUT84), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT24), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT23), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n286), .B2(G107), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n424), .A2(KEYINPUT23), .A3(G20), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G116), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n519), .A2(new_n520), .B1(new_n522), .B2(new_n286), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n516), .A2(new_n517), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n517), .B1(new_n516), .B2(new_n523), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n297), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(G264), .B(new_n251), .C1(new_n470), .C2(new_n478), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(G250), .A2(G1698), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n477), .B2(G1698), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n328), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G294), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n528), .B1(new_n533), .B2(new_n252), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n378), .B1(new_n534), .B2(new_n476), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n534), .A2(new_n476), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n535), .B1(G190), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT86), .B1(new_n315), .B2(G107), .ZN(new_n538));
  XOR2_X1   g0338(.A(KEYINPUT85), .B(KEYINPUT25), .Z(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n315), .A2(KEYINPUT86), .A3(G107), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n540), .B(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(G107), .B2(new_n463), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n526), .A2(new_n537), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n498), .A2(new_n510), .A3(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n260), .A2(G1), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n546), .A2(G250), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n468), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n251), .A3(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(G238), .A2(G1698), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n483), .B2(G1698), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n522), .B1(new_n328), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n368), .B(new_n549), .C1(new_n552), .C2(new_n251), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n339), .A3(new_n242), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n251), .B1(new_n554), .B2(new_n521), .ZN(new_n555));
  INV_X1    g0355(.A(new_n549), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n361), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT81), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT81), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n553), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n205), .A2(new_n511), .B1(new_n248), .B2(new_n286), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT19), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G97), .ZN(new_n564));
  OAI22_X1  g0364(.A1(new_n562), .A2(new_n563), .B1(new_n294), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n339), .A2(new_n286), .A3(G68), .A4(new_n242), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n344), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n417), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(new_n315), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n463), .A2(new_n568), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n559), .A2(new_n561), .A3(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n555), .A2(new_n556), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G190), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n462), .A2(new_n511), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n567), .A2(new_n576), .A3(new_n569), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(G200), .B1(new_n555), .B2(new_n556), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  MUX2_X1   g0381(.A(G257), .B(G264), .S(G1698), .Z(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(new_n339), .A3(new_n242), .ZN(new_n583));
  XNOR2_X1  g0383(.A(KEYINPUT83), .B(G303), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n347), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n251), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT82), .ZN(new_n588));
  OAI211_X1 g0388(.A(G270), .B(new_n251), .C1(new_n470), .C2(new_n478), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n476), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n588), .B1(new_n476), .B2(new_n589), .ZN(new_n592));
  OAI211_X1 g0392(.A(G190), .B(new_n587), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n486), .B(new_n286), .C1(G33), .C2(new_n450), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n594), .B(new_n297), .C1(new_n286), .C2(G116), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n595), .B(KEYINPUT20), .ZN(new_n596));
  INV_X1    g0396(.A(G116), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n287), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n462), .B2(new_n597), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n472), .A2(G41), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n473), .A2(new_n475), .A3(new_n601), .A4(new_n546), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n251), .A2(G274), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n589), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT82), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n586), .B1(new_n606), .B2(new_n590), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n593), .B(new_n600), .C1(new_n378), .C2(new_n607), .ZN(new_n608));
  AOI211_X1 g0408(.A(new_n368), .B(new_n586), .C1(new_n606), .C2(new_n590), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT20), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n595), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n463), .A2(G116), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n598), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT21), .ZN(new_n615));
  OAI21_X1  g0415(.A(G169), .B1(new_n596), .B2(new_n599), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n615), .B1(new_n616), .B2(new_n607), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(new_n613), .A3(KEYINPUT21), .A4(G169), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n608), .A2(new_n614), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n581), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n526), .A2(new_n543), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n534), .A2(new_n476), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n623), .A2(G179), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(new_n361), .B2(new_n623), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n440), .A2(new_n545), .A3(new_n627), .ZN(G372));
  INV_X1    g0428(.A(new_n553), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT87), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n555), .A2(new_n630), .ZN(new_n631));
  AOI211_X1 g0431(.A(KEYINPUT87), .B(new_n251), .C1(new_n554), .C2(new_n521), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n549), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI211_X1 g0433(.A(KEYINPUT88), .B(new_n629), .C1(new_n633), .C2(new_n361), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT88), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n361), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n635), .B1(new_n636), .B2(new_n553), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n572), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n633), .A2(G200), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n578), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n498), .A2(new_n510), .A3(new_n544), .A4(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n614), .A2(new_n617), .A3(new_n619), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n622), .B2(new_n625), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n638), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n509), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n506), .B2(new_n507), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n558), .A2(KEYINPUT81), .B1(new_n570), .B2(new_n571), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n647), .A2(new_n561), .B1(new_n578), .B2(new_n579), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n646), .A2(new_n648), .A3(KEYINPUT26), .ZN(new_n649));
  INV_X1    g0449(.A(new_n466), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n458), .A2(new_n459), .A3(new_n464), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n506), .A2(new_n507), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n638), .A2(new_n640), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n644), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n439), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n377), .A2(new_n371), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n437), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n284), .B2(new_n305), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n309), .B1(new_n387), .B2(new_n385), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT89), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT89), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n665), .B(new_n659), .C1(new_n661), .C2(new_n662), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n412), .A3(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n667), .A2(KEYINPUT90), .A3(new_n415), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT90), .B1(new_n667), .B2(new_n415), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n657), .B1(new_n668), .B2(new_n669), .ZN(G369));
  NAND3_X1  g0470(.A1(new_n254), .A2(new_n286), .A3(G13), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G343), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n626), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n622), .A2(new_n676), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n678), .A2(new_n544), .B1(new_n622), .B2(new_n625), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(new_n677), .ZN(new_n680));
  INV_X1    g0480(.A(new_n642), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n676), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n677), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n676), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n600), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n642), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n620), .B2(new_n685), .ZN(new_n687));
  XOR2_X1   g0487(.A(KEYINPUT91), .B(G330), .Z(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n680), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n683), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n209), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G1), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n212), .B2(new_n696), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n701), .B(new_n684), .C1(new_n644), .C2(new_n655), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n510), .A2(KEYINPUT26), .A3(new_n581), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n653), .B2(KEYINPUT26), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n498), .A2(new_n510), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n626), .A2(new_n681), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n705), .A2(new_n706), .A3(new_n544), .A4(new_n640), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n707), .A3(new_n638), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n708), .A2(new_n684), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n702), .B1(new_n709), .B2(new_n701), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n627), .A2(new_n545), .A3(new_n676), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n607), .A2(G179), .A3(new_n534), .A4(new_n574), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n505), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n534), .A2(new_n574), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n493), .A2(new_n715), .A3(new_n609), .A4(KEYINPUT30), .ZN(new_n716));
  AOI21_X1  g0516(.A(G179), .B1(new_n534), .B2(new_n476), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n505), .A2(new_n717), .A3(new_n618), .A4(new_n633), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n714), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n676), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT31), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g0522(.A(KEYINPUT92), .B(KEYINPUT31), .Z(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n689), .B1(new_n711), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n710), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n700), .B1(new_n728), .B2(G1), .ZN(G364));
  NOR2_X1   g0529(.A1(new_n285), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n254), .B1(new_n730), .B2(G45), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n695), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n390), .A2(G355), .A3(new_n209), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(G116), .B2(new_n209), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT93), .Z(new_n736));
  NAND2_X1  g0536(.A1(new_n335), .A2(new_n340), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n694), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n212), .A2(G45), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n739), .B1(new_n239), .B2(G45), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n736), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT94), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n214), .B1(G20), .B2(new_n361), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n733), .B1(new_n741), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n286), .A2(G179), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G190), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G159), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G190), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n749), .A2(new_n755), .A3(G200), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n754), .A2(KEYINPUT32), .B1(G107), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n749), .A2(G190), .A3(G200), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n758), .B1(new_n511), .B2(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n755), .A2(G179), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n286), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n390), .B1(new_n762), .B2(new_n450), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n286), .A2(new_n368), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G190), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n767), .A2(new_n288), .B1(new_n754), .B2(KEYINPUT32), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n760), .A2(new_n763), .A3(new_n768), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n764), .A2(KEYINPUT95), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n764), .A2(KEYINPUT95), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n755), .A2(G200), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n765), .A2(new_n755), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n774), .A2(G58), .B1(G50), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n770), .A2(new_n750), .A3(new_n771), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n777), .A2(KEYINPUT96), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(KEYINPUT96), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n776), .B1(new_n780), .B2(new_n293), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n781), .A2(KEYINPUT97), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(KEYINPUT97), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n769), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT98), .ZN(new_n785));
  INV_X1    g0585(.A(new_n751), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n390), .B1(new_n786), .B2(G329), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT33), .B(G317), .Z(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n767), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n777), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(G311), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n762), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n792), .A2(G294), .B1(new_n757), .B2(G283), .ZN(new_n793));
  INV_X1    g0593(.A(new_n759), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n775), .A2(G326), .B1(new_n794), .B2(G303), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n774), .A2(G322), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n791), .A2(new_n793), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n784), .A2(KEYINPUT98), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n785), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n748), .B1(new_n799), .B2(new_n745), .ZN(new_n800));
  INV_X1    g0600(.A(new_n744), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n687), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n691), .A2(new_n733), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n689), .B2(new_n687), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  NOR2_X1   g0606(.A1(new_n437), .A2(new_n676), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n433), .B1(new_n434), .B2(new_n684), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(new_n808), .B2(new_n437), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n656), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n811), .B2(new_n676), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n684), .B(new_n809), .C1(new_n644), .C2(new_n655), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n733), .B1(new_n814), .B2(new_n725), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n725), .B2(new_n814), .ZN(new_n816));
  INV_X1    g0616(.A(new_n733), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n745), .A2(new_n742), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(new_n293), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n745), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n780), .A2(new_n597), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n775), .A2(G303), .ZN(new_n822));
  INV_X1    g0622(.A(G283), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n767), .B2(new_n823), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n511), .A2(new_n756), .B1(new_n759), .B2(new_n424), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n390), .B1(new_n786), .B2(G311), .ZN(new_n826));
  INV_X1    g0626(.A(G294), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n826), .B1(new_n450), .B2(new_n762), .C1(new_n773), .C2(new_n827), .ZN(new_n828));
  NOR4_X1   g0628(.A1(new_n821), .A2(new_n824), .A3(new_n825), .A4(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n737), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n792), .A2(G58), .B1(new_n794), .B2(G50), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n288), .B2(new_n756), .C1(new_n832), .C2(new_n751), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n766), .A2(G150), .B1(new_n775), .B2(G137), .ZN(new_n834));
  INV_X1    g0634(.A(G143), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n835), .B2(new_n773), .C1(new_n780), .C2(new_n752), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n830), .B(new_n833), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n829), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n819), .B1(new_n820), .B2(new_n840), .C1(new_n809), .C2(new_n743), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n816), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G384));
  NOR3_X1   g0643(.A1(new_n214), .A2(new_n286), .A3(new_n597), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT35), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n844), .B1(new_n456), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(new_n845), .B2(new_n456), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT36), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n213), .B(G77), .C1(new_n317), .C2(new_n288), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n202), .A2(G68), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n254), .B(G13), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n306), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n684), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n372), .A2(new_n383), .A3(new_n373), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n353), .B2(new_n370), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n353), .A2(new_n674), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT37), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n374), .A2(new_n376), .ZN(new_n860));
  INV_X1    g0660(.A(new_n674), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n374), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n860), .A2(new_n862), .A3(new_n863), .A4(new_n856), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n388), .A2(new_n858), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g0667(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT39), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n323), .B1(new_n342), .B2(new_n288), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n351), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n297), .A3(new_n343), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n674), .B1(new_n873), .B2(new_n373), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n388), .A2(new_n874), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n316), .B(new_n382), .C1(new_n343), .C2(new_n352), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n871), .A2(new_n351), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n343), .A2(new_n297), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n373), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n876), .B1(new_n879), .B2(new_n376), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n861), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n863), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n864), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n875), .B(KEYINPUT38), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n869), .A2(new_n870), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n875), .B1(new_n882), .B2(new_n883), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n870), .B1(new_n888), .B2(new_n884), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n885), .A2(new_n889), .A3(KEYINPUT100), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT100), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n370), .B1(new_n873), .B2(new_n373), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n874), .A2(new_n892), .A3(new_n876), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n864), .B1(new_n893), .B2(new_n863), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n894), .B2(new_n875), .ZN(new_n895));
  INV_X1    g0695(.A(new_n884), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT39), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n869), .A2(new_n870), .A3(new_n884), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n891), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n855), .B1(new_n890), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n807), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n813), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n304), .A2(new_n684), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n306), .A2(new_n309), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n309), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n305), .B(new_n676), .C1(new_n284), .C2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n888), .A2(new_n884), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n909), .A2(new_n911), .B1(new_n659), .B2(new_n861), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n900), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT102), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n701), .B1(new_n708), .B2(new_n684), .ZN(new_n916));
  INV_X1    g0716(.A(new_n702), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n439), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT101), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT101), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n439), .B(new_n920), .C1(new_n916), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n668), .B2(new_n669), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n915), .B(new_n923), .Z(new_n924));
  NOR2_X1   g0724(.A1(new_n627), .A2(new_n545), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n684), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n720), .A2(new_n723), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n439), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT103), .Z(new_n933));
  OAI21_X1  g0733(.A(new_n809), .B1(new_n711), .B2(new_n929), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n905), .B2(new_n907), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT40), .B1(new_n935), .B2(new_n910), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT40), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n869), .B2(new_n884), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n936), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n688), .B1(new_n933), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n939), .B2(new_n933), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n924), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n254), .B2(new_n730), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n924), .A2(new_n941), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n852), .B1(new_n943), .B2(new_n944), .ZN(G367));
  OAI21_X1  g0745(.A(new_n705), .B1(new_n467), .B2(new_n684), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n652), .A2(new_n676), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n683), .A2(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT44), .Z(new_n950));
  NAND2_X1  g0750(.A1(new_n683), .A2(new_n948), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT105), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(KEYINPUT105), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT45), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(KEYINPUT45), .A3(new_n953), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n692), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n680), .B(new_n682), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(new_n690), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n727), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n955), .A2(new_n692), .A3(new_n956), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n959), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n964), .A2(new_n728), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n695), .B(KEYINPUT41), .Z(new_n966));
  OAI21_X1  g0766(.A(new_n731), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n958), .A2(new_n948), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT104), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n577), .A2(new_n684), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n638), .A2(new_n640), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n638), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n969), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n975));
  INV_X1    g0775(.A(new_n948), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n510), .B1(new_n976), .B2(new_n626), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n684), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n948), .A2(new_n680), .A3(new_n682), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT42), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n979), .A2(KEYINPUT42), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n975), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n974), .B(new_n983), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n972), .A2(new_n801), .ZN(new_n985));
  INV_X1    g0785(.A(new_n738), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n746), .B1(new_n209), .B2(new_n417), .C1(new_n986), .C2(new_n232), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n733), .ZN(new_n988));
  INV_X1    g0788(.A(new_n780), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n792), .A2(G68), .ZN(new_n990));
  INV_X1    g0790(.A(new_n775), .ZN(new_n991));
  INV_X1    g0791(.A(G150), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n990), .B1(new_n991), .B2(new_n835), .C1(new_n992), .C2(new_n773), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n989), .A2(G50), .B1(KEYINPUT107), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(G137), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n390), .B1(new_n995), .B2(new_n751), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n767), .A2(new_n752), .B1(new_n759), .B2(new_n317), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n996), .B(new_n997), .C1(G77), .C2(new_n757), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n994), .B(new_n998), .C1(KEYINPUT107), .C2(new_n993), .ZN(new_n999));
  XOR2_X1   g0799(.A(KEYINPUT106), .B(G317), .Z(new_n1000));
  OAI22_X1  g0800(.A1(new_n762), .A2(new_n424), .B1(new_n1000), .B2(new_n751), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n584), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n794), .A2(G116), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT46), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n773), .A2(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1001), .B(new_n1005), .C1(new_n1004), .C2(new_n1003), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n757), .A2(G97), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n767), .B2(new_n827), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n737), .B(new_n1008), .C1(G311), .C2(new_n775), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1006), .B(new_n1009), .C1(new_n823), .C2(new_n780), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n999), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT47), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n988), .B1(new_n1012), .B2(new_n745), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n967), .A2(new_n984), .B1(new_n985), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(G387));
  INV_X1    g0815(.A(new_n962), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n727), .A2(new_n961), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1016), .A2(new_n695), .A3(new_n1017), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1007), .B1(new_n992), .B2(new_n751), .C1(new_n777), .C2(new_n288), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G50), .B2(new_n774), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n762), .A2(new_n417), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G77), .B2(new_n794), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G159), .A2(new_n775), .B1(new_n766), .B2(new_n313), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1020), .A2(new_n737), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n780), .A2(new_n1002), .B1(new_n773), .B2(new_n1000), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1026), .A2(KEYINPUT109), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(KEYINPUT109), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n766), .A2(G311), .B1(new_n775), .B2(G322), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT110), .Z(new_n1030));
  NAND3_X1  g0830(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT48), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n762), .A2(new_n823), .B1(new_n759), .B2(new_n827), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1033), .A2(KEYINPUT49), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n757), .A2(G116), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n786), .A2(G326), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1036), .A2(new_n830), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(KEYINPUT49), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1024), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n820), .B1(new_n1041), .B2(KEYINPUT111), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(KEYINPUT111), .B2(new_n1041), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n680), .A2(new_n801), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n697), .A2(new_n694), .A3(new_n347), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n424), .B2(new_n694), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT108), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n229), .A2(new_n260), .ZN(new_n1048));
  AOI21_X1  g0848(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1049));
  AND3_X1   g0849(.A1(new_n313), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1050));
  AOI21_X1  g0850(.A(KEYINPUT50), .B1(new_n313), .B2(new_n202), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n697), .B(new_n1049), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n738), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1047), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n817), .B(new_n1044), .C1(new_n746), .C2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n961), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1043), .A2(new_n1055), .B1(new_n1056), .B2(new_n732), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1018), .A2(new_n1057), .ZN(G393));
  NAND2_X1  g0858(.A1(new_n964), .A2(new_n695), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT113), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n959), .A2(new_n963), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1060), .B1(new_n1061), .B2(new_n1016), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1060), .A3(new_n1016), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1059), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n959), .A2(new_n732), .A3(new_n963), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n780), .A2(new_n312), .B1(new_n202), .B2(new_n767), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT112), .Z(new_n1068));
  OAI22_X1  g0868(.A1(new_n752), .A2(new_n773), .B1(new_n991), .B2(new_n992), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n756), .A2(new_n511), .B1(new_n751), .B2(new_n835), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n762), .A2(new_n293), .B1(new_n759), .B2(new_n288), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n830), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1068), .A2(new_n1070), .A3(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n774), .A2(G311), .B1(G317), .B2(new_n775), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT52), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n762), .A2(new_n597), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n767), .A2(new_n1002), .B1(new_n759), .B2(new_n823), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n390), .B1(new_n786), .B2(G322), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(new_n424), .B2(new_n756), .C1(new_n777), .C2(new_n827), .ZN(new_n1080));
  OR4_X1    g0880(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n820), .B1(new_n1074), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n746), .B1(new_n450), .B2(new_n209), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n236), .B2(new_n738), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n1082), .A2(new_n817), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n801), .B2(new_n948), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1066), .A2(new_n1086), .ZN(new_n1087));
  OR3_X1    g0887(.A1(new_n1065), .A2(KEYINPUT114), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(KEYINPUT114), .B1(new_n1065), .B2(new_n1087), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(G390));
  OAI21_X1  g0890(.A(KEYINPUT100), .B1(new_n885), .B2(new_n889), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n897), .A2(new_n891), .A3(new_n898), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n909), .A2(new_n854), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n869), .A2(new_n884), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n808), .A2(new_n437), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n807), .B1(new_n709), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n908), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n854), .B(new_n1095), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1094), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n810), .B1(new_n926), .B2(new_n930), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n908), .A2(G330), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n725), .A2(new_n810), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n908), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1094), .A2(new_n1099), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1104), .A2(new_n732), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT115), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1104), .A2(KEYINPUT115), .A3(new_n732), .A4(new_n1107), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n439), .A2(G330), .A3(new_n931), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n922), .B(new_n1113), .C1(new_n668), .C2(new_n669), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(G330), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1098), .B1(new_n1116), .B2(new_n934), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1117), .A2(new_n1097), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1102), .B1(new_n1105), .B2(new_n908), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1118), .A2(new_n1106), .B1(new_n902), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1115), .A2(new_n1121), .A3(new_n1107), .A4(new_n1104), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1107), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1102), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1123), .A2(new_n1124), .B1(new_n1114), .B2(new_n1120), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1122), .A2(new_n695), .A3(new_n1125), .ZN(new_n1126));
  OR3_X1    g0926(.A1(new_n890), .A2(new_n899), .A3(new_n743), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n817), .B1(new_n312), .B2(new_n818), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n780), .A2(new_n1129), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n767), .A2(new_n995), .B1(new_n752), .B2(new_n762), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n756), .A2(new_n202), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n347), .B1(new_n786), .B2(G125), .ZN(new_n1134));
  INV_X1    g0934(.A(G128), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1134), .B1(new_n991), .B2(new_n1135), .C1(new_n832), .C2(new_n773), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n759), .A2(new_n992), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1137), .B(new_n1138), .Z(new_n1139));
  NOR4_X1   g0939(.A1(new_n1130), .A2(new_n1133), .A3(new_n1136), .A4(new_n1139), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n767), .A2(new_n424), .B1(new_n991), .B2(new_n823), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n989), .B2(G97), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT117), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n762), .A2(new_n293), .B1(new_n756), .B2(new_n288), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n347), .B1(new_n751), .B2(new_n827), .C1(new_n511), .C2(new_n759), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(G116), .C2(new_n774), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1140), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1127), .B(new_n1128), .C1(new_n820), .C2(new_n1147), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1112), .A2(new_n1126), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(G378));
  INV_X1    g0950(.A(KEYINPUT121), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1095), .A2(KEYINPUT40), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n907), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n906), .B(new_n903), .C1(new_n284), .C2(new_n305), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1101), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(G330), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n412), .A2(new_n415), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n413), .A2(new_n674), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  OR3_X1    g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1162), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n1156), .A2(new_n936), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1165), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n937), .B1(new_n911), .B2(new_n1155), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1116), .B1(new_n935), .B2(new_n938), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n900), .B(new_n913), .C1(new_n1166), .C2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1165), .B1(new_n1156), .B2(new_n936), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1168), .A2(new_n1169), .A3(new_n1167), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n854), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1172), .B(new_n1173), .C1(new_n1174), .C2(new_n912), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1151), .B1(new_n1171), .B2(new_n1175), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1175), .A2(new_n1151), .ZN(new_n1177));
  OAI21_X1  g0977(.A(KEYINPUT57), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1114), .B1(new_n1179), .B2(new_n1121), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n695), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT122), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT122), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(new_n695), .C1(new_n1178), .C2(new_n1180), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT57), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1185), .B1(new_n1180), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1182), .A2(new_n1184), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n830), .B2(new_n259), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n757), .A2(G58), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n293), .B2(new_n759), .C1(new_n823), .C2(new_n751), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1193), .A2(G41), .A3(new_n737), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT118), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n990), .B1(new_n991), .B2(new_n597), .C1(new_n450), .C2(new_n767), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n424), .A2(new_n773), .B1(new_n777), .B2(new_n417), .ZN(new_n1197));
  NOR3_X1   g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1191), .B1(new_n1198), .B2(KEYINPUT58), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G150), .A2(new_n792), .B1(new_n775), .B2(G125), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n832), .B2(new_n767), .C1(new_n759), .C2(new_n1129), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n1135), .A2(new_n773), .B1(new_n777), .B2(new_n995), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT59), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(KEYINPUT119), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n757), .A2(G159), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G33), .B(G41), .C1(new_n786), .C2(G124), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1205), .A2(KEYINPUT119), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1199), .B1(KEYINPUT58), .B2(new_n1198), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n745), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n817), .B1(new_n202), .B2(new_n818), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n1165), .C2(new_n743), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT120), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n1186), .B2(new_n732), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1189), .A2(new_n1216), .ZN(G375));
  NAND2_X1  g1017(.A1(new_n1098), .A2(new_n742), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n767), .A2(new_n597), .B1(new_n991), .B2(new_n827), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1021), .B1(G303), .B2(new_n786), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n823), .B2(new_n773), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(G97), .C2(new_n794), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n347), .B1(new_n756), .B2(new_n293), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT123), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1222), .B(new_n1224), .C1(new_n424), .C2(new_n780), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n767), .A2(new_n1129), .B1(new_n752), .B2(new_n759), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n991), .A2(new_n832), .B1(new_n202), .B2(new_n762), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1226), .A2(new_n1227), .A3(new_n830), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1192), .B1(new_n1135), .B2(new_n751), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G150), .B2(new_n790), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(new_n995), .C2(new_n773), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n820), .B1(new_n1225), .B2(new_n1231), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n817), .B(new_n1232), .C1(new_n288), .C2(new_n818), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1121), .A2(new_n732), .B1(new_n1218), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1114), .A2(new_n1120), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n966), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n1114), .B2(new_n1120), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1234), .B1(new_n1236), .B2(new_n1238), .ZN(G381));
  NAND3_X1  g1039(.A1(new_n1018), .A2(new_n805), .A3(new_n1057), .ZN(new_n1240));
  OR4_X1    g1040(.A1(G384), .A2(G387), .A3(G381), .A4(new_n1240), .ZN(new_n1241));
  OR4_X1    g1041(.A1(G390), .A2(new_n1241), .A3(G378), .A4(G375), .ZN(G407));
  NAND2_X1  g1042(.A1(new_n675), .A2(G213), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1149), .A2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G407), .B(G213), .C1(G375), .C2(new_n1245), .ZN(G409));
  NAND2_X1  g1046(.A1(G393), .A2(G396), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1247), .A2(new_n1240), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1088), .A2(new_n1089), .A3(new_n1014), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT126), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1014), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1248), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1252), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1248), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1254), .A2(new_n1250), .A3(new_n1255), .A4(new_n1249), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1189), .A2(G378), .A3(new_n1216), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1115), .B1(new_n1259), .B2(new_n1120), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(new_n1237), .A3(new_n1186), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n732), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n1214), .A3(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT124), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1149), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1149), .B2(new_n1263), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1258), .A2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT60), .B1(new_n1114), .B2(new_n1120), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1235), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1114), .A2(KEYINPUT60), .A3(new_n1120), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(new_n695), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1234), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n842), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1272), .A2(G384), .A3(new_n1234), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1268), .A2(new_n1243), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1244), .B1(new_n1258), .B2(new_n1267), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(KEYINPUT63), .A3(new_n1276), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1268), .A2(new_n1243), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1244), .A2(KEYINPUT125), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1274), .A2(new_n1275), .A3(new_n1283), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1244), .A2(G2897), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1284), .B(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT61), .B1(new_n1282), .B2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1257), .A2(new_n1279), .A3(new_n1281), .A4(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT61), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1280), .B2(new_n1286), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1277), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1280), .A2(KEYINPUT62), .A3(new_n1276), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1292), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT127), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1290), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1295), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT62), .B1(new_n1280), .B2(new_n1276), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1297), .B(new_n1288), .C1(new_n1299), .C2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1289), .B1(new_n1298), .B2(new_n1302), .ZN(G405));
  XNOR2_X1  g1103(.A(G375), .B(G378), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(new_n1304), .B(new_n1276), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1305), .B(new_n1257), .ZN(G402));
endmodule


