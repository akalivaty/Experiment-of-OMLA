//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927;
  INV_X1    g000(.A(G15gat), .ZN(new_n202));
  INV_X1    g001(.A(G22gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G15gat), .A2(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT90), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT90), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n208), .A3(new_n205), .ZN(new_n209));
  INV_X1    g008(.A(G1gat), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n207), .A2(new_n209), .B1(KEYINPUT16), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(G8gat), .B1(new_n211), .B2(KEYINPUT91), .ZN(new_n212));
  INV_X1    g011(.A(new_n209), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n208), .B1(new_n204), .B2(new_n205), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT16), .ZN(new_n215));
  OAI22_X1  g014(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(G1gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n207), .A2(new_n210), .A3(new_n209), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n212), .B(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(G43gat), .B(G50gat), .Z(new_n220));
  INV_X1    g019(.A(KEYINPUT15), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT86), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g024(.A(KEYINPUT86), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(G29gat), .A2(G36gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT14), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT87), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(KEYINPUT87), .A3(new_n229), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n227), .A2(KEYINPUT88), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G29gat), .A2(G36gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR4_X1   g035(.A1(new_n231), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT87), .B1(new_n228), .B2(new_n229), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT88), .B1(new_n239), .B2(new_n227), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n222), .B1(new_n236), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n242));
  INV_X1    g041(.A(new_n222), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n230), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n220), .A2(new_n221), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n235), .B(KEYINPUT89), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n243), .A2(new_n244), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n241), .A2(new_n242), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n242), .B1(new_n241), .B2(new_n247), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n219), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G229gat), .A2(G233gat), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n218), .B(G8gat), .C1(KEYINPUT91), .C2(new_n211), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT91), .ZN(new_n253));
  INV_X1    g052(.A(G8gat), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n216), .B(new_n217), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n247), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n250), .A2(new_n251), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT92), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(KEYINPUT18), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n257), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n219), .A2(new_n263), .A3(KEYINPUT93), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT93), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n265), .B1(new_n256), .B2(new_n257), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n266), .A3(new_n258), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n251), .B(KEYINPUT13), .Z(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n261), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n250), .A2(new_n251), .A3(new_n258), .A4(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n262), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(G113gat), .B(G141gat), .Z(new_n273));
  XNOR2_X1  g072(.A(G169gat), .B(G197gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT12), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n262), .A2(new_n269), .A3(new_n271), .A4(new_n278), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G230gat), .ZN(new_n284));
  INV_X1    g083(.A(G233gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G99gat), .A2(G106gat), .ZN(new_n287));
  INV_X1    g086(.A(G85gat), .ZN(new_n288));
  INV_X1    g087(.A(G92gat), .ZN(new_n289));
  AOI22_X1  g088(.A1(KEYINPUT8), .A2(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT7), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(new_n288), .B2(new_n289), .ZN(new_n292));
  NAND3_X1  g091(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G99gat), .B(G106gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G71gat), .A2(G78gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT94), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n298), .A2(G71gat), .A3(G78gat), .ZN(new_n299));
  INV_X1    g098(.A(G71gat), .ZN(new_n300));
  INV_X1    g099(.A(G78gat), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT94), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n297), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT95), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G64gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G57gat), .ZN(new_n307));
  INV_X1    g106(.A(G57gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G64gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT9), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n307), .A2(new_n309), .B1(new_n310), .B2(new_n297), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(G71gat), .A2(G78gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT94), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n298), .B1(G71gat), .B2(G78gat), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT95), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n305), .A2(new_n312), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT96), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n309), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n308), .A2(KEYINPUT96), .A3(G64gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n307), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n300), .A2(new_n301), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n297), .B1(new_n323), .B2(new_n310), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n318), .A2(KEYINPUT100), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT100), .B1(new_n318), .B2(new_n325), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n296), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT10), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n318), .A2(KEYINPUT100), .A3(new_n325), .ZN(new_n330));
  INV_X1    g129(.A(new_n296), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n328), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT98), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n296), .B(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n325), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n316), .A2(KEYINPUT95), .ZN(new_n337));
  AOI211_X1 g136(.A(new_n304), .B(new_n313), .C1(new_n314), .C2(new_n315), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n336), .B1(new_n339), .B2(new_n312), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(KEYINPUT10), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n286), .B1(new_n333), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n286), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n328), .B2(new_n332), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G120gat), .B(G148gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(G204gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(KEYINPUT101), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(G176gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n345), .B(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n283), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT35), .ZN(new_n353));
  INV_X1    g152(.A(G227gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(new_n285), .ZN(new_n355));
  INV_X1    g154(.A(G169gat), .ZN(new_n356));
  INV_X1    g155(.A(G176gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT23), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT64), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n363), .A2(new_n364), .B1(new_n362), .B2(new_n361), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT25), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n358), .B1(KEYINPUT23), .B2(new_n360), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n366), .B1(new_n367), .B2(KEYINPUT64), .ZN(new_n368));
  INV_X1    g167(.A(G183gat), .ZN(new_n369));
  INV_X1    g168(.A(G190gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(KEYINPUT24), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(KEYINPUT24), .B2(new_n372), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT65), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n373), .B(KEYINPUT65), .C1(KEYINPUT24), .C2(new_n372), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n365), .A2(new_n368), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n367), .B1(KEYINPUT23), .B2(new_n360), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n366), .B1(new_n379), .B2(new_n374), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G134gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(KEYINPUT68), .ZN(new_n383));
  XNOR2_X1  g182(.A(G113gat), .B(G120gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(KEYINPUT1), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT1), .ZN(new_n386));
  INV_X1    g185(.A(G113gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n387), .A2(G120gat), .ZN(new_n388));
  INV_X1    g187(.A(G120gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(G113gat), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n386), .B(new_n382), .C1(new_n388), .C2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G127gat), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n385), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n392), .B1(new_n385), .B2(new_n391), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT69), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n372), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n358), .A2(KEYINPUT26), .A3(new_n360), .ZN(new_n398));
  AOI211_X1 g197(.A(new_n397), .B(new_n398), .C1(KEYINPUT26), .C2(new_n360), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT67), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT27), .B(G183gat), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n401), .A2(KEYINPUT28), .A3(new_n370), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT27), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT66), .B1(new_n403), .B2(G183gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n370), .ZN(new_n405));
  INV_X1    g204(.A(new_n401), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT66), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n402), .B1(new_n408), .B2(KEYINPUT28), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n399), .A2(new_n400), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n400), .B1(new_n399), .B2(new_n409), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n381), .B(new_n396), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n399), .A2(new_n409), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT67), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n400), .A3(new_n409), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n414), .A2(new_n415), .B1(new_n380), .B2(new_n378), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n393), .A2(new_n394), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT69), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n355), .B(new_n412), .C1(new_n416), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT70), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n381), .B1(new_n410), .B2(new_n411), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n417), .A2(KEYINPUT69), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(new_n396), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT70), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n424), .A2(new_n425), .A3(new_n355), .A4(new_n412), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT32), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n355), .B1(new_n424), .B2(new_n412), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT34), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI211_X1 g230(.A(KEYINPUT34), .B(new_n355), .C1(new_n424), .C2(new_n412), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n427), .B(KEYINPUT32), .C1(new_n431), .C2(new_n432), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G15gat), .B(G43gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(G71gat), .B(G99gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n437), .B(new_n438), .Z(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n440), .B1(new_n427), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n436), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT29), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT79), .ZN(new_n446));
  NAND2_X1  g245(.A1(G155gat), .A2(G162gat), .ZN(new_n447));
  INV_X1    g246(.A(G155gat), .ZN(new_n448));
  INV_X1    g247(.A(G162gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(KEYINPUT77), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g250(.A(G141gat), .B(G148gat), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n447), .B(new_n450), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n447), .B1(new_n450), .B2(KEYINPUT2), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT78), .ZN(new_n455));
  INV_X1    g254(.A(G141gat), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n455), .B1(new_n456), .B2(G148gat), .ZN(new_n457));
  INV_X1    g256(.A(G148gat), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(KEYINPUT78), .A3(G141gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n458), .A2(G141gat), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n454), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n453), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n446), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n463), .A2(new_n446), .A3(KEYINPUT3), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n445), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT71), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n468), .A2(KEYINPUT22), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(KEYINPUT22), .ZN(new_n470));
  INV_X1    g269(.A(G211gat), .ZN(new_n471));
  INV_X1    g270(.A(G218gat), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n469), .B(new_n470), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G197gat), .B(G204gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  XOR2_X1   g274(.A(G211gat), .B(G218gat), .Z(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT72), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n475), .B(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n467), .A2(new_n478), .ZN(new_n479));
  AND2_X1   g278(.A1(G228gat), .A2(G233gat), .ZN(new_n480));
  INV_X1    g279(.A(new_n463), .ZN(new_n481));
  INV_X1    g280(.A(new_n478), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT3), .B1(new_n482), .B2(new_n445), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n479), .B(new_n480), .C1(new_n481), .C2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n475), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT29), .B1(new_n485), .B2(new_n476), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(new_n476), .B2(new_n485), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT3), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n481), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n489), .B1(new_n467), .B2(new_n478), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n484), .B1(new_n480), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G78gat), .B(G106gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT31), .B(G50gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT84), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n495), .A3(G22gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(G22gat), .B2(new_n494), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n491), .B(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n434), .A2(new_n442), .A3(new_n435), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n444), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G225gat), .A2(G233gat), .ZN(new_n502));
  XOR2_X1   g301(.A(new_n502), .B(KEYINPUT80), .Z(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n417), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n481), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n417), .A2(new_n463), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT83), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT83), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n417), .B(new_n481), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n512), .B(new_n509), .C1(new_n513), .C2(new_n504), .ZN(new_n514));
  OAI221_X1 g313(.A(new_n417), .B1(new_n488), .B2(new_n481), .C1(new_n465), .C2(new_n466), .ZN(new_n515));
  OR3_X1    g314(.A1(new_n417), .A2(KEYINPUT4), .A3(new_n463), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n515), .B(new_n504), .C1(KEYINPUT81), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n518), .A2(KEYINPUT81), .A3(new_n516), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n511), .B(new_n514), .C1(new_n517), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n516), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n521), .A2(new_n515), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n522), .A2(new_n504), .A3(new_n510), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT0), .B(G57gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(G85gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G1gat), .B(G29gat), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n526), .B(new_n527), .Z(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n520), .A2(new_n523), .A3(new_n528), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n524), .A2(KEYINPUT6), .A3(new_n529), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G64gat), .B(G92gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(G36gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT74), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(new_n254), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT76), .ZN(new_n540));
  NAND2_X1  g339(.A1(G226gat), .A2(G233gat), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n541), .B(KEYINPUT73), .Z(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n421), .A2(new_n445), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n378), .A2(new_n380), .B1(new_n399), .B2(new_n409), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n542), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n482), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n421), .A2(new_n542), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n543), .B1(new_n545), .B2(KEYINPUT29), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n478), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI221_X1 g349(.A(new_n539), .B1(new_n540), .B2(KEYINPUT30), .C1(new_n547), .C2(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT76), .B(KEYINPUT30), .Z(new_n552));
  NOR2_X1   g351(.A1(new_n547), .A2(new_n550), .ZN(new_n553));
  INV_X1    g352(.A(new_n539), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT75), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n556), .B1(new_n553), .B2(new_n554), .ZN(new_n557));
  NOR4_X1   g356(.A1(new_n547), .A2(new_n550), .A3(KEYINPUT75), .A4(new_n539), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n551), .B(new_n555), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n535), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n353), .B1(new_n501), .B2(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n434), .A2(new_n442), .A3(new_n435), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n442), .B1(new_n434), .B2(new_n435), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n559), .B1(new_n534), .B2(new_n533), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT35), .A4(new_n499), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n563), .B2(new_n564), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n444), .A2(KEYINPUT36), .A3(new_n500), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n513), .A2(new_n504), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n573), .B(KEYINPUT39), .C1(new_n522), .C2(new_n504), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n504), .B1(new_n521), .B2(new_n515), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT39), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n529), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n574), .A2(KEYINPUT40), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT40), .B1(new_n574), .B2(new_n577), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(new_n559), .A3(new_n530), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n553), .A2(KEYINPUT37), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n544), .A2(new_n482), .A3(new_n546), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n548), .A2(new_n478), .A3(new_n549), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(KEYINPUT37), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n554), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT38), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n553), .B2(KEYINPUT37), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n586), .A2(new_n587), .B1(new_n582), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n553), .A2(new_n587), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(new_n539), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n533), .A2(new_n534), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n581), .B(new_n499), .C1(new_n589), .C2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n561), .A2(new_n498), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n572), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n352), .B1(new_n568), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G127gat), .B(G155gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(G211gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n340), .A2(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n219), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(new_n369), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT97), .B(KEYINPUT21), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n340), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n601), .A2(new_n603), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n598), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n601), .A2(new_n603), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n601), .A2(new_n603), .ZN(new_n608));
  INV_X1    g407(.A(new_n598), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n606), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n606), .B2(new_n610), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n618));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n622), .B(KEYINPUT99), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n248), .A2(new_n249), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n296), .B(KEYINPUT98), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n335), .A2(new_n257), .ZN(new_n629));
  AND4_X1   g428(.A1(new_n624), .A2(new_n627), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n625), .A2(new_n626), .B1(KEYINPUT41), .B2(new_n617), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n624), .B1(new_n631), .B2(new_n629), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n621), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n623), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n631), .A2(new_n624), .A3(new_n629), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(new_n620), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n616), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n596), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n535), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(new_n210), .ZN(G1324gat));
  INV_X1    g442(.A(new_n641), .ZN(new_n644));
  NAND2_X1  g443(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n215), .A2(new_n254), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n644), .A2(new_n559), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT42), .ZN(new_n648));
  OR3_X1    g447(.A1(new_n647), .A2(KEYINPUT102), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n254), .B1(new_n644), .B2(new_n559), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(new_n648), .B2(new_n647), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT102), .B1(new_n647), .B2(new_n648), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(G1325gat));
  NOR3_X1   g452(.A1(new_n641), .A2(new_n202), .A3(new_n572), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n644), .A2(new_n565), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n654), .B1(new_n202), .B2(new_n655), .ZN(G1326gat));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n499), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT43), .B(G22gat), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1327gat));
  AOI21_X1  g458(.A(new_n638), .B1(new_n568), .B2(new_n595), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n614), .A2(new_n615), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n352), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n663), .A2(G29gat), .A3(new_n535), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT45), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n572), .A2(new_n593), .A3(new_n594), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n562), .A2(new_n567), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n639), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI211_X1 g472(.A(KEYINPUT44), .B(new_n639), .C1(new_n669), .C2(new_n670), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n662), .ZN(new_n676));
  OR3_X1    g475(.A1(new_n676), .A2(KEYINPUT104), .A3(new_n535), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT104), .B1(new_n676), .B2(new_n535), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n677), .A2(G29gat), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n666), .A2(new_n667), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n668), .A2(new_n679), .A3(new_n680), .ZN(G1328gat));
  OR3_X1    g480(.A1(new_n663), .A2(G36gat), .A3(new_n560), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(KEYINPUT46), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(KEYINPUT46), .ZN(new_n686));
  OAI21_X1  g485(.A(G36gat), .B1(new_n676), .B2(new_n560), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(G1329gat));
  INV_X1    g487(.A(new_n565), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n663), .A2(G43gat), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n572), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n673), .A2(new_n692), .A3(new_n662), .A4(new_n674), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G43gat), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n691), .A2(new_n694), .A3(KEYINPUT47), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n694), .A2(KEYINPUT107), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n694), .A2(KEYINPUT107), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n696), .A2(new_n697), .A3(new_n690), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n699));
  OAI21_X1  g498(.A(new_n695), .B1(new_n698), .B2(new_n699), .ZN(G1330gat));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT48), .ZN(new_n702));
  OAI21_X1  g501(.A(G50gat), .B1(new_n676), .B2(new_n499), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n663), .A2(G50gat), .A3(new_n499), .ZN(new_n704));
  AOI211_X1 g503(.A(new_n701), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n701), .A2(new_n702), .ZN(new_n707));
  AND4_X1   g506(.A1(new_n706), .A2(new_n703), .A3(new_n707), .A4(new_n704), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n705), .A2(new_n708), .ZN(G1331gat));
  NAND2_X1  g508(.A1(new_n640), .A2(new_n283), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(new_n568), .B2(new_n595), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n350), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n535), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(new_n308), .ZN(G1332gat));
  AOI211_X1 g513(.A(new_n560), .B(new_n712), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1333gat));
  OAI21_X1  g516(.A(new_n300), .B1(new_n712), .B2(new_n689), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n711), .A2(G71gat), .A3(new_n350), .A4(new_n692), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g520(.A1(new_n712), .A2(new_n499), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT109), .B(G78gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1335gat));
  INV_X1    g523(.A(new_n535), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n661), .A2(new_n282), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n673), .A2(new_n350), .A3(new_n674), .A4(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n725), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT111), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT111), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n733), .B(new_n725), .C1(new_n729), .C2(new_n730), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n732), .A2(G85gat), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT112), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n726), .B1(new_n660), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n671), .A2(KEYINPUT112), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT51), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n660), .A2(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n671), .A2(KEYINPUT112), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .A4(new_n726), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n744), .A2(new_n288), .A3(new_n725), .A4(new_n350), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n735), .A2(new_n745), .ZN(G1336gat));
  NOR2_X1   g545(.A1(new_n560), .A2(G92gat), .ZN(new_n747));
  AND4_X1   g546(.A1(new_n350), .A2(new_n739), .A3(new_n743), .A4(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n559), .B1(new_n729), .B2(new_n730), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(G92gat), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751));
  OAI21_X1  g550(.A(G92gat), .B1(new_n727), .B2(new_n560), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n751), .ZN(new_n753));
  OAI22_X1  g552(.A1(new_n750), .A2(new_n751), .B1(new_n748), .B2(new_n753), .ZN(G1337gat));
  NOR2_X1   g553(.A1(new_n729), .A2(new_n730), .ZN(new_n755));
  OAI21_X1  g554(.A(G99gat), .B1(new_n755), .B2(new_n572), .ZN(new_n756));
  INV_X1    g555(.A(G99gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n744), .A2(new_n757), .A3(new_n350), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n756), .B1(new_n689), .B2(new_n758), .ZN(G1338gat));
  NOR2_X1   g558(.A1(new_n499), .A2(G106gat), .ZN(new_n760));
  AND4_X1   g559(.A1(new_n350), .A2(new_n739), .A3(new_n743), .A4(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n498), .B1(new_n729), .B2(new_n730), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(G106gat), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764));
  OAI21_X1  g563(.A(G106gat), .B1(new_n727), .B2(new_n499), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n764), .ZN(new_n766));
  OAI22_X1  g565(.A1(new_n763), .A2(new_n764), .B1(new_n761), .B2(new_n766), .ZN(G1339gat));
  INV_X1    g566(.A(KEYINPUT100), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n337), .A2(new_n338), .A3(new_n311), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n769), .B2(new_n336), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n331), .B1(new_n770), .B2(new_n330), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n296), .B1(new_n340), .B2(KEYINPUT100), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n771), .A2(KEYINPUT10), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n340), .A2(KEYINPUT10), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n626), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n343), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n333), .A2(new_n286), .A3(new_n341), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(KEYINPUT54), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n349), .B1(new_n342), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n778), .A2(new_n780), .A3(KEYINPUT55), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n345), .A2(new_n349), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n778), .A2(new_n780), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n783), .A2(new_n282), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n267), .A2(new_n268), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n251), .B1(new_n250), .B2(new_n258), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n277), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n350), .A2(new_n790), .A3(new_n281), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n639), .B1(new_n787), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n786), .A2(new_n281), .A3(new_n790), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n781), .A2(new_n782), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n793), .A2(new_n638), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n616), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n350), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n661), .A2(new_n638), .A3(new_n797), .A4(new_n283), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n501), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n535), .A2(new_n559), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n283), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(new_n387), .ZN(G1340gat));
  NOR2_X1   g602(.A1(new_n801), .A2(new_n797), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(new_n389), .ZN(G1341gat));
  NOR2_X1   g604(.A1(new_n801), .A2(new_n616), .ZN(new_n806));
  XNOR2_X1  g605(.A(KEYINPUT68), .B(G127gat), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n806), .B(new_n807), .ZN(G1342gat));
  NAND3_X1  g607(.A1(new_n799), .A2(new_n639), .A3(new_n800), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(G134gat), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n812), .A2(KEYINPUT113), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(KEYINPUT113), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n811), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n809), .A2(G134gat), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n813), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(G1343gat));
  AND2_X1   g616(.A1(new_n572), .A2(new_n800), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n796), .A2(new_n798), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n820), .A3(new_n498), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n786), .A2(KEYINPUT114), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n784), .A2(new_n823), .A3(new_n785), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n822), .A2(new_n783), .A3(new_n282), .A4(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n639), .B1(new_n825), .B2(new_n791), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n616), .B1(new_n826), .B2(new_n795), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n499), .B1(new_n827), .B2(new_n798), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n818), .B(new_n821), .C1(new_n828), .C2(new_n820), .ZN(new_n829));
  OAI21_X1  g628(.A(G141gat), .B1(new_n829), .B2(new_n283), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n692), .A2(new_n499), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n831), .A2(new_n800), .A3(new_n819), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(new_n456), .A3(new_n282), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g634(.A1(new_n832), .A2(new_n458), .A3(new_n350), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n829), .A2(new_n797), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(new_n838), .A3(G148gat), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT115), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n827), .A2(new_n841), .A3(new_n798), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n827), .B2(new_n798), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT57), .B1(new_n844), .B2(new_n498), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n820), .B1(new_n796), .B2(new_n798), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n498), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n846), .A2(KEYINPUT116), .A3(new_n498), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n350), .B(new_n818), .C1(new_n845), .C2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n838), .B1(new_n852), .B2(G148gat), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n836), .B1(new_n840), .B2(new_n853), .ZN(G1345gat));
  AOI21_X1  g653(.A(G155gat), .B1(new_n832), .B2(new_n661), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n829), .A2(new_n448), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n661), .ZN(G1346gat));
  AOI21_X1  g656(.A(G162gat), .B1(new_n832), .B2(new_n639), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n829), .A2(new_n449), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(new_n639), .ZN(G1347gat));
  AOI211_X1 g659(.A(new_n725), .B(new_n560), .C1(new_n796), .C2(new_n798), .ZN(new_n861));
  INV_X1    g660(.A(new_n501), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n283), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(new_n356), .ZN(G1348gat));
  NOR2_X1   g664(.A1(new_n863), .A2(new_n797), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(new_n357), .ZN(G1349gat));
  NAND3_X1  g666(.A1(new_n861), .A2(new_n661), .A3(new_n862), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n868), .A2(new_n401), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT60), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT118), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n868), .A2(new_n369), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n869), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI211_X1 g672(.A(KEYINPUT119), .B(new_n871), .C1(new_n869), .C2(new_n872), .ZN(new_n874));
  AOI211_X1 g673(.A(new_n873), .B(new_n874), .C1(KEYINPUT119), .C2(new_n870), .ZN(G1350gat));
  NAND3_X1  g674(.A1(new_n861), .A2(new_n639), .A3(new_n862), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(G190gat), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT120), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(G190gat), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT61), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1351gat));
  AND2_X1   g680(.A1(new_n861), .A2(new_n831), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n883), .A2(G197gat), .A3(new_n283), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n572), .A2(new_n535), .A3(new_n559), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n885), .B(KEYINPUT121), .Z(new_n886));
  NAND2_X1  g685(.A1(new_n822), .A2(new_n824), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n282), .A2(new_n782), .A3(new_n781), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n791), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n795), .B1(new_n889), .B2(new_n638), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n798), .B1(new_n890), .B2(new_n661), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT117), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n827), .A2(new_n841), .A3(new_n798), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n498), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n820), .ZN(new_n895));
  AND4_X1   g694(.A1(KEYINPUT116), .A2(new_n819), .A3(KEYINPUT57), .A4(new_n498), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT116), .B1(new_n846), .B2(new_n498), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n886), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n282), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n884), .B1(new_n900), .B2(G197gat), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n901), .B(new_n902), .ZN(G1352gat));
  XOR2_X1   g702(.A(KEYINPUT123), .B(G204gat), .Z(new_n904));
  NAND2_X1  g703(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n882), .A2(new_n350), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n906), .B(new_n907), .ZN(new_n908));
  AOI211_X1 g707(.A(new_n797), .B(new_n886), .C1(new_n895), .C2(new_n898), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n904), .B2(new_n909), .ZN(G1353gat));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n471), .B1(new_n899), .B2(new_n661), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(KEYINPUT63), .ZN(new_n913));
  INV_X1    g712(.A(new_n886), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n661), .B(new_n914), .C1(new_n845), .C2(new_n851), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n915), .A2(KEYINPUT125), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT63), .ZN(new_n920));
  AOI211_X1 g719(.A(new_n616), .B(new_n886), .C1(new_n895), .C2(new_n898), .ZN(new_n921));
  OAI211_X1 g720(.A(KEYINPUT126), .B(new_n920), .C1(new_n921), .C2(new_n471), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n913), .A2(new_n918), .A3(new_n919), .A4(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n882), .A2(new_n471), .A3(new_n661), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1354gat));
  NAND3_X1  g724(.A1(new_n882), .A2(new_n472), .A3(new_n639), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n899), .A2(new_n639), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n927), .B2(new_n472), .ZN(G1355gat));
endmodule


