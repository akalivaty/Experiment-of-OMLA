

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788;

  BUF_X1 U373 ( .A(n658), .Z(n723) );
  INV_X1 U374 ( .A(n625), .ZN(n354) );
  XNOR2_X1 U375 ( .A(n588), .B(n587), .ZN(n624) );
  XNOR2_X1 U376 ( .A(n520), .B(n521), .ZN(n770) );
  XNOR2_X1 U377 ( .A(n372), .B(G107), .ZN(n562) );
  XNOR2_X1 U378 ( .A(G119), .B(G128), .ZN(n522) );
  INV_X1 U379 ( .A(G116), .ZN(n372) );
  XNOR2_X1 U380 ( .A(n353), .B(n770), .ZN(n662) );
  XNOR2_X1 U381 ( .A(n528), .B(n527), .ZN(n353) );
  AND2_X2 U382 ( .A1(n650), .A2(n438), .ZN(n603) );
  XNOR2_X2 U383 ( .A(n580), .B(KEYINPUT40), .ZN(n787) );
  XNOR2_X2 U384 ( .A(n534), .B(n533), .ZN(n650) );
  INV_X1 U385 ( .A(n418), .ZN(n647) );
  NAND2_X1 U386 ( .A1(n418), .A2(n417), .ZN(n628) );
  XNOR2_X2 U387 ( .A(n626), .B(n354), .ZN(n418) );
  INV_X2 U388 ( .A(KEYINPUT66), .ZN(n470) );
  XNOR2_X1 U389 ( .A(G137), .B(G116), .ZN(n497) );
  AND2_X2 U390 ( .A1(n477), .A2(n473), .ZN(n472) );
  XNOR2_X2 U391 ( .A(G110), .B(KEYINPUT23), .ZN(n523) );
  XNOR2_X2 U392 ( .A(n697), .B(n602), .ZN(n636) );
  NOR2_X2 U393 ( .A1(n457), .A2(n455), .ZN(n454) );
  INV_X2 U394 ( .A(G953), .ZN(n778) );
  XNOR2_X1 U395 ( .A(n612), .B(KEYINPUT48), .ZN(n387) );
  AND2_X1 U396 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U397 ( .A1(n474), .A2(n686), .ZN(n473) );
  AND2_X1 U398 ( .A1(n446), .A2(n447), .ZN(n445) );
  NOR2_X2 U399 ( .A1(n594), .A2(n707), .ZN(n577) );
  XNOR2_X1 U400 ( .A(n608), .B(n441), .ZN(n442) );
  XNOR2_X1 U401 ( .A(n519), .B(n518), .ZN(n693) );
  AND2_X1 U402 ( .A1(n406), .A2(n404), .ZN(n403) );
  AND2_X1 U403 ( .A1(n401), .A2(KEYINPUT80), .ZN(n369) );
  XNOR2_X1 U404 ( .A(n454), .B(KEYINPUT32), .ZN(n783) );
  NAND2_X1 U405 ( .A1(n652), .A2(n651), .ZN(n667) );
  NOR2_X1 U406 ( .A1(n712), .A2(n649), .ZN(n654) );
  NAND2_X1 U407 ( .A1(n445), .A2(n443), .ZN(n638) );
  AND2_X1 U408 ( .A1(n609), .A2(n784), .ZN(n610) );
  NAND2_X1 U409 ( .A1(n444), .A2(n448), .ZN(n443) );
  NAND2_X1 U410 ( .A1(n442), .A2(n633), .ZN(n635) );
  AND2_X1 U411 ( .A1(n644), .A2(n392), .ZN(n391) );
  XNOR2_X1 U412 ( .A(n390), .B(n389), .ZN(n388) );
  OR2_X1 U413 ( .A1(n395), .A2(n394), .ZN(n355) );
  XNOR2_X1 U414 ( .A(n386), .B(n483), .ZN(n510) );
  INV_X1 U415 ( .A(n693), .ZN(n439) );
  XNOR2_X1 U416 ( .A(n370), .B(G101), .ZN(n539) );
  XNOR2_X1 U417 ( .A(n416), .B(n415), .ZN(n542) );
  BUF_X1 U418 ( .A(n646), .Z(n356) );
  NOR2_X1 U419 ( .A1(n654), .A2(n653), .ZN(n488) );
  NOR2_X2 U420 ( .A1(n624), .A2(n623), .ZN(n626) );
  XNOR2_X2 U421 ( .A(G146), .B(G125), .ZN(n543) );
  XNOR2_X1 U422 ( .A(n450), .B(G104), .ZN(n550) );
  XNOR2_X1 U423 ( .A(G113), .B(G122), .ZN(n450) );
  NAND2_X1 U424 ( .A1(n510), .A2(n381), .ZN(n375) );
  OR2_X2 U425 ( .A1(n395), .A2(n394), .ZN(n608) );
  NAND2_X1 U426 ( .A1(n396), .A2(n398), .ZN(n395) );
  NAND2_X1 U427 ( .A1(n509), .A2(n378), .ZN(n397) );
  XNOR2_X1 U428 ( .A(n469), .B(n541), .ZN(n764) );
  XNOR2_X1 U429 ( .A(n419), .B(n542), .ZN(n469) );
  XNOR2_X1 U430 ( .A(n562), .B(n420), .ZN(n419) );
  OR2_X1 U431 ( .A1(n681), .A2(n683), .ZN(n585) );
  INV_X1 U432 ( .A(KEYINPUT68), .ZN(n415) );
  XNOR2_X1 U433 ( .A(G119), .B(KEYINPUT3), .ZN(n416) );
  XNOR2_X1 U434 ( .A(n543), .B(KEYINPUT10), .ZN(n549) );
  XNOR2_X1 U435 ( .A(n550), .B(n360), .ZN(n436) );
  XNOR2_X1 U436 ( .A(G143), .B(G140), .ZN(n553) );
  XOR2_X1 U437 ( .A(KEYINPUT11), .B(KEYINPUT95), .Z(n554) );
  INV_X1 U438 ( .A(KEYINPUT65), .ZN(n370) );
  XNOR2_X1 U439 ( .A(n453), .B(n451), .ZN(n537) );
  XNOR2_X1 U440 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n453) );
  NOR2_X1 U441 ( .A1(n452), .A2(G953), .ZN(n451) );
  INV_X1 U442 ( .A(G224), .ZN(n452) );
  INV_X1 U443 ( .A(KEYINPUT4), .ZN(n494) );
  NOR2_X1 U444 ( .A1(n616), .A2(n571), .ZN(n481) );
  XNOR2_X1 U445 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U446 ( .A(n559), .B(n374), .ZN(n578) );
  XNOR2_X1 U447 ( .A(n558), .B(G475), .ZN(n374) );
  OR2_X2 U448 ( .A1(n379), .A2(n376), .ZN(n697) );
  NAND2_X1 U449 ( .A1(n375), .A2(n380), .ZN(n379) );
  NAND2_X1 U450 ( .A1(n381), .A2(G902), .ZN(n380) );
  INV_X1 U451 ( .A(KEYINPUT1), .ZN(n441) );
  XOR2_X1 U452 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n501) );
  XOR2_X1 U453 ( .A(KEYINPUT5), .B(G113), .Z(n498) );
  XNOR2_X1 U454 ( .A(G134), .B(G122), .ZN(n560) );
  XOR2_X1 U455 ( .A(KEYINPUT98), .B(KEYINPUT9), .Z(n561) );
  XNOR2_X1 U456 ( .A(n540), .B(n361), .ZN(n421) );
  INV_X1 U457 ( .A(n578), .ZN(n592) );
  BUF_X1 U458 ( .A(n697), .Z(n424) );
  XNOR2_X1 U459 ( .A(n741), .B(n365), .ZN(n486) );
  XNOR2_X1 U460 ( .A(n371), .B(KEYINPUT20), .ZN(n530) );
  NAND2_X1 U461 ( .A1(n517), .A2(G234), .ZN(n371) );
  NAND2_X1 U462 ( .A1(n476), .A2(n475), .ZN(n474) );
  INV_X1 U463 ( .A(KEYINPUT79), .ZN(n475) );
  AND2_X1 U464 ( .A1(n687), .A2(KEYINPUT79), .ZN(n478) );
  NOR2_X1 U465 ( .A1(G902), .A2(G237), .ZN(n544) );
  NAND2_X1 U466 ( .A1(n399), .A2(G902), .ZN(n398) );
  NAND2_X1 U467 ( .A1(n511), .A2(n378), .ZN(n377) );
  NOR2_X1 U468 ( .A1(G953), .A2(G237), .ZN(n551) );
  INV_X1 U469 ( .A(KEYINPUT16), .ZN(n420) );
  XNOR2_X1 U470 ( .A(KEYINPUT77), .B(KEYINPUT24), .ZN(n368) );
  XNOR2_X1 U471 ( .A(n513), .B(n512), .ZN(n514) );
  NAND2_X1 U472 ( .A1(G234), .A2(G237), .ZN(n512) );
  XOR2_X1 U473 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n513) );
  XNOR2_X1 U474 ( .A(n515), .B(n427), .ZN(n426) );
  INV_X1 U475 ( .A(KEYINPUT105), .ZN(n427) );
  NAND2_X1 U476 ( .A1(n697), .A2(n710), .ZN(n390) );
  INV_X1 U477 ( .A(KEYINPUT30), .ZN(n389) );
  XNOR2_X1 U478 ( .A(n549), .B(n436), .ZN(n557) );
  XOR2_X1 U479 ( .A(G902), .B(KEYINPUT15), .Z(n657) );
  XNOR2_X1 U480 ( .A(n764), .B(n412), .ZN(n740) );
  AND2_X1 U481 ( .A1(n363), .A2(n435), .ZN(n384) );
  NOR2_X1 U482 ( .A1(n357), .A2(n449), .ZN(n447) );
  INV_X1 U483 ( .A(n637), .ZN(n449) );
  NOR2_X1 U484 ( .A1(n647), .A2(KEYINPUT34), .ZN(n448) );
  XNOR2_X1 U485 ( .A(n579), .B(KEYINPUT100), .ZN(n605) );
  NAND2_X1 U486 ( .A1(n578), .A2(n591), .ZN(n579) );
  NOR2_X2 U487 ( .A1(n689), .A2(n355), .ZN(n644) );
  XNOR2_X1 U488 ( .A(n504), .B(n499), .ZN(n483) );
  XNOR2_X1 U489 ( .A(n411), .B(n565), .ZN(n751) );
  XNOR2_X1 U490 ( .A(n567), .B(n358), .ZN(n411) );
  XOR2_X1 U491 ( .A(KEYINPUT97), .B(KEYINPUT7), .Z(n564) );
  XNOR2_X1 U492 ( .A(G104), .B(G107), .ZN(n505) );
  XNOR2_X1 U493 ( .A(n421), .B(n521), .ZN(n506) );
  XNOR2_X1 U494 ( .A(n382), .B(KEYINPUT110), .ZN(n784) );
  NAND2_X1 U495 ( .A1(n479), .A2(n383), .ZN(n382) );
  NAND2_X1 U496 ( .A1(n480), .A2(KEYINPUT36), .ZN(n479) );
  AND2_X1 U497 ( .A1(n385), .A2(n384), .ZN(n383) );
  NAND2_X1 U498 ( .A1(n435), .A2(n456), .ZN(n455) );
  XNOR2_X1 U499 ( .A(n648), .B(n373), .ZN(n684) );
  XNOR2_X1 U500 ( .A(n413), .B(KEYINPUT94), .ZN(n373) );
  INV_X1 U501 ( .A(KEYINPUT31), .ZN(n413) );
  XNOR2_X1 U502 ( .A(KEYINPUT101), .B(n584), .ZN(n683) );
  INV_X1 U503 ( .A(n664), .ZN(n433) );
  INV_X1 U504 ( .A(KEYINPUT60), .ZN(n463) );
  INV_X1 U505 ( .A(KEYINPUT56), .ZN(n428) );
  INV_X1 U506 ( .A(n435), .ZN(n690) );
  BUF_X1 U507 ( .A(n442), .Z(n435) );
  AND2_X1 U508 ( .A1(n647), .A2(KEYINPUT34), .ZN(n357) );
  XOR2_X1 U509 ( .A(n561), .B(n560), .Z(n358) );
  XOR2_X1 U510 ( .A(n554), .B(n553), .Z(n359) );
  INV_X1 U511 ( .A(n509), .ZN(n399) );
  XNOR2_X1 U512 ( .A(n508), .B(G469), .ZN(n509) );
  INV_X1 U513 ( .A(G902), .ZN(n378) );
  AND2_X1 U514 ( .A1(G214), .A2(n551), .ZN(n360) );
  AND2_X1 U515 ( .A1(n778), .A2(G227), .ZN(n361) );
  AND2_X1 U516 ( .A1(n481), .A2(n482), .ZN(n362) );
  OR2_X1 U517 ( .A1(n481), .A2(n482), .ZN(n363) );
  XOR2_X1 U518 ( .A(KEYINPUT84), .B(KEYINPUT33), .Z(n364) );
  INV_X1 U519 ( .A(KEYINPUT36), .ZN(n482) );
  XOR2_X1 U520 ( .A(n743), .B(n742), .Z(n365) );
  XOR2_X1 U521 ( .A(n750), .B(n749), .Z(n366) );
  XOR2_X1 U522 ( .A(n510), .B(KEYINPUT62), .Z(n367) );
  INV_X1 U523 ( .A(n756), .ZN(n484) );
  NOR2_X1 U524 ( .A1(n600), .A2(n599), .ZN(n611) );
  NAND2_X1 U525 ( .A1(n403), .A2(n400), .ZN(n462) );
  NAND2_X1 U526 ( .A1(n408), .A2(n488), .ZN(n407) );
  NAND2_X1 U527 ( .A1(n462), .A2(n459), .ZN(n458) );
  NAND2_X1 U528 ( .A1(n746), .A2(n399), .ZN(n396) );
  XNOR2_X1 U529 ( .A(n467), .B(n538), .ZN(n412) );
  XNOR2_X1 U530 ( .A(n628), .B(KEYINPUT22), .ZN(n631) );
  XNOR2_X1 U531 ( .A(n632), .B(n461), .ZN(n460) );
  NOR2_X2 U532 ( .A1(n783), .A2(n675), .ZN(n632) );
  NOR2_X1 U533 ( .A1(n775), .A2(n761), .ZN(n724) );
  INV_X1 U534 ( .A(n368), .ZN(n524) );
  NOR2_X1 U535 ( .A1(n662), .A2(G902), .ZN(n534) );
  NAND2_X1 U536 ( .A1(n369), .A2(n402), .ZN(n400) );
  XNOR2_X2 U537 ( .A(n386), .B(n507), .ZN(n746) );
  XNOR2_X1 U538 ( .A(n543), .B(n539), .ZN(n468) );
  NOR2_X1 U539 ( .A1(n707), .A2(n572), .ZN(n573) );
  NAND2_X1 U540 ( .A1(n391), .A2(n388), .ZN(n594) );
  NOR2_X1 U541 ( .A1(n510), .A2(n377), .ZN(n376) );
  INV_X1 U542 ( .A(n511), .ZN(n381) );
  NAND2_X1 U543 ( .A1(n607), .A2(n362), .ZN(n385) );
  XNOR2_X2 U544 ( .A(n771), .B(n496), .ZN(n386) );
  NAND2_X1 U545 ( .A1(n387), .A2(n478), .ZN(n477) );
  OR2_X2 U546 ( .A1(n387), .A2(KEYINPUT79), .ZN(n471) );
  INV_X1 U547 ( .A(n689), .ZN(n633) );
  INV_X1 U548 ( .A(n575), .ZN(n392) );
  OR2_X2 U549 ( .A1(n650), .A2(n627), .ZN(n689) );
  XNOR2_X2 U550 ( .A(n495), .B(n393), .ZN(n771) );
  XNOR2_X1 U551 ( .A(n468), .B(n393), .ZN(n467) );
  XNOR2_X2 U552 ( .A(n440), .B(n494), .ZN(n393) );
  NOR2_X1 U553 ( .A1(n746), .A2(n397), .ZN(n394) );
  NAND2_X1 U554 ( .A1(n640), .A2(KEYINPUT81), .ZN(n401) );
  INV_X1 U555 ( .A(n407), .ZN(n402) );
  NAND2_X1 U556 ( .A1(n640), .A2(n405), .ZN(n404) );
  AND2_X1 U557 ( .A1(n655), .A2(KEYINPUT81), .ZN(n405) );
  NAND2_X1 U558 ( .A1(n407), .A2(n655), .ZN(n406) );
  NAND2_X1 U559 ( .A1(n782), .A2(n642), .ZN(n408) );
  XNOR2_X2 U560 ( .A(n409), .B(n364), .ZN(n734) );
  NAND2_X1 U561 ( .A1(n410), .A2(n636), .ZN(n409) );
  XNOR2_X1 U562 ( .A(n646), .B(KEYINPUT104), .ZN(n410) );
  XNOR2_X2 U563 ( .A(n635), .B(n634), .ZN(n646) );
  XNOR2_X1 U564 ( .A(n574), .B(KEYINPUT42), .ZN(n788) );
  NOR2_X1 U565 ( .A1(n761), .A2(n723), .ZN(n726) );
  XNOR2_X2 U566 ( .A(n458), .B(n656), .ZN(n761) );
  XNOR2_X1 U567 ( .A(n535), .B(KEYINPUT28), .ZN(n437) );
  BUF_X1 U568 ( .A(n679), .Z(n414) );
  NOR2_X1 U569 ( .A1(n709), .A2(n627), .ZN(n417) );
  NOR2_X2 U570 ( .A1(n589), .A2(n624), .ZN(n590) );
  XNOR2_X1 U571 ( .A(n422), .B(n525), .ZN(n528) );
  XNOR2_X1 U572 ( .A(n524), .B(n423), .ZN(n422) );
  INV_X1 U573 ( .A(n523), .ZN(n423) );
  BUF_X1 U574 ( .A(n734), .Z(n425) );
  XNOR2_X1 U575 ( .A(n663), .B(n433), .ZN(n432) );
  NOR2_X1 U576 ( .A1(n426), .A2(G900), .ZN(n516) );
  INV_X1 U577 ( .A(n549), .ZN(n520) );
  NAND2_X1 U578 ( .A1(n679), .A2(n643), .ZN(n601) );
  XNOR2_X2 U579 ( .A(n590), .B(KEYINPUT74), .ZN(n679) );
  XNOR2_X1 U580 ( .A(n429), .B(n428), .ZN(G51) );
  NAND2_X1 U581 ( .A1(n485), .A2(n484), .ZN(n429) );
  NOR2_X1 U582 ( .A1(n575), .A2(n439), .ZN(n438) );
  INV_X1 U583 ( .A(n542), .ZN(n503) );
  NAND2_X1 U584 ( .A1(n432), .A2(n484), .ZN(n665) );
  XNOR2_X1 U585 ( .A(n744), .B(n430), .ZN(n747) );
  XNOR2_X1 U586 ( .A(n746), .B(n745), .ZN(n430) );
  XNOR2_X1 U587 ( .A(n431), .B(n367), .ZN(n489) );
  NAND2_X1 U588 ( .A1(n752), .A2(G472), .ZN(n431) );
  XNOR2_X2 U589 ( .A(n552), .B(G134), .ZN(n495) );
  XNOR2_X2 U590 ( .A(n470), .B(G131), .ZN(n552) );
  NAND2_X1 U591 ( .A1(n434), .A2(n657), .ZN(n660) );
  NAND2_X1 U592 ( .A1(n726), .A2(KEYINPUT2), .ZN(n434) );
  INV_X1 U593 ( .A(n687), .ZN(n476) );
  NAND2_X1 U594 ( .A1(n607), .A2(n710), .ZN(n613) );
  NOR2_X1 U595 ( .A1(n437), .A2(n355), .ZN(n536) );
  NOR2_X2 U596 ( .A1(n659), .A2(n660), .ZN(n752) );
  XNOR2_X1 U597 ( .A(n562), .B(n440), .ZN(n563) );
  NAND2_X2 U598 ( .A1(n492), .A2(n493), .ZN(n440) );
  NAND2_X1 U599 ( .A1(n752), .A2(G210), .ZN(n487) );
  INV_X1 U600 ( .A(n734), .ZN(n444) );
  NAND2_X1 U601 ( .A1(n734), .A2(KEYINPUT34), .ZN(n446) );
  INV_X1 U602 ( .A(n457), .ZN(n652) );
  INV_X1 U603 ( .A(n694), .ZN(n456) );
  OR2_X2 U604 ( .A1(n631), .A2(n636), .ZN(n457) );
  NAND2_X1 U605 ( .A1(n460), .A2(n639), .ZN(n459) );
  INV_X1 U606 ( .A(KEYINPUT44), .ZN(n461) );
  XNOR2_X1 U607 ( .A(n464), .B(n463), .ZN(G60) );
  NAND2_X1 U608 ( .A1(n465), .A2(n484), .ZN(n464) );
  XNOR2_X1 U609 ( .A(n466), .B(n366), .ZN(n465) );
  NAND2_X1 U610 ( .A1(n752), .A2(G475), .ZN(n466) );
  NAND2_X2 U611 ( .A1(n472), .A2(n471), .ZN(n658) );
  INV_X1 U612 ( .A(n607), .ZN(n480) );
  XNOR2_X1 U613 ( .A(n487), .B(n486), .ZN(n485) );
  NOR2_X1 U614 ( .A1(G952), .A2(n778), .ZN(n756) );
  INV_X1 U615 ( .A(KEYINPUT46), .ZN(n581) );
  XNOR2_X1 U616 ( .A(n582), .B(n581), .ZN(n600) );
  INV_X1 U617 ( .A(n667), .ZN(n653) );
  INV_X1 U618 ( .A(KEYINPUT80), .ZN(n655) );
  XNOR2_X1 U619 ( .A(n555), .B(n359), .ZN(n556) );
  XNOR2_X1 U620 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(n748) );
  XNOR2_X1 U622 ( .A(n658), .B(KEYINPUT78), .ZN(n775) );
  INV_X1 U623 ( .A(n740), .ZN(n741) );
  XOR2_X1 U624 ( .A(KEYINPUT38), .B(n593), .Z(n707) );
  BUF_X1 U625 ( .A(n593), .Z(n616) );
  NAND2_X1 U626 ( .A1(n489), .A2(n484), .ZN(n661) );
  INV_X1 U627 ( .A(G128), .ZN(n490) );
  NAND2_X1 U628 ( .A1(n490), .A2(G143), .ZN(n493) );
  INV_X1 U629 ( .A(G143), .ZN(n491) );
  NAND2_X1 U630 ( .A1(n491), .A2(G128), .ZN(n492) );
  XNOR2_X1 U631 ( .A(G146), .B(n539), .ZN(n496) );
  XNOR2_X1 U632 ( .A(n498), .B(n497), .ZN(n499) );
  NAND2_X1 U633 ( .A1(n551), .A2(G210), .ZN(n500) );
  XNOR2_X1 U634 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X2 U635 ( .A(KEYINPUT85), .B(G110), .Z(n540) );
  XOR2_X1 U636 ( .A(G137), .B(G140), .Z(n521) );
  XNOR2_X1 U637 ( .A(n506), .B(n505), .ZN(n507) );
  INV_X1 U638 ( .A(KEYINPUT67), .ZN(n508) );
  XNOR2_X1 U639 ( .A(G472), .B(KEYINPUT69), .ZN(n511) );
  NAND2_X1 U640 ( .A1(G952), .A2(n514), .ZN(n722) );
  NOR2_X1 U641 ( .A1(G953), .A2(n722), .ZN(n622) );
  NAND2_X1 U642 ( .A1(G902), .A2(n514), .ZN(n620) );
  OR2_X1 U643 ( .A1(n778), .A2(n620), .ZN(n515) );
  NOR2_X1 U644 ( .A1(n622), .A2(n516), .ZN(n575) );
  XOR2_X1 U645 ( .A(KEYINPUT90), .B(KEYINPUT21), .Z(n519) );
  INV_X1 U646 ( .A(n657), .ZN(n517) );
  NAND2_X1 U647 ( .A1(n530), .A2(G221), .ZN(n518) );
  XNOR2_X1 U648 ( .A(n522), .B(KEYINPUT89), .ZN(n525) );
  NAND2_X1 U649 ( .A1(G234), .A2(n778), .ZN(n526) );
  XOR2_X1 U650 ( .A(KEYINPUT8), .B(n526), .Z(n566) );
  NAND2_X1 U651 ( .A1(G221), .A2(n566), .ZN(n527) );
  XOR2_X1 U652 ( .A(KEYINPUT25), .B(KEYINPUT72), .Z(n532) );
  NAND2_X1 U653 ( .A1(n530), .A2(G217), .ZN(n531) );
  XNOR2_X1 U654 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U655 ( .A1(n697), .A2(n603), .ZN(n535) );
  XNOR2_X1 U656 ( .A(n536), .B(KEYINPUT109), .ZN(n589) );
  XOR2_X1 U657 ( .A(n537), .B(KEYINPUT73), .Z(n538) );
  XNOR2_X1 U658 ( .A(n550), .B(n540), .ZN(n541) );
  NOR2_X1 U659 ( .A1(n740), .A2(n657), .ZN(n548) );
  XNOR2_X1 U660 ( .A(n544), .B(KEYINPUT71), .ZN(n570) );
  NAND2_X1 U661 ( .A1(G210), .A2(n570), .ZN(n546) );
  INV_X1 U662 ( .A(KEYINPUT86), .ZN(n545) );
  XNOR2_X2 U663 ( .A(n548), .B(n547), .ZN(n593) );
  XNOR2_X1 U664 ( .A(n552), .B(KEYINPUT12), .ZN(n555) );
  NOR2_X1 U665 ( .A1(G902), .A2(n748), .ZN(n559) );
  XNOR2_X1 U666 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n558) );
  XNOR2_X1 U667 ( .A(KEYINPUT99), .B(G478), .ZN(n569) );
  XNOR2_X1 U668 ( .A(n564), .B(n563), .ZN(n565) );
  NAND2_X1 U669 ( .A1(G217), .A2(n566), .ZN(n567) );
  NOR2_X1 U670 ( .A1(G902), .A2(n751), .ZN(n568) );
  XNOR2_X1 U671 ( .A(n569), .B(n568), .ZN(n583) );
  INV_X1 U672 ( .A(n583), .ZN(n591) );
  NAND2_X1 U673 ( .A1(n592), .A2(n591), .ZN(n709) );
  NAND2_X1 U674 ( .A1(G214), .A2(n570), .ZN(n710) );
  INV_X1 U675 ( .A(n710), .ZN(n571) );
  OR2_X1 U676 ( .A1(n709), .A2(n571), .ZN(n572) );
  XNOR2_X1 U677 ( .A(n573), .B(KEYINPUT41), .ZN(n688) );
  NOR2_X1 U678 ( .A1(n589), .A2(n688), .ZN(n574) );
  XNOR2_X1 U679 ( .A(n693), .B(KEYINPUT91), .ZN(n627) );
  INV_X1 U680 ( .A(KEYINPUT39), .ZN(n576) );
  XNOR2_X1 U681 ( .A(n577), .B(n576), .ZN(n618) );
  INV_X1 U682 ( .A(n605), .ZN(n681) );
  AND2_X2 U683 ( .A1(n618), .A2(n681), .ZN(n580) );
  NOR2_X1 U684 ( .A1(n788), .A2(n787), .ZN(n582) );
  NAND2_X1 U685 ( .A1(n583), .A2(n592), .ZN(n584) );
  XNOR2_X1 U686 ( .A(KEYINPUT102), .B(n585), .ZN(n643) );
  INV_X1 U687 ( .A(n593), .ZN(n586) );
  NAND2_X1 U688 ( .A1(n586), .A2(n710), .ZN(n588) );
  INV_X1 U689 ( .A(KEYINPUT19), .ZN(n587) );
  NAND2_X1 U690 ( .A1(n601), .A2(KEYINPUT47), .ZN(n597) );
  NOR2_X1 U691 ( .A1(n592), .A2(n591), .ZN(n637) );
  NOR2_X1 U692 ( .A1(n594), .A2(n616), .ZN(n595) );
  NAND2_X1 U693 ( .A1(n637), .A2(n595), .ZN(n596) );
  XNOR2_X1 U694 ( .A(KEYINPUT108), .B(n596), .ZN(n786) );
  NAND2_X1 U695 ( .A1(n597), .A2(n786), .ZN(n598) );
  XNOR2_X1 U696 ( .A(n598), .B(KEYINPUT76), .ZN(n599) );
  OR2_X1 U697 ( .A1(KEYINPUT47), .A2(n601), .ZN(n609) );
  XNOR2_X1 U698 ( .A(KEYINPUT6), .B(KEYINPUT103), .ZN(n602) );
  NAND2_X1 U699 ( .A1(n636), .A2(n603), .ZN(n604) );
  NOR2_X1 U700 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U701 ( .A(KEYINPUT106), .B(n606), .ZN(n607) );
  XNOR2_X1 U702 ( .A(KEYINPUT107), .B(n613), .ZN(n614) );
  NAND2_X1 U703 ( .A1(n614), .A2(n690), .ZN(n615) );
  XNOR2_X1 U704 ( .A(KEYINPUT43), .B(n615), .ZN(n617) );
  NAND2_X1 U705 ( .A1(n617), .A2(n616), .ZN(n687) );
  NAND2_X1 U706 ( .A1(n618), .A2(n683), .ZN(n686) );
  INV_X1 U707 ( .A(n650), .ZN(n694) );
  NOR2_X1 U708 ( .A1(G898), .A2(n778), .ZN(n619) );
  XOR2_X1 U709 ( .A(KEYINPUT88), .B(n619), .Z(n765) );
  NOR2_X1 U710 ( .A1(n765), .A2(n620), .ZN(n621) );
  NOR2_X1 U711 ( .A1(n622), .A2(n621), .ZN(n623) );
  INV_X1 U712 ( .A(KEYINPUT0), .ZN(n625) );
  NOR2_X1 U713 ( .A1(n424), .A2(n631), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n690), .A2(n629), .ZN(n630) );
  NOR2_X1 U715 ( .A1(n694), .A2(n630), .ZN(n675) );
  INV_X1 U716 ( .A(KEYINPUT70), .ZN(n634) );
  XNOR2_X2 U717 ( .A(n638), .B(KEYINPUT35), .ZN(n782) );
  NAND2_X1 U718 ( .A1(n632), .A2(n782), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n782), .A2(KEYINPUT44), .ZN(n640) );
  INV_X1 U720 ( .A(KEYINPUT81), .ZN(n641) );
  AND2_X1 U721 ( .A1(KEYINPUT44), .A2(n641), .ZN(n642) );
  INV_X1 U722 ( .A(n643), .ZN(n712) );
  NAND2_X1 U723 ( .A1(n644), .A2(n418), .ZN(n645) );
  NOR2_X1 U724 ( .A1(n424), .A2(n645), .ZN(n672) );
  NAND2_X1 U725 ( .A1(n424), .A2(n356), .ZN(n702) );
  NOR2_X1 U726 ( .A1(n647), .A2(n702), .ZN(n648) );
  NOR2_X1 U727 ( .A1(n672), .A2(n684), .ZN(n649) );
  NOR2_X1 U728 ( .A1(n456), .A2(n435), .ZN(n651) );
  INV_X1 U729 ( .A(KEYINPUT45), .ZN(n656) );
  NOR2_X1 U730 ( .A1(KEYINPUT2), .A2(n724), .ZN(n659) );
  XNOR2_X1 U731 ( .A(n661), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U732 ( .A(n662), .B(KEYINPUT122), .ZN(n664) );
  NAND2_X1 U733 ( .A1(G217), .A2(n752), .ZN(n663) );
  XNOR2_X1 U734 ( .A(n665), .B(KEYINPUT123), .ZN(G66) );
  XOR2_X1 U735 ( .A(G101), .B(KEYINPUT111), .Z(n666) );
  XNOR2_X1 U736 ( .A(n667), .B(n666), .ZN(G3) );
  NAND2_X1 U737 ( .A1(n681), .A2(n672), .ZN(n668) );
  XNOR2_X1 U738 ( .A(n668), .B(G104), .ZN(G6) );
  XOR2_X1 U739 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n670) );
  XNOR2_X1 U740 ( .A(G107), .B(KEYINPUT26), .ZN(n669) );
  XNOR2_X1 U741 ( .A(n670), .B(n669), .ZN(n671) );
  XOR2_X1 U742 ( .A(KEYINPUT27), .B(n671), .Z(n674) );
  NAND2_X1 U743 ( .A1(n672), .A2(n683), .ZN(n673) );
  XNOR2_X1 U744 ( .A(n674), .B(n673), .ZN(G9) );
  XOR2_X1 U745 ( .A(G110), .B(n675), .Z(G12) );
  XOR2_X1 U746 ( .A(KEYINPUT29), .B(KEYINPUT114), .Z(n677) );
  NAND2_X1 U747 ( .A1(n683), .A2(n414), .ZN(n676) );
  XNOR2_X1 U748 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U749 ( .A(G128), .B(n678), .ZN(G30) );
  NAND2_X1 U750 ( .A1(n681), .A2(n414), .ZN(n680) );
  XNOR2_X1 U751 ( .A(G146), .B(n680), .ZN(G48) );
  NAND2_X1 U752 ( .A1(n684), .A2(n681), .ZN(n682) );
  XNOR2_X1 U753 ( .A(n682), .B(G113), .ZN(G15) );
  NAND2_X1 U754 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U755 ( .A(n685), .B(G116), .ZN(G18) );
  XNOR2_X1 U756 ( .A(G134), .B(n686), .ZN(G36) );
  XNOR2_X1 U757 ( .A(G140), .B(n687), .ZN(G42) );
  XOR2_X1 U758 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n692) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U760 ( .A(n692), .B(n691), .ZN(n700) );
  NOR2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U762 ( .A(KEYINPUT49), .B(n695), .Z(n696) );
  NOR2_X1 U763 ( .A1(n424), .A2(n696), .ZN(n698) );
  XNOR2_X1 U764 ( .A(n698), .B(KEYINPUT115), .ZN(n699) );
  NOR2_X1 U765 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U766 ( .A(KEYINPUT117), .B(n701), .ZN(n703) );
  NAND2_X1 U767 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U768 ( .A(n704), .B(KEYINPUT118), .ZN(n705) );
  XNOR2_X1 U769 ( .A(n705), .B(KEYINPUT51), .ZN(n706) );
  NOR2_X1 U770 ( .A1(n688), .A2(n706), .ZN(n718) );
  INV_X1 U771 ( .A(n707), .ZN(n711) );
  NOR2_X1 U772 ( .A1(n711), .A2(n710), .ZN(n708) );
  NOR2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n715) );
  NAND2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n713) );
  NOR2_X1 U775 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U776 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U777 ( .A1(n425), .A2(n716), .ZN(n717) );
  NOR2_X1 U778 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U779 ( .A(n719), .B(KEYINPUT52), .Z(n720) );
  XNOR2_X1 U780 ( .A(KEYINPUT119), .B(n720), .ZN(n721) );
  NOR2_X1 U781 ( .A1(n722), .A2(n721), .ZN(n731) );
  INV_X1 U782 ( .A(KEYINPUT2), .ZN(n732) );
  OR2_X1 U783 ( .A1(n723), .A2(n732), .ZN(n725) );
  NAND2_X1 U784 ( .A1(n725), .A2(n724), .ZN(n729) );
  NOR2_X1 U785 ( .A1(n726), .A2(KEYINPUT75), .ZN(n727) );
  NAND2_X1 U786 ( .A1(n727), .A2(KEYINPUT2), .ZN(n728) );
  NAND2_X1 U787 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U788 ( .A1(n731), .A2(n730), .ZN(n738) );
  NAND2_X1 U789 ( .A1(KEYINPUT75), .A2(n732), .ZN(n733) );
  NAND2_X1 U790 ( .A1(n778), .A2(n733), .ZN(n736) );
  NOR2_X1 U791 ( .A1(n425), .A2(n688), .ZN(n735) );
  NOR2_X1 U792 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U793 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U794 ( .A(KEYINPUT53), .B(n739), .Z(G75) );
  XOR2_X1 U795 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n743) );
  XNOR2_X1 U796 ( .A(KEYINPUT82), .B(KEYINPUT83), .ZN(n742) );
  XOR2_X1 U797 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n745) );
  NAND2_X1 U798 ( .A1(n752), .A2(G469), .ZN(n744) );
  NOR2_X1 U799 ( .A1(n756), .A2(n747), .ZN(G54) );
  XOR2_X1 U800 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n750) );
  XNOR2_X1 U801 ( .A(n748), .B(KEYINPUT64), .ZN(n749) );
  XOR2_X1 U802 ( .A(n751), .B(KEYINPUT121), .Z(n754) );
  NAND2_X1 U803 ( .A1(n752), .A2(G478), .ZN(n753) );
  XNOR2_X1 U804 ( .A(n754), .B(n753), .ZN(n755) );
  NOR2_X1 U805 ( .A1(n756), .A2(n755), .ZN(G63) );
  XOR2_X1 U806 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n758) );
  NAND2_X1 U807 ( .A1(G224), .A2(G953), .ZN(n757) );
  XNOR2_X1 U808 ( .A(n758), .B(n757), .ZN(n759) );
  XNOR2_X1 U809 ( .A(KEYINPUT124), .B(n759), .ZN(n760) );
  NAND2_X1 U810 ( .A1(G898), .A2(n760), .ZN(n763) );
  OR2_X1 U811 ( .A1(n761), .A2(G953), .ZN(n762) );
  NAND2_X1 U812 ( .A1(n763), .A2(n762), .ZN(n769) );
  XNOR2_X1 U813 ( .A(n764), .B(G101), .ZN(n766) );
  NAND2_X1 U814 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U815 ( .A(n767), .B(KEYINPUT126), .ZN(n768) );
  XOR2_X1 U816 ( .A(n769), .B(n768), .Z(G69) );
  XOR2_X1 U817 ( .A(n771), .B(n770), .Z(n776) );
  INV_X1 U818 ( .A(n776), .ZN(n772) );
  XNOR2_X1 U819 ( .A(G227), .B(n772), .ZN(n773) );
  NAND2_X1 U820 ( .A1(n773), .A2(G900), .ZN(n774) );
  NAND2_X1 U821 ( .A1(n774), .A2(G953), .ZN(n781) );
  XNOR2_X1 U822 ( .A(n776), .B(n775), .ZN(n777) );
  XNOR2_X1 U823 ( .A(n777), .B(KEYINPUT127), .ZN(n779) );
  NAND2_X1 U824 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U825 ( .A1(n781), .A2(n780), .ZN(G72) );
  XOR2_X1 U826 ( .A(n782), .B(G122), .Z(G24) );
  XOR2_X1 U827 ( .A(n783), .B(G119), .Z(G21) );
  XOR2_X1 U828 ( .A(G125), .B(n784), .Z(n785) );
  XNOR2_X1 U829 ( .A(KEYINPUT37), .B(n785), .ZN(G27) );
  XNOR2_X1 U830 ( .A(n786), .B(G143), .ZN(G45) );
  XOR2_X1 U831 ( .A(n787), .B(G131), .Z(G33) );
  XOR2_X1 U832 ( .A(n788), .B(G137), .Z(G39) );
endmodule

