//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G469), .ZN(new_n192));
  XNOR2_X1  g006(.A(G110), .B(G140), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n194), .A2(G227), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n193), .B(new_n195), .Z(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT76), .B1(new_n197), .B2(G104), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n199));
  INV_X1    g013(.A(G104), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G107), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  OR3_X1    g017(.A1(new_n200), .A2(KEYINPUT3), .A3(G107), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n197), .A2(G104), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT3), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n202), .A2(new_n203), .A3(new_n204), .A4(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT78), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n208), .B1(new_n197), .B2(G104), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n200), .A2(KEYINPUT78), .A3(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n205), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G101), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n207), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G143), .ZN(new_n215));
  INV_X1    g029(.A(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n216), .C2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G128), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT67), .B1(new_n215), .B2(KEYINPUT1), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n218), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(new_n214), .B2(G143), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n215), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n223), .A2(new_n214), .A3(G143), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n225), .A2(new_n226), .A3(G128), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT81), .B1(new_n213), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(new_n227), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n216), .A2(G146), .ZN(new_n232));
  OAI21_X1  g046(.A(G128), .B1(new_n232), .B2(new_n226), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n228), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n213), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n207), .A2(new_n212), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT81), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n237), .A2(new_n238), .A3(new_n228), .A4(new_n222), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n230), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(KEYINPUT65), .A2(G134), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT65), .A2(G134), .ZN(new_n242));
  OAI21_X1  g056(.A(G137), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g059(.A(KEYINPUT66), .B(G137), .C1(new_n241), .C2(new_n242), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OR2_X1    g061(.A1(KEYINPUT65), .A2(G134), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT11), .ZN(new_n249));
  INV_X1    g063(.A(G137), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT65), .A2(G134), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n248), .A2(new_n249), .A3(new_n250), .A4(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G134), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT11), .B1(new_n253), .B2(G137), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n247), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G131), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n247), .A2(new_n258), .A3(new_n255), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n240), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT12), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n240), .A2(KEYINPUT12), .A3(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT80), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n257), .A2(new_n259), .A3(new_n266), .ZN(new_n267));
  AOI221_X4 g081(.A(G131), .B1(new_n252), .B2(new_n254), .C1(new_n245), .C2(new_n246), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n258), .B1(new_n247), .B2(new_n255), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT80), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT10), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n272), .B1(new_n222), .B2(new_n228), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n213), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT79), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n213), .A3(KEYINPUT79), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n207), .A2(KEYINPUT4), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n202), .A2(new_n206), .A3(new_n204), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n203), .A2(KEYINPUT77), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(KEYINPUT4), .A3(new_n281), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT64), .B1(new_n216), .B2(G146), .ZN(new_n286));
  OAI211_X1 g100(.A(G128), .B(new_n227), .C1(new_n286), .C2(new_n232), .ZN(new_n287));
  INV_X1    g101(.A(G128), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n218), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n289), .A3(KEYINPUT0), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n218), .A2(G128), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT0), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n285), .A2(new_n294), .B1(new_n236), .B2(new_n272), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n271), .A2(new_n278), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n196), .B1(new_n265), .B2(new_n296), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n271), .A2(new_n278), .A3(new_n295), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n278), .A2(new_n295), .B1(new_n259), .B2(new_n257), .ZN(new_n299));
  INV_X1    g113(.A(new_n196), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT82), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT82), .ZN(new_n303));
  INV_X1    g117(.A(new_n299), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n296), .A3(new_n196), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n298), .B1(new_n264), .B2(new_n263), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n303), .B(new_n305), .C1(new_n306), .C2(new_n196), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n192), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n300), .B1(new_n298), .B2(new_n299), .ZN(new_n309));
  INV_X1    g123(.A(new_n264), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT12), .B1(new_n240), .B2(new_n260), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n296), .B(new_n196), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n192), .A3(new_n189), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n192), .A2(new_n189), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n191), .B1(new_n308), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT83), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT83), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n320), .B(new_n191), .C1(new_n308), .C2(new_n317), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n248), .A2(new_n251), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(G137), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n250), .A2(G134), .ZN(new_n325));
  OAI21_X1  g139(.A(G131), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n259), .A2(new_n229), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT68), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n328), .B1(new_n260), .B2(new_n294), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n328), .B(new_n294), .C1(new_n268), .C2(new_n269), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n327), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  XOR2_X1   g146(.A(G116), .B(G119), .Z(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT2), .B(G113), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n327), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n294), .B1(new_n268), .B2(new_n269), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT68), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n337), .B1(new_n339), .B2(new_n330), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n333), .B(new_n334), .Z(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n336), .A2(KEYINPUT70), .A3(new_n342), .ZN(new_n343));
  OR3_X1    g157(.A1(new_n340), .A2(KEYINPUT70), .A3(new_n341), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(KEYINPUT28), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n338), .A2(new_n327), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT69), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT69), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n338), .A2(new_n348), .A3(new_n327), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n341), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(G237), .A2(G953), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G210), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(new_n203), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n356));
  XOR2_X1   g170(.A(new_n355), .B(new_n356), .Z(new_n357));
  AND4_X1   g171(.A1(KEYINPUT29), .A2(new_n345), .A3(new_n352), .A4(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n341), .B1(new_n338), .B2(new_n327), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(new_n340), .B2(new_n341), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n352), .B(new_n357), .C1(new_n360), .C2(new_n351), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT29), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI211_X1 g177(.A(new_n335), .B(new_n337), .C1(new_n339), .C2(new_n330), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT30), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n338), .A2(new_n365), .A3(new_n327), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(new_n340), .B2(new_n365), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n364), .B1(new_n367), .B2(new_n335), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(new_n357), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n189), .B1(new_n363), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G472), .B1(new_n358), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n366), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(new_n332), .B2(KEYINPUT30), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n342), .B(new_n357), .C1(new_n373), .C2(new_n341), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT31), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n352), .B1(new_n360), .B2(new_n351), .ZN(new_n376));
  INV_X1    g190(.A(new_n357), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT31), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n368), .A2(new_n379), .A3(new_n357), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n375), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT32), .ZN(new_n382));
  NOR2_X1   g196(.A1(G472), .A2(G902), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n382), .B1(new_n381), .B2(new_n383), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n371), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G110), .B(G122), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n341), .B1(new_n283), .B2(new_n284), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n333), .A2(new_n334), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT5), .ZN(new_n391));
  INV_X1    g205(.A(G119), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G116), .ZN(new_n393));
  OAI211_X1 g207(.A(G113), .B(new_n393), .C1(new_n333), .C2(new_n391), .ZN(new_n394));
  AND4_X1   g208(.A1(new_n390), .A2(new_n394), .A3(new_n207), .A4(new_n212), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n388), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  AOI22_X1  g210(.A1(KEYINPUT4), .A2(new_n207), .B1(new_n280), .B2(new_n281), .ZN(new_n397));
  INV_X1    g211(.A(new_n284), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n335), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n395), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(new_n387), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n396), .A2(new_n401), .A3(KEYINPUT6), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n290), .A2(G125), .A3(new_n293), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n404));
  INV_X1    g218(.A(G125), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n222), .A2(new_n405), .A3(new_n228), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G224), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(G953), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n290), .A2(KEYINPUT84), .A3(G125), .A4(new_n293), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n407), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n410), .B1(new_n407), .B2(new_n411), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n415), .B(new_n388), .C1(new_n389), .C2(new_n395), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n402), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n407), .A2(new_n411), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n409), .B(KEYINPUT86), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(KEYINPUT7), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n410), .A2(KEYINPUT7), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n407), .A2(new_n421), .A3(new_n411), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n387), .B(KEYINPUT85), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(KEYINPUT8), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n213), .B1(new_n390), .B2(new_n394), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n424), .B1(new_n425), .B2(new_n395), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n420), .A2(new_n422), .A3(new_n426), .A4(new_n401), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n417), .A2(new_n189), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G210), .B1(G237), .B2(G902), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n417), .A2(new_n189), .A3(new_n429), .A4(new_n427), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G214), .B1(G237), .B2(G902), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G237), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n194), .A3(G214), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT87), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n216), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n353), .B(G214), .C1(KEYINPUT87), .C2(G143), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G131), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT17), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(new_n258), .A3(new_n440), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n405), .A2(KEYINPUT16), .A3(G140), .ZN(new_n446));
  XNOR2_X1  g260(.A(G125), .B(G140), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n446), .B1(new_n447), .B2(KEYINPUT16), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(G146), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(G146), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n441), .A2(KEYINPUT17), .A3(G131), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n445), .A2(new_n450), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n441), .A2(KEYINPUT18), .A3(G131), .ZN(new_n454));
  AND2_X1   g268(.A1(KEYINPUT18), .A2(G131), .ZN(new_n455));
  XOR2_X1   g269(.A(G125), .B(G140), .Z(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT88), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT88), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n447), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n214), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n456), .A2(G146), .ZN(new_n461));
  OAI221_X1 g275(.A(new_n454), .B1(new_n441), .B2(new_n455), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n453), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G113), .B(G122), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(new_n200), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n465), .A2(KEYINPUT90), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n189), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n463), .A2(new_n466), .ZN(new_n469));
  OAI21_X1  g283(.A(G475), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT20), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n463), .A2(new_n465), .ZN(new_n472));
  INV_X1    g286(.A(new_n451), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n473), .B1(new_n442), .B2(new_n444), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n457), .A2(new_n459), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT19), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n456), .A2(KEYINPUT19), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n214), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n465), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n480), .A3(new_n462), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n472), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(G475), .A2(G902), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(KEYINPUT89), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n471), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n465), .B1(new_n474), .B2(new_n478), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n462), .A2(new_n486), .B1(new_n463), .B2(new_n465), .ZN(new_n487));
  INV_X1    g301(.A(new_n484), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(KEYINPUT20), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n470), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT91), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT91), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n470), .A2(new_n485), .A3(new_n492), .A4(new_n489), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G116), .B(G122), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(G107), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT92), .B1(new_n288), .B2(G143), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT92), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n216), .A3(G128), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT13), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT93), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT13), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n288), .A2(G143), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n500), .A2(new_n506), .A3(new_n501), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n503), .A2(new_n504), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n496), .B1(new_n508), .B2(G134), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n500), .A2(new_n323), .A3(new_n505), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G116), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(KEYINPUT14), .A3(G122), .ZN(new_n514));
  INV_X1    g328(.A(new_n495), .ZN(new_n515));
  OAI211_X1 g329(.A(G107), .B(new_n514), .C1(new_n515), .C2(KEYINPUT14), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n495), .A2(new_n197), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n323), .B1(new_n500), .B2(new_n505), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n516), .B(new_n517), .C1(new_n510), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n188), .A2(G217), .A3(new_n194), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n521), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n512), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n189), .ZN(new_n526));
  INV_X1    g340(.A(G478), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n526), .A2(new_n528), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(G234), .A2(G237), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(G952), .A3(new_n194), .ZN(new_n533));
  XOR2_X1   g347(.A(new_n533), .B(KEYINPUT94), .Z(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  XOR2_X1   g349(.A(KEYINPUT21), .B(G898), .Z(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n532), .A2(G902), .A3(G953), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n535), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n494), .A2(new_n531), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT95), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n494), .A2(new_n531), .A3(KEYINPUT95), .A4(new_n541), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n435), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n392), .A2(G128), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT23), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT72), .B1(new_n288), .B2(G119), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G110), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n288), .A2(G119), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT24), .B(G110), .Z(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n551), .B(new_n555), .C1(new_n473), .C2(new_n449), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT73), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  OAI22_X1  g372(.A1(new_n550), .A2(G110), .B1(new_n553), .B2(new_n554), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n559), .B(new_n451), .C1(G146), .C2(new_n456), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT22), .B(G137), .ZN(new_n561));
  INV_X1    g375(.A(G234), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n187), .A2(new_n562), .A3(G953), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n561), .B(new_n563), .Z(new_n564));
  AND3_X1   g378(.A1(new_n558), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n564), .B1(new_n558), .B2(new_n560), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(KEYINPUT25), .A3(new_n189), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n558), .A2(new_n560), .ZN(new_n569));
  INV_X1    g383(.A(new_n564), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n558), .A2(new_n560), .A3(new_n564), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n189), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT25), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n568), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G217), .B1(new_n562), .B2(G902), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n577), .B(KEYINPUT71), .Z(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(G902), .B1(new_n562), .B2(G217), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n581), .B(KEYINPUT74), .Z(new_n582));
  NAND2_X1  g396(.A1(new_n567), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(KEYINPUT75), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT75), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n578), .B1(new_n568), .B2(new_n575), .ZN(new_n586));
  INV_X1    g400(.A(new_n583), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n322), .A2(new_n386), .A3(new_n546), .A4(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  NAND2_X1  g405(.A1(new_n381), .A2(new_n383), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(G472), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n381), .B2(new_n189), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n322), .A2(new_n589), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT96), .ZN(new_n598));
  INV_X1    g412(.A(new_n434), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n431), .B2(new_n432), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(KEYINPUT97), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n602));
  AOI211_X1 g416(.A(new_n602), .B(new_n599), .C1(new_n431), .C2(new_n432), .ZN(new_n603));
  AOI211_X1 g417(.A(G478), .B(G902), .C1(new_n522), .C2(new_n524), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT33), .B1(new_n523), .B2(KEYINPUT98), .ZN(new_n605));
  INV_X1    g419(.A(new_n524), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n523), .B1(new_n512), .B2(new_n519), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n605), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n522), .A2(new_n524), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n604), .B1(new_n611), .B2(G478), .ZN(new_n612));
  NAND2_X1  g426(.A1(G478), .A2(G902), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n612), .A2(new_n491), .A3(new_n493), .A4(new_n613), .ZN(new_n614));
  NOR4_X1   g428(.A1(new_n601), .A2(new_n603), .A3(new_n614), .A4(new_n540), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n598), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G104), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT99), .B(KEYINPUT34), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  NAND2_X1  g434(.A1(new_n435), .A2(new_n602), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n529), .A2(new_n530), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n600), .A2(KEYINPUT97), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n621), .A2(new_n622), .A3(new_n541), .A4(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n598), .A2(new_n490), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT35), .B(G107), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  INV_X1    g441(.A(new_n582), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n570), .A2(KEYINPUT36), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n569), .B(new_n629), .Z(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n580), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n322), .A2(new_n546), .A3(new_n596), .A4(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT37), .B(G110), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G12));
  INV_X1    g449(.A(G900), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n535), .B1(new_n636), .B2(new_n539), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n531), .A2(new_n490), .A3(new_n637), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n638), .A2(new_n621), .A3(new_n623), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n322), .A2(new_n386), .A3(new_n639), .A4(new_n632), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G128), .ZN(G30));
  NAND2_X1  g455(.A1(new_n592), .A2(KEYINPUT32), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n368), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n357), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n189), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n357), .B1(new_n343), .B2(new_n344), .ZN(new_n648));
  OAI21_X1  g462(.A(G472), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT100), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n644), .A2(new_n652), .A3(new_n649), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NOR4_X1   g468(.A1(new_n632), .A2(new_n531), .A3(new_n494), .A4(new_n599), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n433), .B(KEYINPUT38), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n654), .A2(KEYINPUT101), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n651), .A2(new_n655), .A3(new_n653), .A4(new_n656), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n637), .B(KEYINPUT39), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n322), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT40), .Z(new_n664));
  NAND3_X1  g478(.A1(new_n657), .A2(new_n660), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G143), .ZN(G45));
  AND2_X1   g480(.A1(new_n386), .A2(new_n632), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n601), .A2(new_n603), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n614), .A2(new_n637), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n667), .A2(new_n322), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G146), .ZN(G48));
  AOI21_X1  g485(.A(G902), .B1(new_n309), .B2(new_n312), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n672), .A2(new_n192), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n191), .A3(new_n314), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n386), .A2(new_n615), .A3(new_n589), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT41), .B(G113), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G15));
  NOR2_X1   g492(.A1(new_n624), .A2(new_n490), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n679), .A2(new_n386), .A3(new_n589), .A4(new_n675), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G116), .ZN(G18));
  NAND2_X1  g495(.A1(new_n544), .A2(new_n545), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n674), .A2(new_n601), .A3(new_n603), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n386), .A2(new_n682), .A3(new_n632), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  INV_X1    g499(.A(new_n383), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n375), .A2(new_n380), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n345), .A2(new_n352), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n377), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n686), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n580), .A2(new_n583), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n690), .A2(new_n595), .A3(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n601), .A2(new_n603), .A3(new_n540), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n494), .A2(new_n531), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n692), .A2(new_n693), .A3(new_n694), .A4(new_n675), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G122), .ZN(G24));
  NOR2_X1   g510(.A1(new_n690), .A2(new_n595), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n697), .A2(new_n632), .A3(new_n669), .A4(new_n683), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G125), .ZN(G27));
  NOR2_X1   g513(.A1(new_n433), .A2(new_n599), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n265), .A2(new_n296), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n300), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(G469), .A3(new_n305), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n314), .A3(new_n316), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n700), .A2(new_n704), .A3(new_n191), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n386), .A2(new_n589), .A3(new_n669), .A4(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT42), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n691), .B1(new_n644), .B2(new_n371), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n705), .A2(new_n669), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n707), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n706), .A2(new_n707), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n258), .ZN(G33));
  NAND4_X1  g526(.A1(new_n386), .A2(new_n589), .A3(new_n638), .A4(new_n705), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n713), .A2(KEYINPUT102), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(KEYINPUT102), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G134), .ZN(G36));
  NAND3_X1  g531(.A1(new_n702), .A2(KEYINPUT45), .A3(new_n305), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n719));
  OR2_X1    g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n192), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n302), .A2(new_n307), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n315), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT46), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n314), .B1(new_n725), .B2(KEYINPUT46), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n191), .B(new_n662), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n494), .A2(new_n613), .A3(new_n612), .ZN(new_n730));
  XOR2_X1   g544(.A(new_n730), .B(KEYINPUT43), .Z(new_n731));
  INV_X1    g545(.A(new_n596), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n732), .A3(new_n632), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n700), .B1(new_n733), .B2(new_n734), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n729), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n250), .ZN(G39));
  INV_X1    g552(.A(KEYINPUT47), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(KEYINPUT104), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n720), .A2(new_n721), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(G469), .A3(new_n724), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n316), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n744), .A2(new_n745), .B1(new_n192), .B2(new_n672), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n190), .B1(new_n746), .B2(new_n726), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n739), .A2(KEYINPUT104), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n741), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n700), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n386), .A2(new_n589), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n191), .B1(new_n727), .B2(new_n728), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n740), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n750), .A2(new_n669), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G140), .ZN(G42));
  NAND2_X1  g570(.A1(new_n731), .A2(new_n535), .ZN(new_n757));
  INV_X1    g571(.A(new_n692), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n757), .A2(new_n758), .A3(new_n751), .ZN(new_n759));
  XOR2_X1   g573(.A(new_n759), .B(KEYINPUT111), .Z(new_n760));
  AND2_X1   g574(.A1(new_n750), .A2(new_n754), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n673), .A2(new_n314), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n191), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n760), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n675), .A2(new_n700), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT112), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n765), .A2(KEYINPUT112), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n757), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n632), .A3(new_n697), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n757), .A2(new_n674), .A3(new_n758), .ZN(new_n770));
  INV_X1    g584(.A(new_n656), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n599), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n770), .A2(KEYINPUT50), .A3(new_n599), .A4(new_n771), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n651), .A2(new_n653), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n767), .A2(new_n766), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n589), .A2(new_n776), .A3(new_n535), .A4(new_n777), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n613), .A2(new_n612), .B1(new_n491), .B2(new_n493), .ZN(new_n779));
  AOI22_X1  g593(.A1(new_n774), .A2(new_n775), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n764), .A2(new_n769), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n768), .A2(new_n708), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n784), .A2(KEYINPUT113), .ZN(new_n785));
  OR2_X1    g599(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(KEYINPUT113), .ZN(new_n787));
  NAND2_X1  g601(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n785), .A2(new_n786), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n614), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n778), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n789), .A2(G952), .A3(new_n194), .A4(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n786), .B1(new_n785), .B2(new_n787), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n764), .A2(KEYINPUT51), .A3(new_n769), .A4(new_n780), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n783), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n770), .A2(new_n668), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n680), .A2(new_n684), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n695), .A2(new_n676), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT107), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n680), .A2(new_n695), .A3(new_n676), .A4(new_n684), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT107), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n711), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n322), .A2(new_n386), .A3(new_n632), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n490), .A2(new_n637), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n751), .A2(new_n622), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n806), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n322), .A2(new_n386), .A3(new_n632), .A4(new_n808), .ZN(new_n811));
  INV_X1    g625(.A(new_n809), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT108), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n622), .A2(new_n494), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n540), .B(new_n435), .C1(new_n815), .C2(new_n614), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n322), .A2(new_n816), .A3(new_n589), .A4(new_n596), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n697), .A2(new_n632), .A3(new_n669), .A4(new_n705), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n590), .A2(new_n633), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n714), .B2(new_n715), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n804), .A2(new_n805), .A3(new_n814), .A4(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(KEYINPUT53), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT109), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n322), .A2(new_n386), .A3(new_n668), .A4(new_n632), .ZN(new_n825));
  INV_X1    g639(.A(new_n669), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n640), .B(new_n698), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n191), .A2(new_n668), .A3(new_n694), .A4(new_n704), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n632), .A2(new_n637), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n650), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n824), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n640), .A2(new_n698), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n670), .A3(KEYINPUT52), .A4(new_n830), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n823), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n832), .A2(new_n834), .A3(new_n823), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n822), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n819), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n814), .A2(new_n716), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n832), .A2(new_n834), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n841), .A2(new_n805), .A3(new_n842), .A4(new_n804), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT53), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n839), .A2(KEYINPUT54), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT110), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(new_n802), .B2(new_n711), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT53), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n814), .A2(new_n716), .A3(new_n840), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n802), .A2(new_n711), .A3(new_n846), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n838), .A2(new_n851), .B1(new_n843), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n796), .A2(new_n797), .A3(new_n845), .A4(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(G952), .A2(G953), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT115), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n691), .A2(new_n190), .A3(new_n599), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(KEYINPUT105), .Z(new_n861));
  INV_X1    g675(.A(new_n730), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n762), .A2(KEYINPUT49), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT106), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n771), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n865), .B2(new_n864), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n867), .B(new_n776), .C1(KEYINPUT49), .C2(new_n762), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n859), .A2(new_n868), .ZN(G75));
  NOR2_X1   g683(.A1(new_n848), .A2(new_n849), .ZN(new_n870));
  INV_X1    g684(.A(new_n850), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n832), .A2(new_n823), .A3(new_n834), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n870), .B(new_n871), .C1(new_n835), .C2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n842), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n852), .B1(new_n821), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(G210), .A3(G902), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT56), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n402), .A2(new_n416), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n414), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n194), .A2(G952), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n853), .A2(new_n189), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT56), .B1(new_n887), .B2(G210), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n882), .B1(new_n888), .B2(new_n878), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n878), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(G51));
  XNOR2_X1  g705(.A(new_n853), .B(KEYINPUT54), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n315), .B(KEYINPUT57), .Z(new_n893));
  OAI21_X1  g707(.A(new_n313), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n887), .A2(new_n724), .A3(new_n722), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n884), .B1(new_n894), .B2(new_n895), .ZN(G54));
  NAND3_X1  g710(.A1(new_n887), .A2(KEYINPUT58), .A3(G475), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n897), .A2(new_n482), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n482), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n898), .A2(new_n899), .A3(new_n884), .ZN(G60));
  XOR2_X1   g714(.A(new_n613), .B(KEYINPUT59), .Z(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n855), .B2(new_n845), .ZN(new_n902));
  INV_X1    g716(.A(new_n611), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n885), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n892), .A2(new_n901), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n904), .B1(new_n903), .B2(new_n905), .ZN(G63));
  NAND2_X1  g720(.A1(G217), .A2(G902), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT118), .ZN(new_n908));
  XNOR2_X1  g722(.A(KEYINPUT117), .B(KEYINPUT60), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n908), .B(new_n909), .Z(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n873), .B2(new_n875), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n630), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT61), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n567), .B(KEYINPUT120), .Z(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n885), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(KEYINPUT121), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n876), .A2(new_n910), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n884), .B1(new_n919), .B2(new_n915), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n920), .A2(new_n921), .A3(KEYINPUT61), .A4(new_n913), .ZN(new_n922));
  NOR4_X1   g736(.A1(new_n853), .A2(KEYINPUT119), .A3(new_n631), .A4(new_n911), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT119), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n912), .B2(new_n630), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n917), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n918), .B(new_n922), .C1(new_n926), .C2(KEYINPUT61), .ZN(G66));
  OAI21_X1  g741(.A(G953), .B1(new_n537), .B2(new_n408), .ZN(new_n928));
  INV_X1    g742(.A(new_n804), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n590), .A2(new_n633), .A3(new_n817), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n928), .B1(new_n931), .B2(G953), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n880), .B1(G898), .B2(new_n194), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(G69));
  NOR2_X1   g748(.A1(new_n737), .A2(new_n827), .ZN(new_n935));
  INV_X1    g749(.A(new_n729), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n936), .A2(new_n668), .A3(new_n694), .A4(new_n708), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n711), .B1(new_n714), .B2(new_n715), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n935), .A2(new_n755), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT124), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n476), .A2(new_n477), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n367), .B(new_n942), .ZN(new_n943));
  OR3_X1    g757(.A1(new_n941), .A2(G953), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n827), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n665), .A2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT122), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(KEYINPUT122), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n946), .B2(new_n948), .ZN(new_n951));
  INV_X1    g765(.A(new_n737), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n755), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n663), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n386), .A2(new_n589), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n815), .A2(new_n614), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n954), .A2(new_n955), .A3(new_n700), .A4(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n949), .A2(new_n951), .A3(new_n953), .A4(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n943), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(G953), .B1(new_n943), .B2(new_n636), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT123), .Z(new_n963));
  NAND4_X1  g777(.A1(new_n944), .A2(new_n960), .A3(new_n961), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n636), .A2(KEYINPUT125), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n636), .A2(KEYINPUT125), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n959), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n962), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT126), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n964), .A2(new_n969), .ZN(G72));
  AOI22_X1  g784(.A1(new_n822), .A2(new_n838), .B1(KEYINPUT53), .B2(new_n843), .ZN(new_n971));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT63), .Z(new_n973));
  NAND2_X1  g787(.A1(new_n368), .A2(new_n377), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n971), .A2(new_n646), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n973), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n941), .B2(new_n931), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n975), .B(new_n885), .C1(new_n977), .C2(new_n974), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n979));
  INV_X1    g793(.A(new_n931), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n973), .B1(new_n958), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n646), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n981), .A2(new_n979), .A3(new_n982), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n978), .A2(new_n983), .A3(new_n984), .ZN(G57));
endmodule


