

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U550 ( .A1(n518), .A2(G2105), .ZN(n975) );
  AND2_X2 U551 ( .A1(n518), .A2(G2105), .ZN(n982) );
  NOR2_X2 U552 ( .A1(n613), .A2(n612), .ZN(n1006) );
  NOR2_X2 U553 ( .A1(n667), .A2(n596), .ZN(n598) );
  XNOR2_X2 U554 ( .A(n676), .B(KEYINPUT32), .ZN(n693) );
  AND2_X2 U555 ( .A1(n675), .A2(n674), .ZN(n676) );
  AND2_X1 U556 ( .A1(n715), .A2(G40), .ZN(n587) );
  AND2_X1 U557 ( .A1(n702), .A2(n517), .ZN(n703) );
  NOR2_X1 U558 ( .A1(n734), .A2(n516), .ZN(n735) );
  NOR2_X1 U559 ( .A1(G543), .A2(G651), .ZN(n782) );
  AND2_X1 U560 ( .A1(n736), .A2(n735), .ZN(n515) );
  AND2_X1 U561 ( .A1(n748), .A2(n900), .ZN(n516) );
  OR2_X1 U562 ( .A1(n701), .A2(n700), .ZN(n517) );
  XNOR2_X1 U563 ( .A(n601), .B(KEYINPUT93), .ZN(n614) );
  INV_X1 U564 ( .A(KEYINPUT29), .ZN(n641) );
  INV_X1 U565 ( .A(KEYINPUT71), .ZN(n602) );
  OR2_X1 U566 ( .A1(G1384), .A2(n753), .ZN(n585) );
  XNOR2_X1 U567 ( .A(n603), .B(n602), .ZN(n604) );
  XNOR2_X1 U568 ( .A(n607), .B(KEYINPUT13), .ZN(n609) );
  NAND2_X1 U569 ( .A1(G101), .A2(n975), .ZN(n519) );
  INV_X1 U570 ( .A(G2104), .ZN(n518) );
  NAND2_X1 U571 ( .A1(n982), .A2(G125), .ZN(n521) );
  XOR2_X1 U572 ( .A(KEYINPUT23), .B(n519), .Z(n520) );
  NAND2_X1 U573 ( .A1(n521), .A2(n520), .ZN(n526) );
  NOR2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XOR2_X2 U575 ( .A(KEYINPUT17), .B(n522), .Z(n974) );
  NAND2_X1 U576 ( .A1(G137), .A2(n974), .ZN(n524) );
  AND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n979) );
  NAND2_X1 U578 ( .A1(G113), .A2(n979), .ZN(n523) );
  NAND2_X1 U579 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X2 U580 ( .A1(n526), .A2(n525), .ZN(G160) );
  XNOR2_X1 U581 ( .A(G543), .B(KEYINPUT0), .ZN(n527) );
  XNOR2_X1 U582 ( .A(n527), .B(KEYINPUT65), .ZN(n560) );
  NOR2_X2 U583 ( .A1(n560), .A2(G651), .ZN(n785) );
  NAND2_X1 U584 ( .A1(G52), .A2(n785), .ZN(n530) );
  XOR2_X1 U585 ( .A(G651), .B(KEYINPUT66), .Z(n532) );
  NOR2_X1 U586 ( .A1(G543), .A2(n532), .ZN(n528) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n528), .Z(n610) );
  BUF_X1 U588 ( .A(n610), .Z(n781) );
  NAND2_X1 U589 ( .A1(G64), .A2(n781), .ZN(n529) );
  NAND2_X1 U590 ( .A1(n530), .A2(n529), .ZN(n538) );
  NAND2_X1 U591 ( .A1(n782), .A2(G90), .ZN(n531) );
  XOR2_X1 U592 ( .A(KEYINPUT69), .B(n531), .Z(n535) );
  OR2_X1 U593 ( .A1(n560), .A2(n532), .ZN(n533) );
  XNOR2_X2 U594 ( .A(KEYINPUT67), .B(n533), .ZN(n780) );
  NAND2_X1 U595 ( .A1(n780), .A2(G77), .ZN(n534) );
  NAND2_X1 U596 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U597 ( .A(KEYINPUT9), .B(n536), .Z(n537) );
  NOR2_X1 U598 ( .A1(n538), .A2(n537), .ZN(G171) );
  NAND2_X1 U599 ( .A1(G51), .A2(n785), .ZN(n540) );
  NAND2_X1 U600 ( .A1(G63), .A2(n781), .ZN(n539) );
  NAND2_X1 U601 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U602 ( .A(KEYINPUT6), .B(n541), .ZN(n548) );
  NAND2_X1 U603 ( .A1(n782), .A2(G89), .ZN(n542) );
  XNOR2_X1 U604 ( .A(n542), .B(KEYINPUT4), .ZN(n544) );
  NAND2_X1 U605 ( .A1(G76), .A2(n780), .ZN(n543) );
  NAND2_X1 U606 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U607 ( .A(KEYINPUT5), .B(n545), .Z(n546) );
  XNOR2_X1 U608 ( .A(KEYINPUT76), .B(n546), .ZN(n547) );
  NOR2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U610 ( .A(KEYINPUT7), .B(n549), .Z(G168) );
  XOR2_X1 U611 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U612 ( .A1(G50), .A2(n785), .ZN(n551) );
  NAND2_X1 U613 ( .A1(G88), .A2(n782), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n555) );
  NAND2_X1 U615 ( .A1(G62), .A2(n781), .ZN(n553) );
  NAND2_X1 U616 ( .A1(G75), .A2(n780), .ZN(n552) );
  NAND2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U618 ( .A1(n555), .A2(n554), .ZN(G166) );
  NAND2_X1 U619 ( .A1(G49), .A2(n785), .ZN(n557) );
  NAND2_X1 U620 ( .A1(G74), .A2(G651), .ZN(n556) );
  NAND2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U622 ( .A(KEYINPUT81), .B(n558), .Z(n559) );
  NOR2_X1 U623 ( .A1(n781), .A2(n559), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n560), .A2(G87), .ZN(n561) );
  NAND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(G288) );
  INV_X1 U626 ( .A(G166), .ZN(G303) );
  NAND2_X1 U627 ( .A1(G73), .A2(n780), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT2), .B(n563), .Z(n569) );
  NAND2_X1 U629 ( .A1(n782), .A2(G86), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT82), .ZN(n566) );
  NAND2_X1 U631 ( .A1(G61), .A2(n781), .ZN(n565) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT83), .B(n567), .Z(n568) );
  NOR2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n785), .A2(G48), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(G305) );
  NAND2_X1 U637 ( .A1(n781), .A2(G60), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n785), .A2(G47), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT68), .B(n574), .Z(n578) );
  NAND2_X1 U641 ( .A1(G85), .A2(n782), .ZN(n576) );
  NAND2_X1 U642 ( .A1(G72), .A2(n780), .ZN(n575) );
  AND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(G290) );
  INV_X1 U645 ( .A(G1384), .ZN(n579) );
  AND2_X1 U646 ( .A1(G138), .A2(n579), .ZN(n580) );
  NAND2_X1 U647 ( .A1(n974), .A2(n580), .ZN(n586) );
  AND2_X1 U648 ( .A1(G102), .A2(n975), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G126), .A2(n982), .ZN(n582) );
  NAND2_X1 U650 ( .A1(G114), .A2(n979), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n753) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n715) );
  NAND2_X2 U654 ( .A1(n587), .A2(G160), .ZN(n667) );
  NOR2_X1 U655 ( .A1(G2084), .A2(n667), .ZN(n649) );
  NAND2_X1 U656 ( .A1(G8), .A2(n649), .ZN(n663) );
  NAND2_X1 U657 ( .A1(G8), .A2(n667), .ZN(n701) );
  NOR2_X1 U658 ( .A1(G1966), .A2(n701), .ZN(n661) );
  NAND2_X1 U659 ( .A1(G79), .A2(n780), .ZN(n594) );
  NAND2_X1 U660 ( .A1(G66), .A2(n610), .ZN(n589) );
  NAND2_X1 U661 ( .A1(G92), .A2(n782), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U663 ( .A1(G54), .A2(n785), .ZN(n590) );
  XNOR2_X1 U664 ( .A(KEYINPUT73), .B(n590), .ZN(n591) );
  NOR2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U667 ( .A(n595), .B(KEYINPUT15), .ZN(n1003) );
  INV_X1 U668 ( .A(n1003), .ZN(n758) );
  INV_X1 U669 ( .A(G1996), .ZN(n596) );
  XOR2_X1 U670 ( .A(KEYINPUT26), .B(KEYINPUT92), .Z(n597) );
  XNOR2_X1 U671 ( .A(n598), .B(n597), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n667), .A2(G1341), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U674 ( .A1(G81), .A2(n782), .ZN(n603) );
  XNOR2_X1 U675 ( .A(n604), .B(KEYINPUT12), .ZN(n606) );
  NAND2_X1 U676 ( .A1(G68), .A2(n780), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U678 ( .A1(G43), .A2(n785), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U680 ( .A1(n610), .A2(G56), .ZN(n611) );
  XOR2_X1 U681 ( .A(KEYINPUT14), .B(n611), .Z(n612) );
  NAND2_X1 U682 ( .A1(n614), .A2(n1006), .ZN(n615) );
  XNOR2_X1 U683 ( .A(n615), .B(KEYINPUT64), .ZN(n621) );
  OR2_X2 U684 ( .A1(n758), .A2(n621), .ZN(n619) );
  INV_X1 U685 ( .A(n667), .ZN(n643) );
  NOR2_X1 U686 ( .A1(n643), .A2(G1348), .ZN(n617) );
  NOR2_X1 U687 ( .A1(G2067), .A2(n667), .ZN(n616) );
  NOR2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U690 ( .A(n620), .B(KEYINPUT94), .ZN(n634) );
  NAND2_X1 U691 ( .A1(n621), .A2(n758), .ZN(n632) );
  NAND2_X1 U692 ( .A1(G53), .A2(n785), .ZN(n623) );
  NAND2_X1 U693 ( .A1(G78), .A2(n780), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U695 ( .A1(G65), .A2(n781), .ZN(n625) );
  NAND2_X1 U696 ( .A1(G91), .A2(n782), .ZN(n624) );
  NAND2_X1 U697 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U698 ( .A1(n627), .A2(n626), .ZN(n795) );
  NAND2_X1 U699 ( .A1(n643), .A2(G2072), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n628), .B(KEYINPUT27), .ZN(n630) );
  INV_X1 U701 ( .A(G1956), .ZN(n830) );
  NOR2_X1 U702 ( .A1(n830), .A2(n643), .ZN(n629) );
  NOR2_X1 U703 ( .A1(n630), .A2(n629), .ZN(n636) );
  NOR2_X1 U704 ( .A1(n795), .A2(n636), .ZN(n631) );
  XOR2_X1 U705 ( .A(n631), .B(KEYINPUT28), .Z(n635) );
  AND2_X1 U706 ( .A1(n632), .A2(n635), .ZN(n633) );
  AND2_X1 U707 ( .A1(n634), .A2(n633), .ZN(n640) );
  INV_X1 U708 ( .A(n635), .ZN(n638) );
  NAND2_X1 U709 ( .A1(n795), .A2(n636), .ZN(n637) );
  NOR2_X1 U710 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n642), .B(n641), .ZN(n648) );
  XOR2_X1 U713 ( .A(G2078), .B(KEYINPUT25), .Z(n861) );
  NOR2_X1 U714 ( .A1(n861), .A2(n667), .ZN(n645) );
  NOR2_X1 U715 ( .A1(n643), .A2(G1961), .ZN(n644) );
  NOR2_X1 U716 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U717 ( .A(KEYINPUT91), .B(n646), .ZN(n654) );
  NAND2_X1 U718 ( .A1(n654), .A2(G171), .ZN(n647) );
  NAND2_X1 U719 ( .A1(n648), .A2(n647), .ZN(n659) );
  NOR2_X1 U720 ( .A1(n661), .A2(n649), .ZN(n650) );
  XOR2_X1 U721 ( .A(KEYINPUT95), .B(n650), .Z(n651) );
  NAND2_X1 U722 ( .A1(G8), .A2(n651), .ZN(n652) );
  XNOR2_X1 U723 ( .A(KEYINPUT30), .B(n652), .ZN(n653) );
  NOR2_X1 U724 ( .A1(G168), .A2(n653), .ZN(n656) );
  NOR2_X1 U725 ( .A1(G171), .A2(n654), .ZN(n655) );
  NOR2_X1 U726 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U727 ( .A(KEYINPUT31), .B(n657), .Z(n658) );
  NAND2_X1 U728 ( .A1(n659), .A2(n658), .ZN(n665) );
  XOR2_X1 U729 ( .A(KEYINPUT96), .B(n665), .Z(n660) );
  NOR2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n694) );
  AND2_X1 U732 ( .A1(G286), .A2(G8), .ZN(n664) );
  NAND2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n675) );
  INV_X1 U734 ( .A(G8), .ZN(n673) );
  NOR2_X1 U735 ( .A1(G1971), .A2(n701), .ZN(n666) );
  XNOR2_X1 U736 ( .A(KEYINPUT97), .B(n666), .ZN(n670) );
  NOR2_X1 U737 ( .A1(G2090), .A2(n667), .ZN(n668) );
  NOR2_X1 U738 ( .A1(G166), .A2(n668), .ZN(n669) );
  NAND2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U740 ( .A(n671), .B(KEYINPUT98), .ZN(n672) );
  OR2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n674) );
  INV_X1 U742 ( .A(KEYINPUT33), .ZN(n677) );
  NAND2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n927) );
  AND2_X1 U744 ( .A1(n677), .A2(n927), .ZN(n678) );
  INV_X1 U745 ( .A(n701), .ZN(n683) );
  AND2_X1 U746 ( .A1(n678), .A2(n683), .ZN(n680) );
  AND2_X1 U747 ( .A1(n693), .A2(n680), .ZN(n679) );
  NAND2_X1 U748 ( .A1(n694), .A2(n679), .ZN(n689) );
  INV_X1 U749 ( .A(n680), .ZN(n682) );
  NOR2_X1 U750 ( .A1(G1976), .A2(G288), .ZN(n684) );
  NOR2_X1 U751 ( .A1(G1971), .A2(G303), .ZN(n681) );
  NOR2_X1 U752 ( .A1(n684), .A2(n681), .ZN(n924) );
  OR2_X1 U753 ( .A1(n682), .A2(n924), .ZN(n687) );
  NAND2_X1 U754 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U755 ( .A1(n685), .A2(KEYINPUT33), .ZN(n686) );
  AND2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U758 ( .A(n690), .B(KEYINPUT99), .ZN(n691) );
  XNOR2_X1 U759 ( .A(G1981), .B(G305), .ZN(n919) );
  NOR2_X1 U760 ( .A1(n691), .A2(n919), .ZN(n692) );
  INV_X1 U761 ( .A(n692), .ZN(n704) );
  NAND2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n697) );
  NOR2_X1 U763 ( .A1(G2090), .A2(G303), .ZN(n695) );
  NAND2_X1 U764 ( .A1(G8), .A2(n695), .ZN(n696) );
  NAND2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U766 ( .A1(n701), .A2(n698), .ZN(n702) );
  NOR2_X1 U767 ( .A1(G1981), .A2(G305), .ZN(n699) );
  XOR2_X1 U768 ( .A(n699), .B(KEYINPUT24), .Z(n700) );
  NAND2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n736) );
  NAND2_X1 U770 ( .A1(n975), .A2(G104), .ZN(n705) );
  XNOR2_X1 U771 ( .A(n705), .B(KEYINPUT88), .ZN(n707) );
  NAND2_X1 U772 ( .A1(G140), .A2(n974), .ZN(n706) );
  NAND2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U774 ( .A(KEYINPUT34), .B(n708), .ZN(n713) );
  NAND2_X1 U775 ( .A1(G128), .A2(n982), .ZN(n710) );
  NAND2_X1 U776 ( .A1(G116), .A2(n979), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U778 ( .A(KEYINPUT35), .B(n711), .Z(n712) );
  NOR2_X1 U779 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U780 ( .A(KEYINPUT36), .B(n714), .ZN(n999) );
  XNOR2_X1 U781 ( .A(G2067), .B(KEYINPUT37), .ZN(n746) );
  NOR2_X1 U782 ( .A1(n999), .A2(n746), .ZN(n904) );
  NAND2_X1 U783 ( .A1(G160), .A2(G40), .ZN(n716) );
  NOR2_X1 U784 ( .A1(n715), .A2(n716), .ZN(n748) );
  NAND2_X1 U785 ( .A1(n904), .A2(n748), .ZN(n717) );
  XOR2_X1 U786 ( .A(KEYINPUT89), .B(n717), .Z(n744) );
  INV_X1 U787 ( .A(n744), .ZN(n734) );
  NAND2_X1 U788 ( .A1(G141), .A2(n974), .ZN(n719) );
  NAND2_X1 U789 ( .A1(G129), .A2(n982), .ZN(n718) );
  NAND2_X1 U790 ( .A1(n719), .A2(n718), .ZN(n722) );
  NAND2_X1 U791 ( .A1(n975), .A2(G105), .ZN(n720) );
  XOR2_X1 U792 ( .A(KEYINPUT38), .B(n720), .Z(n721) );
  NOR2_X1 U793 ( .A1(n722), .A2(n721), .ZN(n724) );
  NAND2_X1 U794 ( .A1(n979), .A2(G117), .ZN(n723) );
  NAND2_X1 U795 ( .A1(n724), .A2(n723), .ZN(n989) );
  NAND2_X1 U796 ( .A1(G1996), .A2(n989), .ZN(n725) );
  XNOR2_X1 U797 ( .A(n725), .B(KEYINPUT90), .ZN(n733) );
  NAND2_X1 U798 ( .A1(G131), .A2(n974), .ZN(n727) );
  NAND2_X1 U799 ( .A1(G95), .A2(n975), .ZN(n726) );
  NAND2_X1 U800 ( .A1(n727), .A2(n726), .ZN(n731) );
  NAND2_X1 U801 ( .A1(G119), .A2(n982), .ZN(n729) );
  NAND2_X1 U802 ( .A1(G107), .A2(n979), .ZN(n728) );
  NAND2_X1 U803 ( .A1(n729), .A2(n728), .ZN(n730) );
  OR2_X1 U804 ( .A1(n731), .A2(n730), .ZN(n990) );
  NAND2_X1 U805 ( .A1(G1991), .A2(n990), .ZN(n732) );
  NAND2_X1 U806 ( .A1(n733), .A2(n732), .ZN(n900) );
  XNOR2_X1 U807 ( .A(n515), .B(KEYINPUT100), .ZN(n739) );
  XNOR2_X1 U808 ( .A(G1986), .B(G290), .ZN(n926) );
  NAND2_X1 U809 ( .A1(n748), .A2(n926), .ZN(n737) );
  XOR2_X1 U810 ( .A(KEYINPUT87), .B(n737), .Z(n738) );
  NAND2_X1 U811 ( .A1(n739), .A2(n738), .ZN(n751) );
  NOR2_X1 U812 ( .A1(G1996), .A2(n989), .ZN(n894) );
  NOR2_X1 U813 ( .A1(G1986), .A2(G290), .ZN(n740) );
  NOR2_X1 U814 ( .A1(G1991), .A2(n990), .ZN(n898) );
  NOR2_X1 U815 ( .A1(n740), .A2(n898), .ZN(n741) );
  NOR2_X1 U816 ( .A1(n900), .A2(n741), .ZN(n742) );
  NOR2_X1 U817 ( .A1(n894), .A2(n742), .ZN(n743) );
  XNOR2_X1 U818 ( .A(KEYINPUT39), .B(n743), .ZN(n745) );
  NAND2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n747) );
  NAND2_X1 U820 ( .A1(n999), .A2(n746), .ZN(n907) );
  NAND2_X1 U821 ( .A1(n747), .A2(n907), .ZN(n749) );
  NAND2_X1 U822 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U823 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U824 ( .A(n752), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U825 ( .A1(G138), .A2(n974), .ZN(n754) );
  AND2_X1 U826 ( .A1(n754), .A2(n753), .ZN(G164) );
  AND2_X1 U827 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U828 ( .A(n795), .ZN(G299) );
  INV_X1 U829 ( .A(G57), .ZN(G237) );
  INV_X1 U830 ( .A(G132), .ZN(G219) );
  INV_X1 U831 ( .A(G82), .ZN(G220) );
  NAND2_X1 U832 ( .A1(G7), .A2(G661), .ZN(n755) );
  XNOR2_X1 U833 ( .A(n755), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U834 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n757) );
  INV_X1 U835 ( .A(G223), .ZN(n817) );
  NAND2_X1 U836 ( .A1(G567), .A2(n817), .ZN(n756) );
  XNOR2_X1 U837 ( .A(n757), .B(n756), .ZN(G234) );
  NAND2_X1 U838 ( .A1(n1006), .A2(G860), .ZN(G153) );
  XOR2_X1 U839 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  INV_X1 U840 ( .A(G868), .ZN(n801) );
  NAND2_X1 U841 ( .A1(n758), .A2(n801), .ZN(n759) );
  XNOR2_X1 U842 ( .A(n759), .B(KEYINPUT74), .ZN(n761) );
  NAND2_X1 U843 ( .A1(G301), .A2(G868), .ZN(n760) );
  NAND2_X1 U844 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U845 ( .A(KEYINPUT75), .B(n762), .Z(G284) );
  NOR2_X1 U846 ( .A1(G286), .A2(n801), .ZN(n764) );
  NOR2_X1 U847 ( .A1(G868), .A2(G299), .ZN(n763) );
  NOR2_X1 U848 ( .A1(n764), .A2(n763), .ZN(G297) );
  INV_X1 U849 ( .A(G860), .ZN(n944) );
  NAND2_X1 U850 ( .A1(n944), .A2(G559), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n765), .A2(n1003), .ZN(n766) );
  XNOR2_X1 U852 ( .A(n766), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U853 ( .A1(n1003), .A2(G868), .ZN(n767) );
  NOR2_X1 U854 ( .A1(G559), .A2(n767), .ZN(n769) );
  AND2_X1 U855 ( .A1(n801), .A2(n1006), .ZN(n768) );
  NOR2_X1 U856 ( .A1(n769), .A2(n768), .ZN(G282) );
  XNOR2_X1 U857 ( .A(G2100), .B(KEYINPUT77), .ZN(n778) );
  NAND2_X1 U858 ( .A1(G123), .A2(n982), .ZN(n770) );
  XNOR2_X1 U859 ( .A(n770), .B(KEYINPUT18), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n975), .A2(G99), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n776) );
  NAND2_X1 U862 ( .A1(G135), .A2(n974), .ZN(n774) );
  NAND2_X1 U863 ( .A1(G111), .A2(n979), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n987) );
  XNOR2_X1 U866 ( .A(n987), .B(G2096), .ZN(n777) );
  NAND2_X1 U867 ( .A1(n778), .A2(n777), .ZN(G156) );
  NAND2_X1 U868 ( .A1(G559), .A2(n1003), .ZN(n779) );
  XNOR2_X1 U869 ( .A(n779), .B(n1006), .ZN(n943) );
  NAND2_X1 U870 ( .A1(G80), .A2(n780), .ZN(n790) );
  NAND2_X1 U871 ( .A1(G67), .A2(n781), .ZN(n784) );
  NAND2_X1 U872 ( .A1(G93), .A2(n782), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U874 ( .A1(G55), .A2(n785), .ZN(n786) );
  XNOR2_X1 U875 ( .A(KEYINPUT79), .B(n786), .ZN(n787) );
  NOR2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U878 ( .A(n791), .B(KEYINPUT80), .ZN(n947) );
  XNOR2_X1 U879 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n793) );
  XNOR2_X1 U880 ( .A(G290), .B(KEYINPUT19), .ZN(n792) );
  XNOR2_X1 U881 ( .A(n793), .B(n792), .ZN(n794) );
  XNOR2_X1 U882 ( .A(G288), .B(n794), .ZN(n797) );
  XNOR2_X1 U883 ( .A(n795), .B(G166), .ZN(n796) );
  XNOR2_X1 U884 ( .A(n797), .B(n796), .ZN(n798) );
  XOR2_X1 U885 ( .A(n947), .B(n798), .Z(n799) );
  XNOR2_X1 U886 ( .A(G305), .B(n799), .ZN(n1002) );
  XNOR2_X1 U887 ( .A(n943), .B(n1002), .ZN(n800) );
  NAND2_X1 U888 ( .A1(n800), .A2(G868), .ZN(n803) );
  NAND2_X1 U889 ( .A1(n801), .A2(n947), .ZN(n802) );
  NAND2_X1 U890 ( .A1(n803), .A2(n802), .ZN(G295) );
  NAND2_X1 U891 ( .A1(G2084), .A2(G2078), .ZN(n804) );
  XOR2_X1 U892 ( .A(KEYINPUT20), .B(n804), .Z(n805) );
  NAND2_X1 U893 ( .A1(G2090), .A2(n805), .ZN(n806) );
  XNOR2_X1 U894 ( .A(KEYINPUT21), .B(n806), .ZN(n807) );
  NAND2_X1 U895 ( .A1(n807), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U896 ( .A(KEYINPUT86), .B(G44), .ZN(n808) );
  XNOR2_X1 U897 ( .A(n808), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U898 ( .A1(G220), .A2(G219), .ZN(n809) );
  XOR2_X1 U899 ( .A(KEYINPUT22), .B(n809), .Z(n810) );
  NOR2_X1 U900 ( .A1(G218), .A2(n810), .ZN(n811) );
  NAND2_X1 U901 ( .A1(G96), .A2(n811), .ZN(n941) );
  NAND2_X1 U902 ( .A1(n941), .A2(G2106), .ZN(n815) );
  NAND2_X1 U903 ( .A1(G120), .A2(G108), .ZN(n812) );
  NOR2_X1 U904 ( .A1(G237), .A2(n812), .ZN(n813) );
  NAND2_X1 U905 ( .A1(G69), .A2(n813), .ZN(n942) );
  NAND2_X1 U906 ( .A1(n942), .A2(G567), .ZN(n814) );
  NAND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n948) );
  NAND2_X1 U908 ( .A1(G661), .A2(G483), .ZN(n816) );
  NOR2_X1 U909 ( .A1(n948), .A2(n816), .ZN(n820) );
  NAND2_X1 U910 ( .A1(n820), .A2(G36), .ZN(G176) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n817), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n818) );
  NAND2_X1 U913 ( .A1(G661), .A2(n818), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(G188) );
  XNOR2_X1 U916 ( .A(G108), .B(KEYINPUT115), .ZN(G238) );
  NAND2_X1 U918 ( .A1(G124), .A2(n982), .ZN(n821) );
  XNOR2_X1 U919 ( .A(n821), .B(KEYINPUT44), .ZN(n824) );
  NAND2_X1 U920 ( .A1(G100), .A2(n975), .ZN(n822) );
  XOR2_X1 U921 ( .A(KEYINPUT109), .B(n822), .Z(n823) );
  NAND2_X1 U922 ( .A1(n824), .A2(n823), .ZN(n828) );
  NAND2_X1 U923 ( .A1(G136), .A2(n974), .ZN(n826) );
  NAND2_X1 U924 ( .A1(G112), .A2(n979), .ZN(n825) );
  NAND2_X1 U925 ( .A1(n826), .A2(n825), .ZN(n827) );
  NOR2_X1 U926 ( .A1(n828), .A2(n827), .ZN(G162) );
  XOR2_X1 U927 ( .A(G1348), .B(KEYINPUT59), .Z(n829) );
  XNOR2_X1 U928 ( .A(G4), .B(n829), .ZN(n838) );
  XNOR2_X1 U929 ( .A(G20), .B(n830), .ZN(n833) );
  XOR2_X1 U930 ( .A(G1341), .B(G19), .Z(n831) );
  XNOR2_X1 U931 ( .A(KEYINPUT124), .B(n831), .ZN(n832) );
  NAND2_X1 U932 ( .A1(n833), .A2(n832), .ZN(n835) );
  XNOR2_X1 U933 ( .A(G6), .B(G1981), .ZN(n834) );
  NOR2_X1 U934 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n836), .B(KEYINPUT125), .ZN(n837) );
  NOR2_X1 U936 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U937 ( .A(KEYINPUT60), .B(n839), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n840), .B(KEYINPUT126), .ZN(n844) );
  XNOR2_X1 U939 ( .A(G1966), .B(G21), .ZN(n842) );
  XNOR2_X1 U940 ( .A(G5), .B(G1961), .ZN(n841) );
  NOR2_X1 U941 ( .A1(n842), .A2(n841), .ZN(n843) );
  NAND2_X1 U942 ( .A1(n844), .A2(n843), .ZN(n851) );
  XNOR2_X1 U943 ( .A(G1986), .B(G24), .ZN(n846) );
  XNOR2_X1 U944 ( .A(G1971), .B(G22), .ZN(n845) );
  NOR2_X1 U945 ( .A1(n846), .A2(n845), .ZN(n848) );
  XOR2_X1 U946 ( .A(G1976), .B(G23), .Z(n847) );
  NAND2_X1 U947 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U948 ( .A(KEYINPUT58), .B(n849), .ZN(n850) );
  NOR2_X1 U949 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U950 ( .A(KEYINPUT61), .B(n852), .ZN(n854) );
  INV_X1 U951 ( .A(G16), .ZN(n853) );
  NAND2_X1 U952 ( .A1(n854), .A2(n853), .ZN(n855) );
  NAND2_X1 U953 ( .A1(n855), .A2(G11), .ZN(n880) );
  XNOR2_X1 U954 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n911) );
  XNOR2_X1 U955 ( .A(G2090), .B(G35), .ZN(n872) );
  XNOR2_X1 U956 ( .A(G2067), .B(G26), .ZN(n857) );
  XNOR2_X1 U957 ( .A(G2072), .B(G33), .ZN(n856) );
  NOR2_X1 U958 ( .A1(n857), .A2(n856), .ZN(n866) );
  XOR2_X1 U959 ( .A(G1991), .B(G25), .Z(n858) );
  XNOR2_X1 U960 ( .A(KEYINPUT118), .B(n858), .ZN(n859) );
  NAND2_X1 U961 ( .A1(G28), .A2(n859), .ZN(n860) );
  XOR2_X1 U962 ( .A(KEYINPUT119), .B(n860), .Z(n864) );
  XNOR2_X1 U963 ( .A(G27), .B(n861), .ZN(n862) );
  XNOR2_X1 U964 ( .A(KEYINPUT120), .B(n862), .ZN(n863) );
  NOR2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n869) );
  XOR2_X1 U967 ( .A(KEYINPUT121), .B(G1996), .Z(n867) );
  XNOR2_X1 U968 ( .A(G32), .B(n867), .ZN(n868) );
  NOR2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U970 ( .A(KEYINPUT53), .B(n870), .ZN(n871) );
  NOR2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n875) );
  XOR2_X1 U972 ( .A(G2084), .B(G34), .Z(n873) );
  XNOR2_X1 U973 ( .A(KEYINPUT54), .B(n873), .ZN(n874) );
  NAND2_X1 U974 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U975 ( .A(n911), .B(n876), .Z(n877) );
  NOR2_X1 U976 ( .A1(G29), .A2(n877), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n878), .B(KEYINPUT122), .ZN(n879) );
  NOR2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n915) );
  NAND2_X1 U979 ( .A1(n975), .A2(G103), .ZN(n881) );
  XNOR2_X1 U980 ( .A(KEYINPUT111), .B(n881), .ZN(n889) );
  NAND2_X1 U981 ( .A1(G127), .A2(n982), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G115), .A2(n979), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n884), .B(KEYINPUT112), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n885), .B(KEYINPUT47), .ZN(n887) );
  NAND2_X1 U986 ( .A1(n974), .A2(G139), .ZN(n886) );
  NAND2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n888) );
  NOR2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n973) );
  XOR2_X1 U989 ( .A(G2072), .B(n973), .Z(n891) );
  XOR2_X1 U990 ( .A(G164), .B(G2078), .Z(n890) );
  NOR2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U992 ( .A(KEYINPUT50), .B(n892), .ZN(n897) );
  XOR2_X1 U993 ( .A(G2090), .B(G162), .Z(n893) );
  NOR2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U995 ( .A(KEYINPUT51), .B(n895), .Z(n896) );
  NAND2_X1 U996 ( .A1(n897), .A2(n896), .ZN(n909) );
  NOR2_X1 U997 ( .A1(n898), .A2(n987), .ZN(n902) );
  XOR2_X1 U998 ( .A(G160), .B(G2084), .Z(n899) );
  NOR2_X1 U999 ( .A1(n900), .A2(n899), .ZN(n901) );
  NAND2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n903) );
  NOR2_X1 U1001 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n905), .B(KEYINPUT116), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(n907), .A2(n906), .ZN(n908) );
  NOR2_X1 U1004 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(KEYINPUT52), .B(n910), .ZN(n912) );
  NAND2_X1 U1006 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1007 ( .A1(n913), .A2(G29), .ZN(n914) );
  NAND2_X1 U1008 ( .A1(n915), .A2(n914), .ZN(n939) );
  XOR2_X1 U1009 ( .A(G16), .B(KEYINPUT56), .Z(n937) );
  XNOR2_X1 U1010 ( .A(G1341), .B(n1006), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(n1003), .B(G1348), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(n934) );
  XOR2_X1 U1013 ( .A(G168), .B(G1966), .Z(n918) );
  NOR2_X1 U1014 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1015 ( .A(KEYINPUT57), .B(n920), .Z(n932) );
  XNOR2_X1 U1016 ( .A(G299), .B(G1956), .ZN(n922) );
  AND2_X1 U1017 ( .A1(G1971), .A2(G303), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1020 ( .A1(n926), .A2(n925), .ZN(n928) );
  NAND2_X1 U1021 ( .A1(n928), .A2(n927), .ZN(n930) );
  XOR2_X1 U1022 ( .A(G171), .B(G1961), .Z(n929) );
  NOR2_X1 U1023 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1024 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1025 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1026 ( .A(KEYINPUT123), .B(n935), .Z(n936) );
  NOR2_X1 U1027 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1028 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1029 ( .A(n940), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1030 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1031 ( .A(G120), .ZN(G236) );
  INV_X1 U1032 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1033 ( .A1(n942), .A2(n941), .ZN(G325) );
  INV_X1 U1034 ( .A(G325), .ZN(G261) );
  NAND2_X1 U1035 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1036 ( .A(n945), .B(KEYINPUT78), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(n947), .B(n946), .ZN(G145) );
  INV_X1 U1038 ( .A(n948), .ZN(G319) );
  XOR2_X1 U1039 ( .A(KEYINPUT42), .B(KEYINPUT103), .Z(n950) );
  XNOR2_X1 U1040 ( .A(KEYINPUT104), .B(G2678), .ZN(n949) );
  XNOR2_X1 U1041 ( .A(n950), .B(n949), .ZN(n951) );
  XOR2_X1 U1042 ( .A(n951), .B(G2096), .Z(n953) );
  XNOR2_X1 U1043 ( .A(G2084), .B(G2072), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(n953), .B(n952), .ZN(n957) );
  XOR2_X1 U1045 ( .A(KEYINPUT43), .B(G2100), .Z(n955) );
  XNOR2_X1 U1046 ( .A(G2090), .B(KEYINPUT102), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(n955), .B(n954), .ZN(n956) );
  XOR2_X1 U1048 ( .A(n957), .B(n956), .Z(n959) );
  XNOR2_X1 U1049 ( .A(G2067), .B(G2078), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(n959), .B(n958), .ZN(G227) );
  XOR2_X1 U1051 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n961) );
  XNOR2_X1 U1052 ( .A(G1996), .B(G1991), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(n961), .B(n960), .ZN(n962) );
  XOR2_X1 U1054 ( .A(n962), .B(KEYINPUT105), .Z(n964) );
  XNOR2_X1 U1055 ( .A(G1961), .B(G1956), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(n964), .B(n963), .ZN(n972) );
  XOR2_X1 U1057 ( .A(KEYINPUT41), .B(G2474), .Z(n966) );
  XNOR2_X1 U1058 ( .A(G1971), .B(G1981), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(n966), .B(n965), .ZN(n970) );
  XOR2_X1 U1060 ( .A(KEYINPUT106), .B(G1976), .Z(n968) );
  XNOR2_X1 U1061 ( .A(G1986), .B(G1966), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(n968), .B(n967), .ZN(n969) );
  XOR2_X1 U1063 ( .A(n970), .B(n969), .Z(n971) );
  XNOR2_X1 U1064 ( .A(n972), .B(n971), .ZN(G229) );
  XNOR2_X1 U1065 ( .A(G160), .B(n973), .ZN(n998) );
  NAND2_X1 U1066 ( .A1(G142), .A2(n974), .ZN(n977) );
  NAND2_X1 U1067 ( .A1(G106), .A2(n975), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(n978), .B(KEYINPUT45), .ZN(n981) );
  NAND2_X1 U1070 ( .A1(G118), .A2(n979), .ZN(n980) );
  NAND2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n985) );
  NAND2_X1 U1072 ( .A1(n982), .A2(G130), .ZN(n983) );
  XOR2_X1 U1073 ( .A(KEYINPUT110), .B(n983), .Z(n984) );
  NOR2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1075 ( .A(n987), .B(n986), .Z(n988) );
  XNOR2_X1 U1076 ( .A(n989), .B(n988), .ZN(n994) );
  XNOR2_X1 U1077 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n992) );
  XNOR2_X1 U1078 ( .A(n990), .B(KEYINPUT46), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(n992), .B(n991), .ZN(n993) );
  XOR2_X1 U1080 ( .A(n994), .B(n993), .Z(n996) );
  XNOR2_X1 U1081 ( .A(G164), .B(G162), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(n996), .B(n995), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(n998), .B(n997), .ZN(n1000) );
  XOR2_X1 U1084 ( .A(n1000), .B(n999), .Z(n1001) );
  NOR2_X1 U1085 ( .A1(G37), .A2(n1001), .ZN(G395) );
  XOR2_X1 U1086 ( .A(KEYINPUT114), .B(n1002), .Z(n1005) );
  XNOR2_X1 U1087 ( .A(n1003), .B(G286), .ZN(n1004) );
  XNOR2_X1 U1088 ( .A(n1005), .B(n1004), .ZN(n1008) );
  XNOR2_X1 U1089 ( .A(n1006), .B(G171), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(n1008), .B(n1007), .ZN(n1009) );
  NOR2_X1 U1091 ( .A1(G37), .A2(n1009), .ZN(G397) );
  XOR2_X1 U1092 ( .A(G2443), .B(G2454), .Z(n1011) );
  XNOR2_X1 U1093 ( .A(G1341), .B(G2435), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(n1011), .B(n1010), .ZN(n1018) );
  XOR2_X1 U1095 ( .A(KEYINPUT101), .B(G2446), .Z(n1013) );
  XNOR2_X1 U1096 ( .A(G1348), .B(G2430), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(n1013), .B(n1012), .ZN(n1014) );
  XOR2_X1 U1098 ( .A(n1014), .B(G2451), .Z(n1016) );
  XNOR2_X1 U1099 ( .A(G2438), .B(G2427), .ZN(n1015) );
  XNOR2_X1 U1100 ( .A(n1016), .B(n1015), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(n1018), .B(n1017), .ZN(n1019) );
  NAND2_X1 U1102 ( .A1(n1019), .A2(G14), .ZN(n1025) );
  NAND2_X1 U1103 ( .A1(G319), .A2(n1025), .ZN(n1022) );
  NOR2_X1 U1104 ( .A1(G227), .A2(G229), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(KEYINPUT49), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  NOR2_X1 U1107 ( .A1(G395), .A2(G397), .ZN(n1023) );
  NAND2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(G225) );
  INV_X1 U1109 ( .A(G225), .ZN(G308) );
  INV_X1 U1110 ( .A(G69), .ZN(G235) );
  INV_X1 U1111 ( .A(n1025), .ZN(G401) );
endmodule

