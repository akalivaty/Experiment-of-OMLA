

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U323 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n415) );
  XOR2_X1 U324 ( .A(G148GAT), .B(KEYINPUT69), .Z(n291) );
  XOR2_X1 U325 ( .A(n304), .B(n303), .Z(n292) );
  XNOR2_X1 U326 ( .A(n390), .B(n446), .ZN(n299) );
  XNOR2_X1 U327 ( .A(n378), .B(n291), .ZN(n357) );
  XNOR2_X1 U328 ( .A(n358), .B(n357), .ZN(n362) );
  INV_X1 U329 ( .A(KEYINPUT7), .ZN(n296) );
  XNOR2_X1 U330 ( .A(n305), .B(n292), .ZN(n306) );
  XNOR2_X1 U331 ( .A(n297), .B(n296), .ZN(n390) );
  XNOR2_X1 U332 ( .A(n307), .B(n306), .ZN(n410) );
  XNOR2_X1 U333 ( .A(n455), .B(KEYINPUT124), .ZN(n456) );
  XNOR2_X1 U334 ( .A(n461), .B(G176GAT), .ZN(n462) );
  XNOR2_X1 U335 ( .A(n457), .B(n456), .ZN(G1355GAT) );
  XNOR2_X1 U336 ( .A(n463), .B(n462), .ZN(G1349GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n294) );
  NAND2_X1 U338 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U340 ( .A(n295), .B(G92GAT), .Z(n300) );
  XOR2_X1 U341 ( .A(G43GAT), .B(KEYINPUT8), .Z(n297) );
  XNOR2_X1 U342 ( .A(G29GAT), .B(G134GAT), .ZN(n298) );
  XNOR2_X1 U343 ( .A(n298), .B(KEYINPUT70), .ZN(n446) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n302) );
  XNOR2_X1 U345 ( .A(G36GAT), .B(G190GAT), .ZN(n301) );
  XOR2_X1 U346 ( .A(n301), .B(G218GAT), .Z(n426) );
  XNOR2_X1 U347 ( .A(n302), .B(n426), .ZN(n307) );
  XOR2_X1 U348 ( .A(G50GAT), .B(G162GAT), .Z(n333) );
  XOR2_X1 U349 ( .A(G99GAT), .B(G85GAT), .Z(n354) );
  XNOR2_X1 U350 ( .A(n333), .B(n354), .ZN(n305) );
  XOR2_X1 U351 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n304) );
  XNOR2_X1 U352 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n303) );
  XOR2_X1 U353 ( .A(KEYINPUT36), .B(n410), .Z(n488) );
  XOR2_X1 U354 ( .A(KEYINPUT26), .B(KEYINPUT99), .Z(n351) );
  XOR2_X1 U355 ( .A(KEYINPUT79), .B(KEYINPUT20), .Z(n309) );
  XNOR2_X1 U356 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U358 ( .A(G120GAT), .B(G176GAT), .Z(n311) );
  XNOR2_X1 U359 ( .A(G134GAT), .B(G190GAT), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n330) );
  XOR2_X1 U362 ( .A(G99GAT), .B(G43GAT), .Z(n315) );
  NAND2_X1 U363 ( .A1(G227GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n318) );
  XOR2_X1 U365 ( .A(G127GAT), .B(KEYINPUT78), .Z(n317) );
  XNOR2_X1 U366 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n317), .B(n316), .ZN(n447) );
  XOR2_X1 U368 ( .A(n318), .B(n447), .Z(n328) );
  XOR2_X1 U369 ( .A(KEYINPUT18), .B(KEYINPUT82), .Z(n320) );
  XNOR2_X1 U370 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U372 ( .A(n321), .B(KEYINPUT83), .Z(n323) );
  XNOR2_X1 U373 ( .A(G169GAT), .B(G183GAT), .ZN(n322) );
  XNOR2_X1 U374 ( .A(n323), .B(n322), .ZN(n421) );
  XOR2_X1 U375 ( .A(G71GAT), .B(KEYINPUT81), .Z(n325) );
  XNOR2_X1 U376 ( .A(G15GAT), .B(KEYINPUT80), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n421), .B(n326), .ZN(n327) );
  XNOR2_X1 U379 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U380 ( .A(n330), .B(n329), .Z(n531) );
  INV_X1 U381 ( .A(n531), .ZN(n522) );
  XOR2_X1 U382 ( .A(KEYINPUT23), .B(KEYINPUT87), .Z(n332) );
  XNOR2_X1 U383 ( .A(KEYINPUT88), .B(KEYINPUT22), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n345) );
  XOR2_X1 U385 ( .A(KEYINPUT24), .B(G218GAT), .Z(n335) );
  XOR2_X1 U386 ( .A(G106GAT), .B(G78GAT), .Z(n363) );
  XNOR2_X1 U387 ( .A(n333), .B(n363), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U389 ( .A(n336), .B(G204GAT), .Z(n343) );
  XOR2_X1 U390 ( .A(G211GAT), .B(KEYINPUT86), .Z(n338) );
  XNOR2_X1 U391 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n425) );
  XOR2_X1 U393 ( .A(n425), .B(KEYINPUT89), .Z(n340) );
  NAND2_X1 U394 ( .A1(G228GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U396 ( .A(G22GAT), .B(n341), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U399 ( .A(KEYINPUT2), .B(G155GAT), .Z(n347) );
  XNOR2_X1 U400 ( .A(KEYINPUT3), .B(G148GAT), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U402 ( .A(G141GAT), .B(n348), .Z(n435) );
  XOR2_X1 U403 ( .A(n349), .B(n435), .Z(n466) );
  NAND2_X1 U404 ( .A1(n522), .A2(n466), .ZN(n350) );
  XOR2_X1 U405 ( .A(n351), .B(n350), .Z(n548) );
  INV_X1 U406 ( .A(n548), .ZN(n451) );
  XOR2_X1 U407 ( .A(G64GAT), .B(G92GAT), .Z(n353) );
  XNOR2_X1 U408 ( .A(G176GAT), .B(G204GAT), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n419) );
  XOR2_X1 U410 ( .A(n419), .B(n354), .Z(n356) );
  NAND2_X1 U411 ( .A1(G230GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n356), .B(n355), .ZN(n358) );
  XOR2_X1 U413 ( .A(G71GAT), .B(KEYINPUT13), .Z(n378) );
  XOR2_X1 U414 ( .A(KEYINPUT68), .B(KEYINPUT32), .Z(n360) );
  XNOR2_X1 U415 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U417 ( .A(n362), .B(n361), .Z(n365) );
  XOR2_X1 U418 ( .A(G120GAT), .B(G57GAT), .Z(n441) );
  XNOR2_X1 U419 ( .A(n363), .B(n441), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n574) );
  XOR2_X1 U421 ( .A(KEYINPUT72), .B(KEYINPUT75), .Z(n367) );
  XNOR2_X1 U422 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n386) );
  XOR2_X1 U424 ( .A(G78GAT), .B(G211GAT), .Z(n369) );
  XNOR2_X1 U425 ( .A(G183GAT), .B(G155GAT), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U427 ( .A(KEYINPUT76), .B(G64GAT), .Z(n371) );
  XNOR2_X1 U428 ( .A(G127GAT), .B(G57GAT), .ZN(n370) );
  XNOR2_X1 U429 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U430 ( .A(n373), .B(n372), .Z(n384) );
  XOR2_X1 U431 ( .A(KEYINPUT15), .B(KEYINPUT74), .Z(n375) );
  XNOR2_X1 U432 ( .A(KEYINPUT71), .B(KEYINPUT73), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n375), .B(n374), .ZN(n382) );
  XOR2_X1 U434 ( .A(G8GAT), .B(G1GAT), .Z(n377) );
  XNOR2_X1 U435 ( .A(G22GAT), .B(G15GAT), .ZN(n376) );
  XNOR2_X1 U436 ( .A(n377), .B(n376), .ZN(n391) );
  XOR2_X1 U437 ( .A(n378), .B(n391), .Z(n380) );
  NAND2_X1 U438 ( .A1(G231GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n578) );
  INV_X1 U443 ( .A(n578), .ZN(n556) );
  NOR2_X1 U444 ( .A1(n556), .A2(n488), .ZN(n387) );
  XOR2_X1 U445 ( .A(KEYINPUT45), .B(n387), .Z(n388) );
  NOR2_X1 U446 ( .A1(n574), .A2(n388), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n389), .B(KEYINPUT110), .ZN(n405) );
  XOR2_X1 U448 ( .A(n391), .B(n390), .Z(n404) );
  XOR2_X1 U449 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n393) );
  NAND2_X1 U450 ( .A1(G229GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U452 ( .A(n394), .B(KEYINPUT30), .Z(n402) );
  XOR2_X1 U453 ( .A(G141GAT), .B(G36GAT), .Z(n396) );
  XNOR2_X1 U454 ( .A(G50GAT), .B(G29GAT), .ZN(n395) );
  XNOR2_X1 U455 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U456 ( .A(KEYINPUT66), .B(G113GAT), .Z(n398) );
  XNOR2_X1 U457 ( .A(G169GAT), .B(G197GAT), .ZN(n397) );
  XNOR2_X1 U458 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U461 ( .A(n404), .B(n403), .Z(n569) );
  AND2_X1 U462 ( .A1(n405), .A2(n569), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n406), .B(KEYINPUT111), .ZN(n414) );
  XOR2_X1 U464 ( .A(KEYINPUT41), .B(n574), .Z(n538) );
  INV_X1 U465 ( .A(n538), .ZN(n551) );
  NOR2_X1 U466 ( .A1(n569), .A2(n551), .ZN(n408) );
  XNOR2_X1 U467 ( .A(KEYINPUT46), .B(KEYINPUT109), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n408), .B(n407), .ZN(n409) );
  NAND2_X1 U469 ( .A1(n409), .A2(n556), .ZN(n411) );
  INV_X1 U470 ( .A(n410), .ZN(n559) );
  NOR2_X1 U471 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U472 ( .A(KEYINPUT47), .B(n412), .ZN(n413) );
  AND2_X1 U473 ( .A1(n414), .A2(n413), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n416), .B(n415), .ZN(n530) );
  XOR2_X1 U475 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n418) );
  NAND2_X1 U476 ( .A1(G226GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U477 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U478 ( .A(n420), .B(n419), .Z(n423) );
  XNOR2_X1 U479 ( .A(G8GAT), .B(n421), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n427) );
  XOR2_X1 U482 ( .A(n427), .B(n426), .Z(n498) );
  INV_X1 U483 ( .A(n498), .ZN(n520) );
  NOR2_X1 U484 ( .A1(n530), .A2(n520), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n428), .B(KEYINPUT54), .ZN(n450) );
  XOR2_X1 U486 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n430) );
  XNOR2_X1 U487 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U489 ( .A(KEYINPUT6), .B(n431), .Z(n433) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U492 ( .A(n434), .B(KEYINPUT92), .Z(n437) );
  XNOR2_X1 U493 ( .A(G1GAT), .B(n435), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n437), .B(n436), .ZN(n445) );
  XOR2_X1 U495 ( .A(KEYINPUT95), .B(KEYINPUT93), .Z(n439) );
  XNOR2_X1 U496 ( .A(KEYINPUT4), .B(KEYINPUT94), .ZN(n438) );
  XNOR2_X1 U497 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U498 ( .A(n440), .B(G85GAT), .Z(n443) );
  XNOR2_X1 U499 ( .A(G162GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U501 ( .A(n445), .B(n444), .Z(n449) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n449), .B(n448), .ZN(n473) );
  XOR2_X1 U504 ( .A(KEYINPUT96), .B(n473), .Z(n494) );
  INV_X1 U505 ( .A(n494), .ZN(n517) );
  NAND2_X1 U506 ( .A1(n450), .A2(n517), .ZN(n458) );
  NOR2_X1 U507 ( .A1(n451), .A2(n458), .ZN(n452) );
  XNOR2_X1 U508 ( .A(n452), .B(KEYINPUT120), .ZN(n579) );
  INV_X1 U509 ( .A(n579), .ZN(n570) );
  NOR2_X1 U510 ( .A1(n488), .A2(n570), .ZN(n457) );
  XOR2_X1 U511 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n454) );
  XNOR2_X1 U512 ( .A(G218GAT), .B(KEYINPUT125), .ZN(n453) );
  XOR2_X1 U513 ( .A(n454), .B(n453), .Z(n455) );
  NOR2_X1 U514 ( .A1(n458), .A2(n466), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n459), .B(KEYINPUT55), .ZN(n460) );
  NOR2_X2 U516 ( .A1(n522), .A2(n460), .ZN(n566) );
  NAND2_X1 U517 ( .A1(n566), .A2(n538), .ZN(n463) );
  XOR2_X1 U518 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n461) );
  XNOR2_X1 U519 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n481) );
  NOR2_X1 U520 ( .A1(n569), .A2(n574), .ZN(n492) );
  XOR2_X1 U521 ( .A(KEYINPUT28), .B(n466), .Z(n525) );
  INV_X1 U522 ( .A(n525), .ZN(n535) );
  XNOR2_X1 U523 ( .A(KEYINPUT27), .B(n498), .ZN(n469) );
  NAND2_X1 U524 ( .A1(n494), .A2(n469), .ZN(n529) );
  NOR2_X1 U525 ( .A1(n535), .A2(n529), .ZN(n464) );
  NAND2_X1 U526 ( .A1(n522), .A2(n464), .ZN(n475) );
  XNOR2_X1 U527 ( .A(KEYINPUT25), .B(KEYINPUT100), .ZN(n468) );
  NOR2_X1 U528 ( .A1(n522), .A2(n520), .ZN(n465) );
  NOR2_X1 U529 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U530 ( .A(n468), .B(n467), .ZN(n471) );
  NAND2_X1 U531 ( .A1(n548), .A2(n469), .ZN(n470) );
  NAND2_X1 U532 ( .A1(n471), .A2(n470), .ZN(n472) );
  NAND2_X1 U533 ( .A1(n473), .A2(n472), .ZN(n474) );
  NAND2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n489) );
  NOR2_X1 U535 ( .A1(n556), .A2(n410), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n476), .B(KEYINPUT16), .ZN(n477) );
  XOR2_X1 U537 ( .A(KEYINPUT77), .B(n477), .Z(n478) );
  AND2_X1 U538 ( .A1(n489), .A2(n478), .ZN(n506) );
  NAND2_X1 U539 ( .A1(n492), .A2(n506), .ZN(n479) );
  XNOR2_X1 U540 ( .A(KEYINPUT101), .B(n479), .ZN(n486) );
  NAND2_X1 U541 ( .A1(n494), .A2(n486), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(G1324GAT) );
  NAND2_X1 U543 ( .A1(n486), .A2(n498), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n482), .B(KEYINPUT102), .ZN(n483) );
  XNOR2_X1 U545 ( .A(G8GAT), .B(n483), .ZN(G1325GAT) );
  XOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT35), .Z(n485) );
  NAND2_X1 U547 ( .A1(n486), .A2(n531), .ZN(n484) );
  XNOR2_X1 U548 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NAND2_X1 U549 ( .A1(n486), .A2(n535), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n487), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n496) );
  NOR2_X1 U552 ( .A1(n488), .A2(n578), .ZN(n490) );
  NAND2_X1 U553 ( .A1(n490), .A2(n489), .ZN(n491) );
  XNOR2_X1 U554 ( .A(KEYINPUT37), .B(n491), .ZN(n516) );
  NAND2_X1 U555 ( .A1(n492), .A2(n516), .ZN(n493) );
  XOR2_X1 U556 ( .A(KEYINPUT38), .B(n493), .Z(n503) );
  NAND2_X1 U557 ( .A1(n494), .A2(n503), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U559 ( .A(G29GAT), .B(n497), .Z(G1328GAT) );
  NAND2_X1 U560 ( .A1(n498), .A2(n503), .ZN(n499) );
  XNOR2_X1 U561 ( .A(G36GAT), .B(n499), .ZN(G1329GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT104), .B(KEYINPUT40), .Z(n501) );
  NAND2_X1 U563 ( .A1(n503), .A2(n531), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U565 ( .A(G43GAT), .B(n502), .Z(G1330GAT) );
  XOR2_X1 U566 ( .A(G50GAT), .B(KEYINPUT105), .Z(n505) );
  NAND2_X1 U567 ( .A1(n535), .A2(n503), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(G1331GAT) );
  INV_X1 U569 ( .A(n569), .ZN(n562) );
  NOR2_X1 U570 ( .A1(n562), .A2(n551), .ZN(n515) );
  NAND2_X1 U571 ( .A1(n506), .A2(n515), .ZN(n512) );
  NOR2_X1 U572 ( .A1(n517), .A2(n512), .ZN(n507) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n507), .Z(n508) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(n508), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n520), .A2(n512), .ZN(n509) );
  XOR2_X1 U576 ( .A(G64GAT), .B(n509), .Z(G1333GAT) );
  NOR2_X1 U577 ( .A1(n522), .A2(n512), .ZN(n510) );
  XOR2_X1 U578 ( .A(KEYINPUT106), .B(n510), .Z(n511) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(n511), .ZN(G1334GAT) );
  NOR2_X1 U580 ( .A1(n525), .A2(n512), .ZN(n514) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n513) );
  XNOR2_X1 U582 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NAND2_X1 U583 ( .A1(n516), .A2(n515), .ZN(n524) );
  NOR2_X1 U584 ( .A1(n517), .A2(n524), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(G1336GAT) );
  NOR2_X1 U587 ( .A1(n520), .A2(n524), .ZN(n521) );
  XOR2_X1 U588 ( .A(G92GAT), .B(n521), .Z(G1337GAT) );
  NOR2_X1 U589 ( .A1(n522), .A2(n524), .ZN(n523) );
  XOR2_X1 U590 ( .A(G99GAT), .B(n523), .Z(G1338GAT) );
  NOR2_X1 U591 ( .A1(n525), .A2(n524), .ZN(n527) );
  XNOR2_X1 U592 ( .A(KEYINPUT108), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U594 ( .A(G106GAT), .B(n528), .Z(G1339GAT) );
  INV_X1 U595 ( .A(KEYINPUT113), .ZN(n533) );
  NOR2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n549) );
  NAND2_X1 U597 ( .A1(n549), .A2(n531), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n534) );
  NOR2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(KEYINPUT114), .B(n536), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n562), .A2(n545), .ZN(n537) );
  XNOR2_X1 U602 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n540) );
  NAND2_X1 U604 ( .A1(n538), .A2(n545), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(n542) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT115), .Z(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  NAND2_X1 U608 ( .A1(n545), .A2(n578), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n543), .B(KEYINPUT50), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U612 ( .A1(n410), .A2(n545), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n558) );
  NOR2_X1 U615 ( .A1(n569), .A2(n558), .ZN(n550) );
  XOR2_X1 U616 ( .A(G141GAT), .B(n550), .Z(G1344GAT) );
  NOR2_X1 U617 ( .A1(n558), .A2(n551), .ZN(n555) );
  XOR2_X1 U618 ( .A(KEYINPUT117), .B(KEYINPUT52), .Z(n553) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n556), .A2(n558), .ZN(n557) );
  XOR2_X1 U623 ( .A(G155GAT), .B(n557), .Z(G1346GAT) );
  NOR2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT118), .B(n560), .Z(n561) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(n561), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n566), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n563), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U629 ( .A(G183GAT), .B(KEYINPUT119), .Z(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n578), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n410), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(KEYINPUT58), .ZN(n568) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(n568), .ZN(G1351GAT) );
  NOR2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n573) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT59), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT121), .B(KEYINPUT61), .Z(n576) );
  NAND2_X1 U640 ( .A1(n579), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(G204GAT), .B(n577), .Z(G1353GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n581) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n582), .ZN(G1354GAT) );
endmodule

