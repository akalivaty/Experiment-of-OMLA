//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1256, new_n1257, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT64), .Z(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n222), .B1(new_n202), .B2(new_n223), .C1(new_n203), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n207), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n210), .B1(new_n214), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G226), .B(G232), .Z(new_n229));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  XOR2_X1   g0044(.A(KEYINPUT8), .B(G58), .Z(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G13), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n247), .A2(G1), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G20), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n252), .A2(new_n211), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(G1), .B2(new_n212), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n251), .B1(new_n246), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n202), .A2(new_n203), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G58), .A2(G68), .ZN(new_n257));
  OAI21_X1  g0057(.A(G20), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G159), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(KEYINPUT7), .B1(new_n266), .B2(new_n212), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT72), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n203), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT7), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(G20), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT72), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n261), .B1(new_n269), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n253), .B1(new_n275), .B2(KEYINPUT16), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT16), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n270), .A2(G20), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n262), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n265), .ZN(new_n280));
  AOI21_X1  g0080(.A(KEYINPUT73), .B1(new_n262), .B2(KEYINPUT3), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n278), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n203), .B1(new_n282), .B2(new_n272), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n277), .B1(new_n283), .B2(new_n261), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n255), .B1(new_n276), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G169), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G1), .A3(G13), .ZN(new_n288));
  OR2_X1    g0088(.A1(G223), .A2(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G226), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G1698), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n263), .A2(new_n289), .A3(new_n265), .A4(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G87), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n288), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  INV_X1    g0096(.A(G45), .ZN(new_n297));
  AOI21_X1  g0097(.A(G1), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n298), .A2(new_n288), .A3(G274), .ZN(new_n299));
  INV_X1    g0099(.A(G1), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(G41), .B2(G45), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n288), .A2(G232), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n286), .B1(new_n295), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n294), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT18), .B1(new_n285), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n261), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT72), .ZN(new_n311));
  OAI21_X1  g0111(.A(G68), .B1(new_n272), .B2(KEYINPUT72), .ZN(new_n312));
  OAI211_X1 g0112(.A(KEYINPUT16), .B(new_n310), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n252), .A2(new_n211), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(new_n284), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n255), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT18), .ZN(new_n318));
  INV_X1    g0118(.A(new_n308), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT17), .ZN(new_n321));
  INV_X1    g0121(.A(G190), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n295), .A2(new_n322), .A3(new_n304), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n294), .B2(new_n303), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n321), .B1(new_n285), .B2(new_n326), .ZN(new_n327));
  AND4_X1   g0127(.A1(new_n321), .A2(new_n315), .A3(new_n316), .A4(new_n326), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n309), .B(new_n320), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT67), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n262), .B2(G20), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n212), .A2(KEYINPUT67), .A3(G33), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G77), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n259), .A2(G50), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n203), .A2(G20), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n314), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT11), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n338), .A2(KEYINPUT11), .A3(new_n314), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n248), .A2(KEYINPUT12), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n250), .A2(KEYINPUT12), .B1(new_n337), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n254), .A2(KEYINPUT12), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n344), .B1(new_n345), .B2(G68), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n341), .A2(new_n342), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n223), .A2(G1698), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n271), .B(new_n349), .C1(G226), .C2(G1698), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G97), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n288), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n288), .A2(new_n301), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n299), .B1(new_n224), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT13), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT70), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT13), .B1(new_n352), .B2(new_n354), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT14), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n355), .A2(KEYINPUT70), .A3(new_n356), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n360), .A2(new_n361), .A3(G169), .A4(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n357), .A2(KEYINPUT71), .A3(G179), .A4(new_n359), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n357), .A2(G179), .A3(new_n359), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT71), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n363), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n360), .A2(G169), .A3(new_n362), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT14), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n348), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n322), .B1(new_n355), .B2(new_n356), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n347), .B1(new_n359), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n360), .A2(G200), .A3(new_n362), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n334), .A2(new_n245), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n259), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n253), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n250), .A2(new_n201), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n254), .B2(new_n201), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT9), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT9), .B1(new_n379), .B2(new_n381), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n299), .B1(new_n290), .B2(new_n353), .ZN(new_n386));
  NOR2_X1   g0186(.A1(G222), .A2(G1698), .ZN(new_n387));
  INV_X1    g0187(.A(G1698), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(G223), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n271), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n266), .A2(new_n217), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT66), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n288), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n390), .A2(KEYINPUT66), .A3(new_n391), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n386), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n384), .A2(new_n385), .B1(new_n396), .B2(G190), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n396), .A2(new_n324), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT10), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n384), .A2(new_n385), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT69), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n396), .A2(G190), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n399), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n397), .B(new_n398), .C1(new_n402), .C2(KEYINPUT10), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n299), .ZN(new_n409));
  INV_X1    g0209(.A(new_n353), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n409), .B1(G244), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G238), .A2(G1698), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n271), .B(new_n412), .C1(new_n223), .C2(G1698), .ZN(new_n413));
  INV_X1    g0213(.A(new_n288), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n413), .B(new_n414), .C1(G107), .C2(new_n271), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n416), .A2(new_n322), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(G200), .B2(new_n416), .ZN(new_n418));
  XNOR2_X1  g0218(.A(KEYINPUT15), .B(G87), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT68), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n334), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n245), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n253), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n250), .A2(new_n217), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n254), .B2(new_n217), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n382), .B1(new_n396), .B2(new_n306), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G169), .B2(new_n396), .ZN(new_n430));
  INV_X1    g0230(.A(new_n427), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n416), .A2(new_n286), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n411), .A2(new_n415), .A3(new_n306), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n428), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  AND4_X1   g0235(.A1(new_n330), .A2(new_n376), .A3(new_n408), .A4(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT76), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n438), .A2(new_n296), .A3(KEYINPUT5), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT5), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(KEYINPUT76), .B2(G41), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n297), .A2(G1), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n288), .A2(G274), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G270), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n443), .A2(new_n288), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(G257), .A2(G1698), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n388), .A2(G264), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n271), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(G303), .B2(new_n271), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT78), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n288), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n452), .B(KEYINPUT78), .C1(G303), .C2(new_n271), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n449), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G190), .ZN(new_n458));
  INV_X1    g0258(.A(G116), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n250), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n300), .A2(G33), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n253), .A2(new_n249), .A3(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n460), .B1(new_n462), .B2(new_n459), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G283), .ZN(new_n464));
  INV_X1    g0264(.A(G97), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n464), .B(new_n212), .C1(G33), .C2(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n466), .B(new_n314), .C1(new_n212), .C2(G116), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT20), .ZN(new_n468));
  OR2_X1    g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n468), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n458), .B(new_n471), .C1(new_n324), .C2(new_n457), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n453), .A2(new_n454), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(new_n414), .A3(new_n456), .ZN(new_n474));
  INV_X1    g0274(.A(new_n449), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n476), .A2(new_n306), .A3(new_n471), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n286), .B1(new_n474), .B2(new_n475), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT21), .ZN(new_n480));
  INV_X1    g0280(.A(new_n471), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n480), .B1(new_n479), .B2(new_n481), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n472), .B(new_n478), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n271), .A2(G250), .A3(new_n388), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G294), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n263), .A2(new_n265), .A3(G257), .A4(G1698), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n414), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n443), .A2(G264), .A3(new_n288), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n446), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G169), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT80), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n493), .A2(KEYINPUT80), .A3(G169), .ZN(new_n497));
  INV_X1    g0297(.A(new_n448), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n414), .A2(new_n490), .B1(new_n498), .B2(G264), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(G179), .A3(new_n446), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n496), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n249), .A2(G107), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n502), .B(KEYINPUT25), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n462), .A2(KEYINPUT74), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT74), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n253), .A2(new_n249), .A3(new_n505), .A4(new_n461), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(G107), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n271), .A2(new_n212), .A3(G87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT22), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT22), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n271), .A2(new_n511), .A3(new_n212), .A4(G87), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT23), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n212), .B2(G107), .ZN(new_n515));
  INV_X1    g0315(.A(G107), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(KEYINPUT23), .A3(G20), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(KEYINPUT79), .A2(KEYINPUT24), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G116), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(G20), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(KEYINPUT79), .A2(KEYINPUT24), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n253), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n513), .B(new_n522), .C1(KEYINPUT79), .C2(KEYINPUT24), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n508), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n501), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(KEYINPUT81), .B1(new_n493), .B2(G190), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT81), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n499), .A2(new_n531), .A3(new_n322), .A4(new_n446), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n493), .A2(new_n324), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n527), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n220), .B1(new_n297), .B2(G1), .ZN(new_n537));
  INV_X1    g0337(.A(G274), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n300), .A2(new_n538), .A3(G45), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n288), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT77), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT77), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n288), .A2(new_n537), .A3(new_n539), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n218), .A2(G1698), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(G238), .B2(G1698), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n520), .B1(new_n545), .B2(new_n266), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n541), .A2(new_n543), .B1(new_n546), .B2(new_n414), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(G169), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n306), .B2(new_n547), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT19), .B1(new_n334), .B2(G97), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n271), .A2(new_n212), .A3(G68), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT19), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n212), .B1(new_n351), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n219), .A2(new_n465), .A3(new_n516), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n314), .B1(new_n550), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n504), .A2(new_n421), .A3(new_n506), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n419), .B(KEYINPUT68), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n250), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n549), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n504), .A2(G87), .A3(new_n506), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n557), .A2(new_n563), .A3(new_n560), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n541), .A2(new_n543), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n546), .A2(new_n414), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G200), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n565), .B(new_n569), .C1(new_n322), .C2(new_n568), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n562), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT75), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n282), .A2(new_n272), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G107), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n516), .A2(KEYINPUT6), .A3(G97), .ZN(new_n576));
  XOR2_X1   g0376(.A(G97), .B(G107), .Z(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(KEYINPUT6), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n253), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n504), .A2(G97), .A3(new_n506), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n250), .A2(new_n465), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n573), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n575), .A2(new_n579), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n314), .ZN(new_n586));
  INV_X1    g0386(.A(new_n583), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT75), .ZN(new_n588));
  INV_X1    g0388(.A(G257), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n446), .B1(new_n589), .B2(new_n448), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n266), .A2(new_n220), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT4), .ZN(new_n592));
  OAI21_X1  g0392(.A(G1698), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n266), .B2(new_n218), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n271), .A2(KEYINPUT4), .A3(G244), .A4(new_n388), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n593), .A2(new_n464), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n590), .B1(new_n596), .B2(new_n414), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n597), .A2(G200), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n594), .A2(new_n595), .A3(new_n464), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n271), .A2(G250), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n388), .B1(new_n600), .B2(KEYINPUT4), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n414), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n445), .B1(new_n498), .B2(G257), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(G190), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n584), .B(new_n588), .C1(new_n598), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(G169), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n306), .B2(new_n604), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n586), .A2(new_n587), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n486), .A2(new_n536), .A3(new_n572), .A4(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n437), .A2(new_n612), .ZN(G372));
  INV_X1    g0413(.A(KEYINPUT83), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n407), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT83), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n285), .A2(new_n321), .A3(new_n326), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n315), .A2(new_n316), .A3(new_n326), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT17), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n373), .A2(new_n374), .ZN(new_n622));
  INV_X1    g0422(.A(new_n434), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n621), .B1(new_n371), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n318), .B1(new_n317), .B2(new_n319), .ZN(new_n627));
  AOI211_X1 g0427(.A(KEYINPUT18), .B(new_n308), .C1(new_n315), .C2(new_n316), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n617), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n430), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT84), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n615), .A2(new_n616), .ZN(new_n633));
  INV_X1    g0433(.A(new_n629), .ZN(new_n634));
  INV_X1    g0434(.A(new_n370), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n363), .A2(new_n364), .A3(new_n367), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n347), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n637), .A2(new_n624), .B1(new_n620), .B2(new_n618), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n633), .B1(new_n634), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT84), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(new_n640), .A3(new_n430), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n632), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n564), .B1(G190), .B2(new_n547), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n569), .A2(KEYINPUT82), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT82), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n568), .A2(new_n645), .A3(G200), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n534), .A2(new_n527), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n648), .A2(new_n606), .A3(new_n610), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n476), .A2(new_n481), .A3(G169), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT21), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n477), .B1(new_n651), .B2(new_n482), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n529), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n562), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT26), .B1(new_n571), .B2(new_n610), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n643), .A2(new_n647), .B1(new_n549), .B2(new_n561), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n588), .A2(new_n584), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n657), .A2(new_n658), .A3(new_n608), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n436), .B1(new_n655), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n642), .A2(new_n662), .ZN(G369));
  INV_X1    g0463(.A(new_n652), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n248), .A2(new_n212), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(G213), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(new_n471), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n485), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n536), .B1(new_n527), .B2(new_n671), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n529), .B2(new_n671), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n529), .A2(new_n670), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n652), .A2(new_n670), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n536), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT85), .ZN(G399));
  NOR2_X1   g0484(.A1(new_n554), .A2(G116), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n208), .A2(new_n296), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n686), .A3(G1), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n215), .B2(new_n686), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  INV_X1    g0489(.A(G330), .ZN(new_n690));
  AND4_X1   g0490(.A1(G179), .A2(new_n547), .A3(new_n492), .A4(new_n491), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(new_n457), .A3(new_n597), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT86), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(KEYINPUT86), .A3(KEYINPUT30), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT31), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT88), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT87), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n568), .A2(new_n306), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n457), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n701), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n476), .A2(KEYINPUT87), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n604), .A2(new_n493), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n699), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  AOI211_X1 g0508(.A(KEYINPUT88), .B(new_n706), .C1(new_n702), .C2(new_n704), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n697), .B(new_n698), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n670), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n652), .A2(new_n472), .A3(new_n610), .A4(new_n606), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n572), .A2(new_n529), .A3(new_n535), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT31), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n457), .A2(new_n700), .A3(new_n701), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT87), .B1(new_n476), .B2(new_n703), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n707), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n697), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n690), .B1(new_n715), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n671), .B1(new_n655), .B2(new_n661), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n657), .A2(KEYINPUT26), .A3(new_n608), .A4(new_n659), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT89), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n659), .A2(new_n608), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n728), .A2(KEYINPUT89), .A3(new_n657), .A4(KEYINPUT26), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n658), .B1(new_n571), .B2(new_n610), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n562), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n649), .B2(new_n653), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n670), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT29), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n721), .B1(new_n724), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n689), .B1(new_n736), .B2(G1), .ZN(G364));
  NOR2_X1   g0537(.A1(new_n247), .A2(G20), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G45), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n686), .A2(G1), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n674), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n212), .A2(new_n306), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G190), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n747), .A2(new_n322), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n749), .A2(new_n203), .B1(new_n751), .B2(new_n201), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n322), .A2(G179), .A3(G200), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n212), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n465), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  OR3_X1    g0556(.A1(new_n212), .A2(KEYINPUT91), .A3(G190), .ZN(new_n757));
  OAI21_X1  g0557(.A(KEYINPUT91), .B1(new_n212), .B2(G190), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n324), .A2(G179), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G107), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n759), .A2(G20), .A3(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n266), .B1(new_n764), .B2(G87), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n746), .A2(G190), .A3(new_n324), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G190), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n746), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n767), .A2(G58), .B1(new_n770), .B2(G77), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n756), .A2(new_n762), .A3(new_n765), .A4(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G179), .A2(G200), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n757), .A2(new_n758), .A3(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G159), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT32), .ZN(new_n777));
  INV_X1    g0577(.A(G317), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n748), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G294), .ZN(new_n782));
  INV_X1    g0582(.A(G326), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n781), .B1(new_n782), .B2(new_n754), .C1(new_n783), .C2(new_n751), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n761), .A2(G283), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n767), .A2(G322), .B1(new_n770), .B2(G311), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n775), .A2(G329), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n271), .B1(new_n764), .B2(G303), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n785), .A2(new_n786), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n772), .A2(new_n777), .B1(new_n784), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n211), .B1(G20), .B2(new_n286), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n743), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n266), .A2(new_n208), .ZN(new_n793));
  INV_X1    g0593(.A(new_n215), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n793), .B1(new_n297), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n240), .B2(new_n297), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n271), .A2(new_n208), .ZN(new_n797));
  INV_X1    g0597(.A(G355), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n797), .A2(new_n798), .B1(G116), .B2(new_n208), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n799), .A2(KEYINPUT90), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(KEYINPUT90), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n796), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n790), .A2(new_n791), .B1(new_n792), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n740), .B1(new_n745), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n740), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n674), .A2(G330), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(new_n806), .B2(new_n675), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT92), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  INV_X1    g0610(.A(new_n661), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n670), .B1(new_n733), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT96), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n434), .B(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n431), .A2(KEYINPUT97), .A3(new_n670), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT97), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n427), .B2(new_n671), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n815), .A2(new_n817), .B1(new_n427), .B2(new_n418), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n812), .A2(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n814), .A2(new_n818), .B1(new_n623), .B2(new_n670), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n821), .B1(new_n812), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n721), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT98), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n824), .A2(new_n825), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n824), .A2(new_n825), .A3(KEYINPUT98), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n828), .A2(new_n829), .A3(new_n740), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n761), .A2(G68), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n201), .B2(new_n763), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT94), .Z(new_n834));
  AOI21_X1  g0634(.A(new_n266), .B1(new_n775), .B2(G132), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(KEYINPUT95), .B2(new_n835), .C1(new_n202), .C2(new_n754), .ZN(new_n836));
  XOR2_X1   g0636(.A(KEYINPUT93), .B(G143), .Z(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n767), .A2(new_n838), .B1(new_n770), .B2(G159), .ZN(new_n839));
  INV_X1    g0639(.A(G150), .ZN(new_n840));
  INV_X1    g0640(.A(G137), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n839), .B1(new_n749), .B2(new_n840), .C1(new_n841), .C2(new_n751), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT34), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n842), .A2(new_n843), .B1(KEYINPUT95), .B2(new_n835), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n843), .B2(new_n842), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n755), .B1(G283), .B2(new_n748), .ZN(new_n846));
  INV_X1    g0646(.A(G303), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n847), .B2(new_n751), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n516), .A2(new_n763), .B1(new_n769), .B2(new_n459), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n271), .B(new_n849), .C1(G294), .C2(new_n767), .ZN(new_n850));
  INV_X1    g0650(.A(G311), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n219), .B2(new_n760), .C1(new_n851), .C2(new_n774), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n836), .A2(new_n845), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n791), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n791), .A2(new_n741), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n740), .B1(new_n217), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n741), .B2(new_n822), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n831), .A2(new_n859), .ZN(G384));
  AND2_X1   g0660(.A1(new_n578), .A2(KEYINPUT35), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n578), .A2(KEYINPUT35), .ZN(new_n862));
  NOR4_X1   g0662(.A1(new_n861), .A2(new_n862), .A3(new_n459), .A4(new_n214), .ZN(new_n863));
  XNOR2_X1  g0663(.A(KEYINPUT99), .B(KEYINPUT36), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n863), .B(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n794), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n201), .A2(G68), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n300), .B(G13), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n634), .A2(new_n668), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n619), .A2(new_n872), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n315), .A2(new_n316), .B1(new_n308), .B2(new_n668), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT101), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n313), .A2(new_n284), .A3(new_n314), .ZN(new_n876));
  INV_X1    g0676(.A(new_n668), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n876), .A2(new_n255), .B1(new_n319), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT101), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(new_n879), .A3(new_n872), .A4(new_n619), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n275), .A2(KEYINPUT16), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n255), .B1(new_n882), .B2(new_n276), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n619), .B1(new_n883), .B2(new_n668), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n308), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n871), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT100), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n883), .A2(new_n668), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n888), .B(new_n889), .C1(new_n629), .C2(new_n621), .ZN(new_n890));
  INV_X1    g0690(.A(new_n889), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT100), .B1(new_n329), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n887), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT102), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n887), .B(KEYINPUT102), .C1(new_n890), .C2(new_n892), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n881), .A2(new_n886), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n890), .B2(new_n892), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n895), .A2(new_n896), .B1(new_n871), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n814), .A2(new_n670), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n812), .B2(new_n820), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n348), .A2(new_n671), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n637), .A2(new_n622), .A3(new_n904), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n370), .A2(new_n363), .A3(new_n364), .A4(new_n367), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n347), .B(new_n670), .C1(new_n906), .C2(new_n375), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n285), .B(new_n668), .C1(new_n629), .C2(new_n621), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n285), .A2(KEYINPUT104), .A3(new_n326), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT104), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n619), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n912), .A2(new_n914), .A3(new_n878), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n880), .A2(new_n875), .B1(new_n915), .B2(KEYINPUT37), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n910), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT39), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n893), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n898), .A2(new_n871), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n329), .A2(new_n891), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n888), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n329), .A2(KEYINPUT100), .A3(new_n891), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT102), .B1(new_n925), .B2(new_n887), .ZN(new_n926));
  INV_X1    g0726(.A(new_n896), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n921), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n920), .B1(new_n928), .B2(KEYINPUT39), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n371), .A2(new_n671), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n870), .B1(new_n899), .B2(new_n909), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n724), .A2(new_n436), .A3(new_n735), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n642), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n931), .B(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT40), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n822), .B1(new_n905), .B2(new_n907), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n612), .A2(KEYINPUT31), .B1(new_n710), .B2(new_n670), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n670), .A2(KEYINPUT31), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n718), .A2(KEYINPUT88), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n705), .A2(new_n699), .A3(new_n707), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n938), .B1(new_n941), .B2(new_n697), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n936), .B1(new_n937), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n935), .B1(new_n899), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n942), .B1(new_n711), .B2(new_n714), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n893), .A2(new_n917), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n946), .A2(new_n947), .A3(KEYINPUT40), .A4(new_n936), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n437), .A2(new_n945), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n690), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n950), .B2(new_n949), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n934), .A2(new_n952), .B1(new_n300), .B2(new_n738), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT105), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n934), .A2(new_n952), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n953), .B2(new_n954), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n869), .B1(new_n955), .B2(new_n957), .ZN(G367));
  INV_X1    g0758(.A(new_n236), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n792), .B1(new_n559), .B2(new_n208), .C1(new_n959), .C2(new_n793), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n805), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT111), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n565), .A2(new_n671), .ZN(new_n963));
  MUX2_X1   g0763(.A(new_n657), .B(new_n732), .S(new_n963), .Z(new_n964));
  NOR2_X1   g0764(.A1(new_n763), .A2(new_n459), .ZN(new_n965));
  AOI22_X1  g0765(.A1(KEYINPUT46), .A2(new_n965), .B1(new_n748), .B2(G294), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n516), .B2(new_n754), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n465), .A2(new_n760), .B1(new_n774), .B2(new_n778), .ZN(new_n968));
  INV_X1    g0768(.A(G283), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n266), .B1(new_n769), .B2(new_n969), .C1(new_n847), .C2(new_n766), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n751), .A2(new_n851), .B1(KEYINPUT46), .B2(new_n965), .ZN(new_n971));
  NOR4_X1   g0771(.A1(new_n967), .A2(new_n968), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT112), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n202), .A2(new_n763), .B1(new_n769), .B2(new_n201), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n266), .B(new_n974), .C1(G150), .C2(new_n767), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n761), .A2(G77), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n975), .B(new_n976), .C1(new_n841), .C2(new_n774), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n754), .A2(new_n203), .ZN(new_n978));
  INV_X1    g0778(.A(G159), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n751), .A2(new_n837), .B1(new_n749), .B2(new_n979), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n973), .A2(new_n981), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n982), .A2(KEYINPUT47), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n791), .B1(new_n982), .B2(KEYINPUT47), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n962), .B1(new_n744), .B2(new_n964), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n659), .A2(new_n670), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n611), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n728), .A2(new_n670), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT106), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT106), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n529), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT107), .ZN(new_n997));
  INV_X1    g0797(.A(new_n610), .ZN(new_n998));
  OR3_X1    g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n997), .B1(new_n996), .B2(new_n998), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n999), .A2(new_n1000), .A3(new_n671), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n681), .A2(new_n536), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n992), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT42), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n986), .B(new_n987), .C1(new_n1001), .C2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1001), .A2(new_n1004), .A3(new_n987), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT108), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1005), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n679), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n993), .A2(new_n995), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n739), .A2(G1), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n1016));
  XNOR2_X1  g0816(.A(new_n686), .B(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n682), .A2(new_n991), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT44), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n682), .A2(new_n991), .ZN(new_n1021));
  XOR2_X1   g0821(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n1022));
  XNOR2_X1  g0822(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n1011), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1020), .A2(new_n679), .A3(new_n1023), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1002), .B1(new_n678), .B2(new_n681), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(new_n676), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n736), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1018), .B1(new_n1031), .B2(new_n736), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n1010), .A2(new_n1014), .B1(new_n1015), .B2(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n985), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(KEYINPUT113), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT113), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1037), .B(new_n985), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(G387));
  OR2_X1    g0840(.A1(new_n678), .A2(new_n744), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n797), .A2(new_n685), .B1(G107), .B2(new_n208), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n233), .A2(G45), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n245), .A2(new_n201), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT50), .Z(new_n1045));
  INV_X1    g0845(.A(new_n685), .ZN(new_n1046));
  AOI211_X1 g0846(.A(G45), .B(new_n1046), .C1(G68), .C2(G77), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n793), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1042), .B1(new_n1043), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n792), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n805), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n766), .A2(new_n201), .B1(new_n769), .B2(new_n203), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n266), .B(new_n1052), .C1(G77), .C2(new_n764), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G159), .A2(new_n750), .B1(new_n748), .B2(new_n245), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n754), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n421), .A2(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G97), .A2(new_n761), .B1(new_n775), .B2(G150), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1053), .A2(new_n1054), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n767), .A2(G317), .B1(new_n770), .B2(G303), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n750), .A2(G322), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(new_n851), .C2(new_n749), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1055), .A2(G283), .B1(new_n764), .B2(G294), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT114), .Z(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(KEYINPUT49), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n266), .B1(new_n760), .B2(new_n459), .C1(new_n783), .C2(new_n774), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT115), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1067), .A2(KEYINPUT49), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1058), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1051), .B1(new_n1073), .B2(new_n791), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1029), .A2(new_n1015), .B1(new_n1041), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n686), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1030), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1029), .A2(new_n736), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(G393));
  NAND2_X1  g0879(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1031), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1015), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1027), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n993), .A2(new_n743), .A3(new_n995), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n792), .B1(new_n465), .B2(new_n208), .C1(new_n243), .C2(new_n793), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n805), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n266), .B1(new_n769), .B2(new_n782), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n749), .A2(new_n847), .B1(new_n459), .B2(new_n754), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(G283), .C2(new_n764), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n751), .A2(new_n778), .B1(new_n851), .B2(new_n766), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT52), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n775), .A2(G322), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1089), .A2(new_n762), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n751), .A2(new_n840), .B1(new_n979), .B2(new_n766), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT51), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n271), .B1(new_n763), .B2(new_n203), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n761), .B2(G87), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1095), .B(new_n1097), .C1(new_n774), .C2(new_n837), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n754), .A2(new_n217), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n246), .B2(new_n769), .C1(new_n201), .C2(new_n749), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT116), .Z(new_n1102));
  OAI21_X1  g0902(.A(new_n1093), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1086), .B1(new_n1103), .B2(new_n791), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1083), .B1(new_n1084), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1081), .A2(new_n1105), .ZN(G390));
  AOI21_X1  g0906(.A(new_n908), .B1(new_n721), .B2(new_n823), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n908), .A2(new_n823), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n945), .A2(new_n1108), .A3(new_n690), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n902), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n715), .A2(new_n720), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1111), .A2(new_n908), .A3(G330), .A4(new_n823), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n900), .B1(new_n734), .B2(new_n820), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n945), .A2(new_n690), .A3(new_n822), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1112), .B(new_n1113), .C1(new_n1114), .C2(new_n908), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n946), .A2(G330), .A3(new_n436), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n642), .A2(new_n932), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n908), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n930), .B1(new_n901), .B2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1122), .B(new_n919), .C1(new_n899), .C2(new_n918), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n930), .B(new_n947), .C1(new_n1113), .C2(new_n1121), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n1112), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1109), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1120), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1118), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1123), .A2(new_n1124), .A3(new_n1112), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1124), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n929), .B2(new_n1122), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1129), .B(new_n1130), .C1(new_n1132), .C2(new_n1126), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1128), .A2(new_n1133), .A3(new_n1076), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT117), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1128), .A2(new_n1133), .A3(KEYINPUT117), .A4(new_n1076), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n767), .A2(G116), .B1(new_n770), .B2(G97), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n271), .B1(new_n764), .B2(G87), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n832), .A3(new_n1139), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1100), .B1(new_n749), .B2(new_n516), .C1(new_n969), .C2(new_n751), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1140), .B(new_n1141), .C1(G294), .C2(new_n775), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1143), .A2(KEYINPUT118), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n764), .A2(G150), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT53), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(G159), .B2(new_n1055), .ZN(new_n1147));
  INV_X1    g0947(.A(G132), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n271), .B1(new_n766), .B2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT54), .B(G143), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1149), .B1(new_n770), .B2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G128), .A2(new_n750), .B1(new_n748), .B2(G137), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G50), .A2(new_n761), .B1(new_n775), .B2(G125), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1147), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT118), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1155), .B1(new_n1142), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n791), .B1(new_n1144), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n855), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1158), .B(new_n805), .C1(new_n245), .C2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n929), .B2(new_n741), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1161), .B1(new_n1162), .B2(new_n1015), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1136), .A2(new_n1137), .A3(new_n1163), .ZN(G378));
  INV_X1    g0964(.A(new_n791), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n262), .B(new_n296), .C1(new_n760), .C2(new_n979), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G128), .A2(new_n767), .B1(new_n764), .B2(new_n1151), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n841), .B2(new_n769), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G150), .A2(new_n1055), .B1(new_n750), .B2(G125), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1169), .B(new_n1170), .C1(new_n1148), .C2(new_n749), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1166), .B(new_n1172), .C1(G124), .C2(new_n775), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(KEYINPUT59), .B2(new_n1171), .ZN(new_n1174));
  AOI211_X1 g0974(.A(G41), .B(new_n271), .C1(new_n764), .C2(G77), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n516), .B2(new_n766), .C1(new_n969), .C2(new_n774), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n978), .B1(G116), .B2(new_n750), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n465), .B2(new_n749), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n559), .A2(new_n769), .B1(new_n202), .B2(new_n760), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT58), .Z(new_n1181));
  AOI21_X1  g0981(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1174), .B(new_n1181), .C1(G50), .C2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1165), .B1(new_n1183), .B2(KEYINPUT119), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(KEYINPUT119), .B2(new_n1183), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n740), .B1(new_n201), .B2(new_n855), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1187));
  OR3_X1    g0987(.A1(new_n617), .A2(new_n631), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n617), .B2(new_n631), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n382), .B2(new_n668), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n382), .A2(new_n668), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1188), .A2(new_n1192), .A3(new_n1189), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1185), .B(new_n1186), .C1(new_n1194), .C2(new_n742), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n895), .A2(new_n896), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n943), .B1(new_n1197), .B2(new_n921), .ZN(new_n1198));
  OAI211_X1 g0998(.A(G330), .B(new_n948), .C1(new_n1198), .C2(KEYINPUT40), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1194), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1194), .A2(new_n944), .A3(G330), .A4(new_n948), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n931), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n870), .B1(new_n909), .B2(new_n899), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n930), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n919), .B1(new_n899), .B2(new_n918), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1208), .A2(new_n1202), .A3(new_n1201), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1204), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1196), .B1(new_n1210), .B2(new_n1015), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1204), .A2(new_n1209), .B1(new_n1119), .B2(new_n1133), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1076), .B1(new_n1212), .B2(KEYINPUT57), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1133), .A2(new_n1119), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1210), .A2(KEYINPUT57), .A3(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1211), .B1(new_n1213), .B2(new_n1215), .ZN(G375));
  NAND2_X1  g1016(.A1(new_n1116), .A2(new_n1015), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1121), .A2(new_n741), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n805), .B1(G68), .B2(new_n1159), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n774), .A2(new_n847), .B1(new_n763), .B2(new_n465), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT120), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G116), .A2(new_n748), .B1(new_n750), .B2(G294), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n271), .B1(new_n770), .B2(G107), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(new_n969), .C2(new_n766), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1056), .A2(new_n976), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1221), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT121), .Z(new_n1227));
  AOI22_X1  g1027(.A1(G132), .A2(new_n750), .B1(new_n767), .B2(G137), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n749), .B2(new_n1150), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(KEYINPUT122), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(KEYINPUT122), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n271), .B1(new_n769), .B2(new_n840), .C1(new_n979), .C2(new_n763), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G50), .B2(new_n1055), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G58), .A2(new_n761), .B1(new_n775), .B2(G128), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1231), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1227), .B1(new_n1230), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT123), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1165), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1219), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1218), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1217), .A2(KEYINPUT124), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT124), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1082), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1241), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1243), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1129), .A2(new_n1018), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1110), .A2(new_n1118), .A3(new_n1115), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1242), .A2(new_n1246), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(G381));
  AOI21_X1  g1050(.A(G390), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1134), .A2(new_n1163), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1251), .A2(new_n1249), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1254), .A2(G375), .ZN(G407));
  NAND2_X1  g1055(.A1(new_n669), .A2(G213), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1252), .A2(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G407), .B(G213), .C1(G375), .C2(new_n1258), .ZN(G409));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT126), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1081), .A2(new_n1105), .A3(new_n1261), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n985), .B(new_n1262), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G390), .A2(KEYINPUT126), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1264), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n985), .B(new_n1266), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(G393), .B(new_n809), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1265), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1035), .A2(G390), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1268), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1260), .B(new_n1269), .C1(new_n1251), .C2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1242), .A2(new_n1246), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT60), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1248), .A2(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1110), .A2(new_n1118), .A3(new_n1115), .A4(KEYINPUT60), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1277), .A2(new_n1120), .A3(new_n1076), .A4(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1275), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1275), .A2(G384), .A3(new_n1279), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(G2897), .A3(new_n1257), .A4(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1257), .A2(G2897), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1282), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1284), .B1(new_n1285), .B2(new_n1280), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  XOR2_X1   g1087(.A(new_n1287), .B(KEYINPUT125), .Z(new_n1288));
  OAI211_X1 g1088(.A(G378), .B(new_n1211), .C1(new_n1213), .C2(new_n1215), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1212), .A2(new_n1017), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1209), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1208), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1015), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1195), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1252), .B1(new_n1290), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1289), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1256), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1288), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1257), .B1(new_n1289), .B2(new_n1295), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1285), .A2(new_n1280), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1299), .A2(KEYINPUT63), .A3(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1296), .A2(new_n1256), .A3(new_n1300), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1274), .A2(new_n1298), .A3(new_n1301), .A4(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1269), .B1(new_n1251), .B2(new_n1272), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1287), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1260), .B1(new_n1299), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1302), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1299), .A2(KEYINPUT62), .A3(new_n1300), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1308), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1306), .B1(new_n1312), .B2(KEYINPUT127), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT61), .B1(new_n1297), .B2(new_n1287), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1311), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT62), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1316));
  OAI211_X1 g1116(.A(KEYINPUT127), .B(new_n1314), .C1(new_n1315), .C2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1305), .B1(new_n1313), .B2(new_n1318), .ZN(G405));
  NAND2_X1  g1119(.A1(G375), .A2(new_n1252), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1289), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1321), .B(new_n1300), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1322), .B(new_n1306), .ZN(G402));
endmodule


