

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(G2105), .A2(n519), .ZN(n883) );
  XNOR2_X1 U549 ( .A(n540), .B(KEYINPUT23), .ZN(n541) );
  XOR2_X1 U550 ( .A(n523), .B(KEYINPUT80), .Z(n516) );
  AND2_X1 U551 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X2 U552 ( .A1(n701), .A2(n700), .ZN(n731) );
  INV_X1 U553 ( .A(n731), .ZN(n747) );
  NOR2_X1 U554 ( .A1(G1384), .A2(G164), .ZN(n699) );
  INV_X1 U555 ( .A(KEYINPUT66), .ZN(n540) );
  NOR2_X1 U556 ( .A1(G651), .A2(G543), .ZN(n635) );
  NOR2_X1 U557 ( .A1(G651), .A2(n627), .ZN(n641) );
  XNOR2_X1 U558 ( .A(n542), .B(n541), .ZN(n544) );
  NOR2_X1 U559 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U560 ( .A1(n548), .A2(n547), .ZN(G160) );
  NOR2_X1 U561 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  XOR2_X2 U562 ( .A(KEYINPUT17), .B(n517), .Z(n882) );
  NAND2_X1 U563 ( .A1(G138), .A2(n882), .ZN(n518) );
  XNOR2_X1 U564 ( .A(n518), .B(KEYINPUT81), .ZN(n526) );
  INV_X1 U565 ( .A(G2104), .ZN(n519) );
  NAND2_X1 U566 ( .A1(G102), .A2(n883), .ZN(n522) );
  NAND2_X1 U567 ( .A1(n519), .A2(G2105), .ZN(n520) );
  XNOR2_X2 U568 ( .A(n520), .B(KEYINPUT65), .ZN(n879) );
  NAND2_X1 U569 ( .A1(G126), .A2(n879), .ZN(n521) );
  NAND2_X1 U570 ( .A1(n522), .A2(n521), .ZN(n524) );
  AND2_X2 U571 ( .A1(G2105), .A2(G2104), .ZN(n878) );
  NAND2_X1 U572 ( .A1(n878), .A2(G114), .ZN(n523) );
  OR2_X1 U573 ( .A1(n524), .A2(n516), .ZN(n525) );
  XNOR2_X1 U574 ( .A(KEYINPUT82), .B(n527), .ZN(G164) );
  NAND2_X1 U575 ( .A1(n635), .A2(G89), .ZN(n528) );
  XNOR2_X1 U576 ( .A(n528), .B(KEYINPUT4), .ZN(n530) );
  XOR2_X1 U577 ( .A(KEYINPUT0), .B(G543), .Z(n627) );
  INV_X1 U578 ( .A(G651), .ZN(n532) );
  NOR2_X1 U579 ( .A1(n627), .A2(n532), .ZN(n630) );
  NAND2_X1 U580 ( .A1(G76), .A2(n630), .ZN(n529) );
  NAND2_X1 U581 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U582 ( .A(n531), .B(KEYINPUT5), .ZN(n538) );
  NOR2_X1 U583 ( .A1(G543), .A2(n532), .ZN(n533) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n533), .Z(n633) );
  NAND2_X1 U585 ( .A1(G63), .A2(n633), .ZN(n535) );
  NAND2_X1 U586 ( .A1(G51), .A2(n641), .ZN(n534) );
  NAND2_X1 U587 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U588 ( .A(KEYINPUT6), .B(n536), .Z(n537) );
  NAND2_X1 U589 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U590 ( .A(n539), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U591 ( .A1(G101), .A2(n883), .ZN(n542) );
  NAND2_X1 U592 ( .A1(G113), .A2(n878), .ZN(n543) );
  NAND2_X1 U593 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U594 ( .A1(G137), .A2(n882), .ZN(n546) );
  NAND2_X1 U595 ( .A1(G125), .A2(n879), .ZN(n545) );
  NAND2_X1 U596 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U597 ( .A1(G65), .A2(n633), .ZN(n550) );
  NAND2_X1 U598 ( .A1(G91), .A2(n635), .ZN(n549) );
  NAND2_X1 U599 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U600 ( .A1(G78), .A2(n630), .ZN(n552) );
  NAND2_X1 U601 ( .A1(G53), .A2(n641), .ZN(n551) );
  NAND2_X1 U602 ( .A1(n552), .A2(n551), .ZN(n553) );
  OR2_X1 U603 ( .A1(n554), .A2(n553), .ZN(G299) );
  NAND2_X1 U604 ( .A1(G85), .A2(n635), .ZN(n556) );
  NAND2_X1 U605 ( .A1(G72), .A2(n630), .ZN(n555) );
  NAND2_X1 U606 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U607 ( .A1(G60), .A2(n633), .ZN(n558) );
  NAND2_X1 U608 ( .A1(G47), .A2(n641), .ZN(n557) );
  NAND2_X1 U609 ( .A1(n558), .A2(n557), .ZN(n559) );
  OR2_X1 U610 ( .A1(n560), .A2(n559), .ZN(G290) );
  NAND2_X1 U611 ( .A1(G64), .A2(n633), .ZN(n562) );
  NAND2_X1 U612 ( .A1(G52), .A2(n641), .ZN(n561) );
  NAND2_X1 U613 ( .A1(n562), .A2(n561), .ZN(n567) );
  NAND2_X1 U614 ( .A1(G90), .A2(n635), .ZN(n564) );
  NAND2_X1 U615 ( .A1(G77), .A2(n630), .ZN(n563) );
  NAND2_X1 U616 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U617 ( .A(KEYINPUT9), .B(n565), .Z(n566) );
  NOR2_X1 U618 ( .A1(n567), .A2(n566), .ZN(G171) );
  INV_X1 U619 ( .A(G171), .ZN(G301) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U621 ( .A(G57), .ZN(G237) );
  INV_X1 U622 ( .A(G120), .ZN(G236) );
  NAND2_X1 U623 ( .A1(G7), .A2(G661), .ZN(n568) );
  XOR2_X1 U624 ( .A(n568), .B(KEYINPUT10), .Z(n906) );
  NAND2_X1 U625 ( .A1(n906), .A2(G567), .ZN(n569) );
  XOR2_X1 U626 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  NAND2_X1 U627 ( .A1(G56), .A2(n633), .ZN(n570) );
  XOR2_X1 U628 ( .A(KEYINPUT14), .B(n570), .Z(n577) );
  NAND2_X1 U629 ( .A1(G81), .A2(n635), .ZN(n571) );
  XOR2_X1 U630 ( .A(KEYINPUT67), .B(n571), .Z(n572) );
  XNOR2_X1 U631 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U632 ( .A1(G68), .A2(n630), .ZN(n573) );
  NAND2_X1 U633 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U634 ( .A(KEYINPUT13), .B(n575), .Z(n576) );
  NOR2_X1 U635 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U636 ( .A1(n641), .A2(G43), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n579), .A2(n578), .ZN(n911) );
  INV_X1 U638 ( .A(G860), .ZN(n592) );
  OR2_X1 U639 ( .A1(n911), .A2(n592), .ZN(G153) );
  NAND2_X1 U640 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U641 ( .A1(G66), .A2(n633), .ZN(n581) );
  NAND2_X1 U642 ( .A1(G92), .A2(n635), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U644 ( .A1(G79), .A2(n630), .ZN(n583) );
  NAND2_X1 U645 ( .A1(G54), .A2(n641), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U647 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U648 ( .A(KEYINPUT15), .B(n586), .Z(n907) );
  OR2_X1 U649 ( .A1(n907), .A2(G868), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n588), .A2(n587), .ZN(G284) );
  XOR2_X1 U651 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U652 ( .A(G868), .ZN(n654) );
  NOR2_X1 U653 ( .A1(G286), .A2(n654), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(KEYINPUT68), .ZN(n591) );
  NOR2_X1 U655 ( .A1(G299), .A2(G868), .ZN(n590) );
  NOR2_X1 U656 ( .A1(n591), .A2(n590), .ZN(G297) );
  NAND2_X1 U657 ( .A1(n592), .A2(G559), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n593), .A2(n907), .ZN(n594) );
  XNOR2_X1 U659 ( .A(n594), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U660 ( .A1(G868), .A2(n911), .ZN(n595) );
  XOR2_X1 U661 ( .A(KEYINPUT69), .B(n595), .Z(n599) );
  NAND2_X1 U662 ( .A1(n907), .A2(G868), .ZN(n596) );
  NOR2_X1 U663 ( .A1(G559), .A2(n596), .ZN(n597) );
  XNOR2_X1 U664 ( .A(KEYINPUT70), .B(n597), .ZN(n598) );
  NOR2_X1 U665 ( .A1(n599), .A2(n598), .ZN(G282) );
  NAND2_X1 U666 ( .A1(G111), .A2(n878), .ZN(n601) );
  NAND2_X1 U667 ( .A1(G99), .A2(n883), .ZN(n600) );
  NAND2_X1 U668 ( .A1(n601), .A2(n600), .ZN(n607) );
  NAND2_X1 U669 ( .A1(G123), .A2(n879), .ZN(n602) );
  XOR2_X1 U670 ( .A(KEYINPUT18), .B(n602), .Z(n603) );
  XNOR2_X1 U671 ( .A(n603), .B(KEYINPUT71), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G135), .A2(n882), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U674 ( .A1(n607), .A2(n606), .ZN(n984) );
  XNOR2_X1 U675 ( .A(G2096), .B(n984), .ZN(n608) );
  INV_X1 U676 ( .A(G2100), .ZN(n833) );
  NAND2_X1 U677 ( .A1(n608), .A2(n833), .ZN(G156) );
  NAND2_X1 U678 ( .A1(n907), .A2(G559), .ZN(n651) );
  XNOR2_X1 U679 ( .A(n911), .B(n651), .ZN(n609) );
  NOR2_X1 U680 ( .A1(n609), .A2(G860), .ZN(n616) );
  NAND2_X1 U681 ( .A1(G67), .A2(n633), .ZN(n611) );
  NAND2_X1 U682 ( .A1(G93), .A2(n635), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U684 ( .A1(G80), .A2(n630), .ZN(n613) );
  NAND2_X1 U685 ( .A1(G55), .A2(n641), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n653) );
  XNOR2_X1 U688 ( .A(n616), .B(n653), .ZN(G145) );
  NAND2_X1 U689 ( .A1(G62), .A2(n633), .ZN(n618) );
  NAND2_X1 U690 ( .A1(G88), .A2(n635), .ZN(n617) );
  NAND2_X1 U691 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U692 ( .A1(G75), .A2(n630), .ZN(n620) );
  NAND2_X1 U693 ( .A1(G50), .A2(n641), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U696 ( .A(KEYINPUT75), .B(n623), .ZN(G303) );
  NAND2_X1 U697 ( .A1(G49), .A2(n641), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n633), .A2(n626), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n627), .A2(G87), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n629), .A2(n628), .ZN(G288) );
  XOR2_X1 U703 ( .A(KEYINPUT2), .B(KEYINPUT74), .Z(n632) );
  NAND2_X1 U704 ( .A1(G73), .A2(n630), .ZN(n631) );
  XNOR2_X1 U705 ( .A(n632), .B(n631), .ZN(n640) );
  NAND2_X1 U706 ( .A1(n633), .A2(G61), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n634), .B(KEYINPUT72), .ZN(n637) );
  NAND2_X1 U708 ( .A1(G86), .A2(n635), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U710 ( .A(KEYINPUT73), .B(n638), .Z(n639) );
  NOR2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U712 ( .A1(n641), .A2(G48), .ZN(n642) );
  NAND2_X1 U713 ( .A1(n643), .A2(n642), .ZN(G305) );
  XOR2_X1 U714 ( .A(G303), .B(n653), .Z(n648) );
  XOR2_X1 U715 ( .A(KEYINPUT19), .B(KEYINPUT76), .Z(n644) );
  XNOR2_X1 U716 ( .A(G299), .B(n644), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n645), .B(G290), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n646), .B(G288), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n649), .B(G305), .ZN(n650) );
  XNOR2_X1 U721 ( .A(n650), .B(n911), .ZN(n895) );
  XNOR2_X1 U722 ( .A(n895), .B(n651), .ZN(n652) );
  NOR2_X1 U723 ( .A1(n654), .A2(n652), .ZN(n656) );
  AND2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U725 ( .A1(n656), .A2(n655), .ZN(G295) );
  NAND2_X1 U726 ( .A1(G2084), .A2(G2078), .ZN(n657) );
  XOR2_X1 U727 ( .A(KEYINPUT20), .B(n657), .Z(n658) );
  NAND2_X1 U728 ( .A1(G2090), .A2(n658), .ZN(n659) );
  XNOR2_X1 U729 ( .A(KEYINPUT21), .B(n659), .ZN(n660) );
  NAND2_X1 U730 ( .A1(n660), .A2(G2072), .ZN(n661) );
  XOR2_X1 U731 ( .A(KEYINPUT77), .B(n661), .Z(G158) );
  XNOR2_X1 U732 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U733 ( .A1(G236), .A2(G237), .ZN(n662) );
  NAND2_X1 U734 ( .A1(G69), .A2(n662), .ZN(n663) );
  XNOR2_X1 U735 ( .A(KEYINPUT79), .B(n663), .ZN(n664) );
  NAND2_X1 U736 ( .A1(n664), .A2(G108), .ZN(n826) );
  NAND2_X1 U737 ( .A1(n826), .A2(G567), .ZN(n670) );
  NAND2_X1 U738 ( .A1(G132), .A2(G82), .ZN(n665) );
  XNOR2_X1 U739 ( .A(n665), .B(KEYINPUT22), .ZN(n666) );
  XNOR2_X1 U740 ( .A(n666), .B(KEYINPUT78), .ZN(n667) );
  NOR2_X1 U741 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U742 ( .A1(G96), .A2(n668), .ZN(n827) );
  NAND2_X1 U743 ( .A1(n827), .A2(G2106), .ZN(n669) );
  NAND2_X1 U744 ( .A1(n670), .A2(n669), .ZN(n828) );
  NAND2_X1 U745 ( .A1(G661), .A2(G483), .ZN(n671) );
  NOR2_X1 U746 ( .A1(n828), .A2(n671), .ZN(n824) );
  NAND2_X1 U747 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U748 ( .A1(G160), .A2(G40), .ZN(n700) );
  NOR2_X1 U749 ( .A1(n699), .A2(n700), .ZN(n672) );
  XOR2_X1 U750 ( .A(KEYINPUT83), .B(n672), .Z(n804) );
  NAND2_X1 U751 ( .A1(n882), .A2(G140), .ZN(n673) );
  XNOR2_X1 U752 ( .A(n673), .B(KEYINPUT84), .ZN(n675) );
  NAND2_X1 U753 ( .A1(G104), .A2(n883), .ZN(n674) );
  NAND2_X1 U754 ( .A1(n675), .A2(n674), .ZN(n677) );
  XOR2_X1 U755 ( .A(KEYINPUT34), .B(KEYINPUT85), .Z(n676) );
  XNOR2_X1 U756 ( .A(n677), .B(n676), .ZN(n682) );
  NAND2_X1 U757 ( .A1(G116), .A2(n878), .ZN(n679) );
  NAND2_X1 U758 ( .A1(G128), .A2(n879), .ZN(n678) );
  NAND2_X1 U759 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U760 ( .A(KEYINPUT35), .B(n680), .Z(n681) );
  NOR2_X1 U761 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U762 ( .A(KEYINPUT36), .B(n683), .ZN(n876) );
  XNOR2_X1 U763 ( .A(KEYINPUT37), .B(G2067), .ZN(n802) );
  NOR2_X1 U764 ( .A1(n876), .A2(n802), .ZN(n1004) );
  NAND2_X1 U765 ( .A1(n804), .A2(n1004), .ZN(n800) );
  XOR2_X1 U766 ( .A(KEYINPUT38), .B(KEYINPUT86), .Z(n685) );
  NAND2_X1 U767 ( .A1(G105), .A2(n883), .ZN(n684) );
  XNOR2_X1 U768 ( .A(n685), .B(n684), .ZN(n689) );
  NAND2_X1 U769 ( .A1(G117), .A2(n878), .ZN(n687) );
  NAND2_X1 U770 ( .A1(G129), .A2(n879), .ZN(n686) );
  NAND2_X1 U771 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U772 ( .A1(n689), .A2(n688), .ZN(n691) );
  NAND2_X1 U773 ( .A1(n882), .A2(G141), .ZN(n690) );
  NAND2_X1 U774 ( .A1(n691), .A2(n690), .ZN(n873) );
  AND2_X1 U775 ( .A1(n873), .A2(G1996), .ZN(n985) );
  NAND2_X1 U776 ( .A1(G107), .A2(n878), .ZN(n693) );
  NAND2_X1 U777 ( .A1(G95), .A2(n883), .ZN(n692) );
  NAND2_X1 U778 ( .A1(n693), .A2(n692), .ZN(n697) );
  NAND2_X1 U779 ( .A1(G131), .A2(n882), .ZN(n695) );
  NAND2_X1 U780 ( .A1(G119), .A2(n879), .ZN(n694) );
  NAND2_X1 U781 ( .A1(n695), .A2(n694), .ZN(n696) );
  OR2_X1 U782 ( .A1(n697), .A2(n696), .ZN(n889) );
  AND2_X1 U783 ( .A1(n889), .A2(G1991), .ZN(n987) );
  OR2_X1 U784 ( .A1(n985), .A2(n987), .ZN(n698) );
  NAND2_X1 U785 ( .A1(n804), .A2(n698), .ZN(n793) );
  NAND2_X1 U786 ( .A1(n800), .A2(n793), .ZN(n790) );
  INV_X1 U787 ( .A(n699), .ZN(n701) );
  NAND2_X1 U788 ( .A1(G8), .A2(n747), .ZN(n782) );
  NOR2_X1 U789 ( .A1(G1981), .A2(G305), .ZN(n702) );
  XOR2_X1 U790 ( .A(n702), .B(KEYINPUT24), .Z(n703) );
  NOR2_X1 U791 ( .A1(n782), .A2(n703), .ZN(n704) );
  XNOR2_X1 U792 ( .A(n704), .B(KEYINPUT87), .ZN(n767) );
  AND2_X1 U793 ( .A1(n731), .A2(G1996), .ZN(n705) );
  XNOR2_X1 U794 ( .A(n705), .B(KEYINPUT26), .ZN(n709) );
  NAND2_X1 U795 ( .A1(n747), .A2(G1341), .ZN(n707) );
  INV_X1 U796 ( .A(n911), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n711) );
  NOR2_X1 U799 ( .A1(n711), .A2(n907), .ZN(n710) );
  XNOR2_X1 U800 ( .A(n710), .B(KEYINPUT89), .ZN(n718) );
  NAND2_X1 U801 ( .A1(n711), .A2(n907), .ZN(n716) );
  NAND2_X1 U802 ( .A1(G1348), .A2(n747), .ZN(n713) );
  NAND2_X1 U803 ( .A1(G2067), .A2(n731), .ZN(n712) );
  NAND2_X1 U804 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U805 ( .A(KEYINPUT88), .B(n714), .ZN(n715) );
  NAND2_X1 U806 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U807 ( .A1(n718), .A2(n717), .ZN(n724) );
  NAND2_X1 U808 ( .A1(n731), .A2(G2072), .ZN(n719) );
  XOR2_X1 U809 ( .A(KEYINPUT27), .B(n719), .Z(n721) );
  NAND2_X1 U810 ( .A1(G1956), .A2(n747), .ZN(n720) );
  NAND2_X1 U811 ( .A1(n721), .A2(n720), .ZN(n725) );
  NOR2_X1 U812 ( .A1(G299), .A2(n725), .ZN(n722) );
  XOR2_X1 U813 ( .A(KEYINPUT90), .B(n722), .Z(n723) );
  NAND2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n728) );
  NAND2_X1 U815 ( .A1(G299), .A2(n725), .ZN(n726) );
  XNOR2_X1 U816 ( .A(n726), .B(KEYINPUT28), .ZN(n727) );
  NAND2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n730) );
  XNOR2_X1 U818 ( .A(KEYINPUT91), .B(KEYINPUT29), .ZN(n729) );
  XNOR2_X1 U819 ( .A(n730), .B(n729), .ZN(n735) );
  INV_X1 U820 ( .A(G1961), .ZN(n950) );
  NAND2_X1 U821 ( .A1(n747), .A2(n950), .ZN(n733) );
  XNOR2_X1 U822 ( .A(G2078), .B(KEYINPUT25), .ZN(n965) );
  NAND2_X1 U823 ( .A1(n731), .A2(n965), .ZN(n732) );
  NAND2_X1 U824 ( .A1(n733), .A2(n732), .ZN(n740) );
  NAND2_X1 U825 ( .A1(n740), .A2(G171), .ZN(n734) );
  NAND2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n746) );
  NOR2_X1 U827 ( .A1(G1966), .A2(n782), .ZN(n736) );
  NOR2_X1 U828 ( .A1(G2084), .A2(n747), .ZN(n759) );
  NOR2_X1 U829 ( .A1(n736), .A2(n759), .ZN(n737) );
  NAND2_X1 U830 ( .A1(n737), .A2(G8), .ZN(n738) );
  XNOR2_X1 U831 ( .A(n738), .B(KEYINPUT30), .ZN(n739) );
  NOR2_X1 U832 ( .A1(n739), .A2(G168), .ZN(n742) );
  NOR2_X1 U833 ( .A1(G171), .A2(n740), .ZN(n741) );
  NOR2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n744) );
  INV_X1 U835 ( .A(KEYINPUT31), .ZN(n743) );
  XNOR2_X1 U836 ( .A(n744), .B(n743), .ZN(n745) );
  NAND2_X1 U837 ( .A1(n746), .A2(n745), .ZN(n756) );
  NAND2_X1 U838 ( .A1(G286), .A2(n756), .ZN(n753) );
  NOR2_X1 U839 ( .A1(G1971), .A2(n782), .ZN(n749) );
  NOR2_X1 U840 ( .A1(G2090), .A2(n747), .ZN(n748) );
  NOR2_X1 U841 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U842 ( .A(KEYINPUT93), .B(n750), .Z(n751) );
  NAND2_X1 U843 ( .A1(n751), .A2(G303), .ZN(n752) );
  NAND2_X1 U844 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U845 ( .A1(G8), .A2(n754), .ZN(n755) );
  XNOR2_X1 U846 ( .A(n755), .B(KEYINPUT32), .ZN(n771) );
  OR2_X1 U847 ( .A1(G1966), .A2(n782), .ZN(n757) );
  XNOR2_X1 U848 ( .A(n758), .B(KEYINPUT92), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n759), .A2(G8), .ZN(n760) );
  NAND2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n770) );
  NAND2_X1 U851 ( .A1(n771), .A2(n770), .ZN(n764) );
  NOR2_X1 U852 ( .A1(G2090), .A2(G303), .ZN(n762) );
  NAND2_X1 U853 ( .A1(G8), .A2(n762), .ZN(n763) );
  NAND2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n765), .A2(n782), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n788) );
  NAND2_X1 U857 ( .A1(G1976), .A2(G288), .ZN(n917) );
  INV_X1 U858 ( .A(n917), .ZN(n768) );
  OR2_X1 U859 ( .A1(n782), .A2(n768), .ZN(n775) );
  INV_X1 U860 ( .A(n775), .ZN(n769) );
  AND2_X1 U861 ( .A1(n770), .A2(n769), .ZN(n772) );
  NAND2_X1 U862 ( .A1(n772), .A2(n771), .ZN(n777) );
  NOR2_X1 U863 ( .A1(G1976), .A2(G288), .ZN(n918) );
  NOR2_X1 U864 ( .A1(G1971), .A2(G303), .ZN(n773) );
  NOR2_X1 U865 ( .A1(n918), .A2(n773), .ZN(n774) );
  OR2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U868 ( .A(n778), .B(KEYINPUT64), .ZN(n779) );
  NOR2_X1 U869 ( .A1(KEYINPUT33), .A2(n779), .ZN(n786) );
  NAND2_X1 U870 ( .A1(KEYINPUT33), .A2(n918), .ZN(n780) );
  XNOR2_X1 U871 ( .A(KEYINPUT94), .B(n780), .ZN(n781) );
  NOR2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U873 ( .A(KEYINPUT95), .B(n783), .ZN(n784) );
  XOR2_X1 U874 ( .A(G1981), .B(G305), .Z(n926) );
  NAND2_X1 U875 ( .A1(n784), .A2(n926), .ZN(n785) );
  NOR2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n792) );
  XNOR2_X1 U879 ( .A(G1986), .B(G290), .ZN(n909) );
  NAND2_X1 U880 ( .A1(n909), .A2(n804), .ZN(n791) );
  NAND2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n807) );
  NOR2_X1 U882 ( .A1(G1996), .A2(n873), .ZN(n995) );
  INV_X1 U883 ( .A(n793), .ZN(n796) );
  NOR2_X1 U884 ( .A1(G1986), .A2(G290), .ZN(n794) );
  NOR2_X1 U885 ( .A1(G1991), .A2(n889), .ZN(n986) );
  NOR2_X1 U886 ( .A1(n794), .A2(n986), .ZN(n795) );
  NOR2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U888 ( .A(n797), .B(KEYINPUT96), .ZN(n798) );
  NOR2_X1 U889 ( .A1(n995), .A2(n798), .ZN(n799) );
  XNOR2_X1 U890 ( .A(n799), .B(KEYINPUT39), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U892 ( .A1(n876), .A2(n802), .ZN(n992) );
  NAND2_X1 U893 ( .A1(n803), .A2(n992), .ZN(n805) );
  NAND2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n810) );
  XOR2_X1 U896 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n808) );
  XNOR2_X1 U897 ( .A(KEYINPUT40), .B(n808), .ZN(n809) );
  XNOR2_X1 U898 ( .A(n810), .B(n809), .ZN(G329) );
  XOR2_X1 U899 ( .A(KEYINPUT99), .B(G2451), .Z(n812) );
  XNOR2_X1 U900 ( .A(G2446), .B(G2427), .ZN(n811) );
  XNOR2_X1 U901 ( .A(n812), .B(n811), .ZN(n819) );
  XOR2_X1 U902 ( .A(G2438), .B(G2435), .Z(n814) );
  XNOR2_X1 U903 ( .A(G2443), .B(G2430), .ZN(n813) );
  XNOR2_X1 U904 ( .A(n814), .B(n813), .ZN(n815) );
  XOR2_X1 U905 ( .A(n815), .B(G2454), .Z(n817) );
  XNOR2_X1 U906 ( .A(G1341), .B(G1348), .ZN(n816) );
  XNOR2_X1 U907 ( .A(n817), .B(n816), .ZN(n818) );
  XNOR2_X1 U908 ( .A(n819), .B(n818), .ZN(n820) );
  NAND2_X1 U909 ( .A1(n820), .A2(G14), .ZN(n900) );
  XOR2_X1 U910 ( .A(KEYINPUT100), .B(n900), .Z(G401) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n906), .ZN(G217) );
  NAND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n821) );
  XNOR2_X1 U913 ( .A(KEYINPUT101), .B(n821), .ZN(n822) );
  NAND2_X1 U914 ( .A1(n822), .A2(G661), .ZN(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n823) );
  XNOR2_X1 U916 ( .A(KEYINPUT102), .B(n823), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n825), .A2(n824), .ZN(G188) );
  INV_X1 U919 ( .A(G132), .ZN(G219) );
  INV_X1 U920 ( .A(G108), .ZN(G238) );
  INV_X1 U921 ( .A(G82), .ZN(G220) );
  NOR2_X1 U922 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U923 ( .A(G325), .ZN(G261) );
  INV_X1 U924 ( .A(n828), .ZN(G319) );
  XOR2_X1 U925 ( .A(KEYINPUT43), .B(G2090), .Z(n830) );
  XNOR2_X1 U926 ( .A(G2067), .B(G2072), .ZN(n829) );
  XNOR2_X1 U927 ( .A(n830), .B(n829), .ZN(n841) );
  XOR2_X1 U928 ( .A(KEYINPUT42), .B(G2096), .Z(n832) );
  XNOR2_X1 U929 ( .A(G2678), .B(KEYINPUT106), .ZN(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(n837) );
  XNOR2_X1 U931 ( .A(KEYINPUT103), .B(n833), .ZN(n835) );
  XNOR2_X1 U932 ( .A(KEYINPUT105), .B(KEYINPUT104), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U934 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U935 ( .A(G2084), .B(G2078), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U937 ( .A(n841), .B(n840), .Z(G227) );
  XOR2_X1 U938 ( .A(G1956), .B(G1971), .Z(n843) );
  XNOR2_X1 U939 ( .A(G1996), .B(G1976), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n847) );
  XNOR2_X1 U941 ( .A(n950), .B(G1966), .ZN(n845) );
  XNOR2_X1 U942 ( .A(G1986), .B(G1981), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U944 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U945 ( .A(G2474), .B(KEYINPUT41), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U947 ( .A(KEYINPUT107), .B(n850), .ZN(n851) );
  XOR2_X1 U948 ( .A(n851), .B(G1991), .Z(G229) );
  NAND2_X1 U949 ( .A1(G136), .A2(n882), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n852), .B(KEYINPUT108), .ZN(n858) );
  NAND2_X1 U951 ( .A1(n878), .A2(G112), .ZN(n853) );
  XOR2_X1 U952 ( .A(KEYINPUT109), .B(n853), .Z(n855) );
  NAND2_X1 U953 ( .A1(n883), .A2(G100), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U955 ( .A(KEYINPUT110), .B(n856), .Z(n857) );
  NAND2_X1 U956 ( .A1(n858), .A2(n857), .ZN(n861) );
  NAND2_X1 U957 ( .A1(n879), .A2(G124), .ZN(n859) );
  XOR2_X1 U958 ( .A(KEYINPUT44), .B(n859), .Z(n860) );
  NOR2_X1 U959 ( .A1(n861), .A2(n860), .ZN(G162) );
  XOR2_X1 U960 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n871) );
  NAND2_X1 U961 ( .A1(G139), .A2(n882), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G103), .A2(n883), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n868) );
  NAND2_X1 U964 ( .A1(G115), .A2(n878), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G127), .A2(n879), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U967 ( .A(KEYINPUT47), .B(n866), .Z(n867) );
  NOR2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U969 ( .A(KEYINPUT111), .B(n869), .Z(n999) );
  XNOR2_X1 U970 ( .A(n999), .B(n984), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U972 ( .A(G162), .B(n872), .ZN(n875) );
  XOR2_X1 U973 ( .A(G164), .B(n873), .Z(n874) );
  XNOR2_X1 U974 ( .A(n875), .B(n874), .ZN(n877) );
  XNOR2_X1 U975 ( .A(n877), .B(n876), .ZN(n893) );
  NAND2_X1 U976 ( .A1(G118), .A2(n878), .ZN(n881) );
  NAND2_X1 U977 ( .A1(G130), .A2(n879), .ZN(n880) );
  NAND2_X1 U978 ( .A1(n881), .A2(n880), .ZN(n888) );
  NAND2_X1 U979 ( .A1(G142), .A2(n882), .ZN(n885) );
  NAND2_X1 U980 ( .A1(G106), .A2(n883), .ZN(n884) );
  NAND2_X1 U981 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U982 ( .A(n886), .B(KEYINPUT45), .Z(n887) );
  NOR2_X1 U983 ( .A1(n888), .A2(n887), .ZN(n890) );
  XNOR2_X1 U984 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U985 ( .A(G160), .B(n891), .ZN(n892) );
  XNOR2_X1 U986 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U987 ( .A1(G37), .A2(n894), .ZN(G395) );
  XOR2_X1 U988 ( .A(n895), .B(G286), .Z(n897) );
  XOR2_X1 U989 ( .A(n907), .B(G301), .Z(n896) );
  XNOR2_X1 U990 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U991 ( .A1(n898), .A2(G37), .ZN(n899) );
  XNOR2_X1 U992 ( .A(n899), .B(KEYINPUT112), .ZN(G397) );
  NAND2_X1 U993 ( .A1(G319), .A2(n900), .ZN(n903) );
  NOR2_X1 U994 ( .A1(G227), .A2(G229), .ZN(n901) );
  XNOR2_X1 U995 ( .A(KEYINPUT49), .B(n901), .ZN(n902) );
  NOR2_X1 U996 ( .A1(n903), .A2(n902), .ZN(n905) );
  NOR2_X1 U997 ( .A1(G395), .A2(G397), .ZN(n904) );
  NAND2_X1 U998 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U999 ( .A(G225), .ZN(G308) );
  INV_X1 U1000 ( .A(G96), .ZN(G221) );
  INV_X1 U1001 ( .A(G69), .ZN(G235) );
  INV_X1 U1002 ( .A(n906), .ZN(G223) );
  XNOR2_X1 U1003 ( .A(G16), .B(KEYINPUT56), .ZN(n932) );
  XOR2_X1 U1004 ( .A(n907), .B(G1348), .Z(n908) );
  NOR2_X1 U1005 ( .A1(n909), .A2(n908), .ZN(n915) );
  XOR2_X1 U1006 ( .A(G1341), .B(KEYINPUT119), .Z(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n913) );
  XOR2_X1 U1008 ( .A(G301), .B(n950), .Z(n912) );
  NOR2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(n925) );
  XOR2_X1 U1011 ( .A(G1956), .B(G299), .Z(n916) );
  NAND2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(n922) );
  XNOR2_X1 U1013 ( .A(n918), .B(KEYINPUT117), .ZN(n920) );
  XOR2_X1 U1014 ( .A(G303), .B(G1971), .Z(n919) );
  NAND2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1017 ( .A(KEYINPUT118), .B(n923), .Z(n924) );
  NOR2_X1 U1018 ( .A1(n925), .A2(n924), .ZN(n930) );
  XNOR2_X1 U1019 ( .A(G1966), .B(G168), .ZN(n927) );
  NAND2_X1 U1020 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1021 ( .A(n928), .B(KEYINPUT57), .ZN(n929) );
  NAND2_X1 U1022 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1023 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1024 ( .A(KEYINPUT120), .B(n933), .ZN(n1014) );
  XOR2_X1 U1025 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n943) );
  XNOR2_X1 U1026 ( .A(G1341), .B(G19), .ZN(n935) );
  XNOR2_X1 U1027 ( .A(G1956), .B(G20), .ZN(n934) );
  NOR2_X1 U1028 ( .A1(n935), .A2(n934), .ZN(n941) );
  XOR2_X1 U1029 ( .A(KEYINPUT122), .B(G4), .Z(n937) );
  XNOR2_X1 U1030 ( .A(G1348), .B(KEYINPUT59), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(n937), .B(n936), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(G1981), .B(G6), .ZN(n938) );
  NOR2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1035 ( .A(n943), .B(n942), .ZN(n956) );
  XNOR2_X1 U1036 ( .A(G1976), .B(G23), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(G1971), .B(G22), .ZN(n944) );
  NOR2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n947) );
  XOR2_X1 U1039 ( .A(G1986), .B(G24), .Z(n946) );
  NAND2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n949) );
  XOR2_X1 U1041 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n948) );
  XNOR2_X1 U1042 ( .A(n949), .B(n948), .ZN(n954) );
  XNOR2_X1 U1043 ( .A(G1966), .B(G21), .ZN(n952) );
  XOR2_X1 U1044 ( .A(n950), .B(G5), .Z(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1046 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1047 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1048 ( .A(KEYINPUT61), .B(n957), .Z(n958) );
  XNOR2_X1 U1049 ( .A(n958), .B(KEYINPUT125), .ZN(n960) );
  XNOR2_X1 U1050 ( .A(G16), .B(KEYINPUT121), .ZN(n959) );
  NAND2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1052 ( .A1(G11), .A2(n961), .ZN(n1012) );
  XOR2_X1 U1053 ( .A(G2090), .B(G35), .Z(n978) );
  XOR2_X1 U1054 ( .A(G2072), .B(G33), .Z(n962) );
  NAND2_X1 U1055 ( .A1(n962), .A2(G28), .ZN(n974) );
  XNOR2_X1 U1056 ( .A(G25), .B(G1991), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(n963), .B(KEYINPUT113), .ZN(n972) );
  XNOR2_X1 U1058 ( .A(G2067), .B(G26), .ZN(n970) );
  XNOR2_X1 U1059 ( .A(G1996), .B(G32), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(n964), .B(KEYINPUT114), .ZN(n967) );
  XOR2_X1 U1061 ( .A(G27), .B(n965), .Z(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n968), .B(KEYINPUT115), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1067 ( .A(KEYINPUT116), .B(n975), .Z(n976) );
  XNOR2_X1 U1068 ( .A(n976), .B(KEYINPUT53), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G34), .B(G2084), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(KEYINPUT54), .B(n979), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1073 ( .A1(G29), .A2(n982), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(n983), .B(KEYINPUT55), .ZN(n1010) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n989) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n991) );
  XOR2_X1 U1078 ( .A(G160), .B(G2084), .Z(n990) );
  NOR2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n993) );
  NAND2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n998) );
  XOR2_X1 U1081 ( .A(G2090), .B(G162), .Z(n994) );
  NOR2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(n996), .B(KEYINPUT51), .ZN(n997) );
  NOR2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n1006) );
  XOR2_X1 U1085 ( .A(G2072), .B(n999), .Z(n1001) );
  XOR2_X1 U1086 ( .A(G164), .B(G2078), .Z(n1000) );
  NOR2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1088 ( .A(KEYINPUT50), .B(n1002), .Z(n1003) );
  NOR2_X1 U1089 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1090 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1091 ( .A(KEYINPUT52), .B(n1007), .ZN(n1008) );
  NAND2_X1 U1092 ( .A1(G29), .A2(n1008), .ZN(n1009) );
  NAND2_X1 U1093 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1094 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1095 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1096 ( .A(KEYINPUT62), .B(n1015), .Z(G311) );
  XOR2_X1 U1097 ( .A(KEYINPUT126), .B(G311), .Z(G150) );
  INV_X1 U1098 ( .A(G303), .ZN(G166) );
endmodule

