//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT78), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT78), .ZN(new_n189));
  INV_X1    g003(.A(G113), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G122), .ZN(new_n191));
  INV_X1    g005(.A(G122), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G113), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n189), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT77), .B(G104), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n188), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n195), .B1(new_n188), .B2(new_n194), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G125), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(new_n202), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT18), .A2(G131), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(G237), .A2(G953), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n210), .A2(G143), .A3(G214), .ZN(new_n211));
  AOI21_X1  g025(.A(G143), .B1(new_n210), .B2(G214), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G237), .ZN(new_n214));
  INV_X1    g028(.A(G953), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G214), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n210), .A2(G143), .A3(G214), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(new_n208), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n207), .A2(new_n213), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT65), .B(G131), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n211), .B2(new_n212), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT17), .ZN(new_n224));
  AND2_X1   g038(.A1(KEYINPUT65), .A2(G131), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT65), .A2(G131), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n218), .A2(new_n227), .A3(new_n219), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n223), .A2(new_n224), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n200), .A2(new_n202), .A3(KEYINPUT16), .ZN(new_n230));
  OR3_X1    g044(.A1(new_n201), .A2(KEYINPUT16), .A3(G140), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n205), .ZN(new_n233));
  OAI211_X1 g047(.A(KEYINPUT17), .B(new_n222), .C1(new_n211), .C2(new_n212), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(new_n231), .A3(G146), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n198), .B(new_n221), .C1(new_n229), .C2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n207), .A2(new_n213), .A3(new_n220), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n223), .A2(new_n224), .A3(new_n228), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT79), .B1(new_n242), .B2(new_n198), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n221), .B1(new_n229), .B2(new_n236), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT79), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n244), .B(new_n245), .C1(new_n196), .C2(new_n197), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n238), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(G475), .B1(new_n247), .B2(G902), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n223), .A2(new_n228), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n200), .A2(new_n202), .A3(KEYINPUT19), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT19), .B1(new_n200), .B2(new_n202), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n205), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n235), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n198), .B1(new_n253), .B2(new_n221), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(new_n242), .B2(new_n198), .ZN(new_n255));
  NOR2_X1   g069(.A1(G475), .A2(G902), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT20), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n253), .A2(new_n221), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n237), .B1(new_n259), .B2(new_n198), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT20), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(new_n256), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n248), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT13), .ZN(new_n266));
  INV_X1    g080(.A(G128), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(G143), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n217), .A2(KEYINPUT13), .A3(G128), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(G143), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G134), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n217), .A2(G128), .ZN(new_n274));
  INV_X1    g088(.A(G134), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n270), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n192), .A2(G116), .ZN(new_n277));
  INV_X1    g091(.A(G116), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G122), .ZN(new_n279));
  INV_X1    g093(.A(G107), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n280), .B1(new_n277), .B2(new_n279), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n276), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(G116), .B(G122), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n280), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n274), .A2(new_n270), .A3(new_n275), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n275), .B1(new_n274), .B2(new_n270), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n278), .A2(KEYINPUT14), .A3(G122), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G107), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT14), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n290), .B1(new_n291), .B2(new_n284), .ZN(new_n292));
  OAI22_X1  g106(.A1(new_n273), .A2(new_n283), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT9), .B(G234), .ZN(new_n294));
  INV_X1    g108(.A(G217), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n294), .A2(new_n295), .A3(G953), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n272), .B(new_n276), .C1(new_n282), .C2(new_n281), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n299), .B(new_n296), .C1(new_n292), .C2(new_n288), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n300), .A3(KEYINPUT80), .ZN(new_n301));
  INV_X1    g115(.A(G902), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT80), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n293), .A2(new_n303), .A3(new_n297), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G478), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(KEYINPUT15), .ZN(new_n307));
  OR2_X1    g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n215), .A2(G952), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(G234), .B2(G237), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT21), .B(G898), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(G234), .A2(G237), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(G902), .A3(G953), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  XOR2_X1   g130(.A(new_n316), .B(KEYINPUT81), .Z(new_n317));
  NAND2_X1  g131(.A1(new_n305), .A2(new_n307), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n308), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n265), .A2(new_n320), .A3(KEYINPUT82), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT82), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(new_n264), .B2(new_n319), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G469), .ZN(new_n325));
  INV_X1    g139(.A(G104), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT3), .B1(new_n326), .B2(G107), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n280), .A3(G104), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(G107), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G101), .ZN(new_n332));
  INV_X1    g146(.A(G101), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n327), .A2(new_n329), .A3(new_n333), .A4(new_n330), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(KEYINPUT4), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n205), .A2(G143), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n217), .A2(G146), .ZN(new_n337));
  AND2_X1   g151(.A1(KEYINPUT0), .A2(G128), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT64), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(new_n217), .B2(G146), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n205), .A2(KEYINPUT64), .A3(G143), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n336), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(KEYINPUT0), .A2(G128), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n338), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n340), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n333), .A2(KEYINPUT4), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n331), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n335), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT11), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(new_n275), .B2(G137), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n275), .A2(G137), .ZN(new_n353));
  INV_X1    g167(.A(G137), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(KEYINPUT11), .A3(G134), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G131), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n227), .A2(new_n353), .A3(new_n352), .A4(new_n355), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n280), .A2(G104), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n326), .A2(G107), .ZN(new_n362));
  OAI21_X1  g176(.A(G101), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT1), .B1(new_n217), .B2(G146), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n364), .A2(G128), .B1(new_n336), .B2(new_n337), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n267), .A2(KEYINPUT1), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n366), .A2(new_n336), .A3(new_n337), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n334), .B(new_n363), .C1(new_n365), .C2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n334), .A2(new_n363), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n366), .A2(new_n336), .A3(new_n337), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n217), .A2(G146), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT64), .B1(new_n205), .B2(G143), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n341), .A2(new_n217), .A3(G146), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n267), .B1(new_n336), .B2(KEYINPUT1), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n372), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n371), .A2(new_n378), .A3(KEYINPUT10), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n350), .A2(new_n360), .A3(new_n370), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n215), .A2(G227), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT71), .ZN(new_n382));
  XNOR2_X1  g196(.A(G110), .B(G140), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n368), .B1(new_n378), .B2(new_n371), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT12), .A3(new_n359), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n359), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT12), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n385), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n350), .A2(new_n370), .A3(new_n379), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n359), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n384), .B1(new_n393), .B2(new_n380), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n325), .B(new_n302), .C1(new_n391), .C2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n385), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n393), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n350), .A2(new_n370), .A3(new_n379), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n387), .A2(new_n390), .B1(new_n398), .B2(new_n360), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n397), .B(G469), .C1(new_n399), .C2(new_n384), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n325), .A2(new_n302), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n395), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G221), .ZN(new_n404));
  INV_X1    g218(.A(new_n294), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n302), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G214), .B1(G237), .B2(G902), .ZN(new_n410));
  XOR2_X1   g224(.A(new_n410), .B(KEYINPUT72), .Z(new_n411));
  INV_X1    g225(.A(G224), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(G953), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT7), .ZN(new_n415));
  INV_X1    g229(.A(new_n346), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n339), .B1(new_n376), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n415), .B1(new_n417), .B2(G125), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n201), .B(new_n372), .C1(new_n376), .C2(new_n377), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT75), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n419), .A2(new_n420), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n418), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n190), .A2(KEYINPUT2), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT2), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G113), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G116), .B(G119), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G119), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G116), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n278), .A2(G119), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT5), .ZN(new_n433));
  OAI21_X1  g247(.A(G113), .B1(new_n431), .B2(KEYINPUT5), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n429), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n334), .A2(new_n363), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n278), .A2(G119), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT5), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n190), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT5), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n442), .A2(new_n429), .A3(new_n334), .A4(new_n363), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G110), .B(G122), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT8), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n423), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n377), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n344), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n450), .A2(KEYINPUT75), .A3(new_n201), .A4(new_n372), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n419), .A2(new_n420), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n417), .A2(G125), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n453), .A2(new_n454), .B1(KEYINPUT7), .B2(new_n414), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT76), .B1(new_n448), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT74), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n431), .A2(new_n432), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n424), .A3(new_n426), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n459), .A2(new_n429), .B1(new_n331), .B2(new_n348), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n440), .A2(new_n441), .B1(new_n428), .B2(new_n427), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n335), .A2(new_n460), .B1(new_n371), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n457), .B1(new_n462), .B2(new_n445), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n457), .A3(new_n445), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n454), .B1(new_n421), .B2(new_n422), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n415), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT76), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n453), .A2(new_n418), .B1(new_n444), .B2(new_n446), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n456), .A2(new_n466), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n335), .A2(new_n460), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n443), .ZN(new_n475));
  XOR2_X1   g289(.A(new_n445), .B(KEYINPUT73), .Z(new_n476));
  AOI21_X1  g290(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n462), .A2(new_n457), .A3(new_n445), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n477), .B1(new_n478), .B2(new_n463), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n467), .A2(new_n413), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n453), .A2(new_n454), .A3(new_n414), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n475), .A2(new_n473), .A3(new_n476), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n479), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n472), .A2(new_n302), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G210), .B1(G237), .B2(G902), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n472), .A2(new_n484), .A3(new_n302), .A4(new_n486), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n411), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n324), .A2(new_n409), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT83), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G110), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n267), .A2(KEYINPUT23), .A3(G119), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n430), .A2(G128), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n430), .A2(G128), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n495), .B(new_n496), .C1(new_n497), .C2(KEYINPUT23), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n494), .B1(new_n498), .B2(KEYINPUT69), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(KEYINPUT69), .B2(new_n498), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n233), .A2(new_n235), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n267), .A2(G119), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT24), .B(G110), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n500), .B(new_n501), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n504), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(new_n498), .B2(G110), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n235), .A3(new_n206), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n508), .A2(KEYINPUT70), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(KEYINPUT70), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT22), .B(G137), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n215), .A2(G221), .A3(G234), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n514), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n505), .B(new_n516), .C1(new_n509), .C2(new_n510), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n295), .B1(G234), .B2(new_n302), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(G902), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n518), .B2(G902), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n515), .A2(KEYINPUT25), .A3(new_n302), .A4(new_n517), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n522), .B1(new_n526), .B2(new_n519), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT68), .B(KEYINPUT32), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n459), .A2(new_n429), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n347), .A2(new_n359), .ZN(new_n531));
  INV_X1    g345(.A(G131), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n354), .A2(G134), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n532), .B1(new_n353), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(new_n227), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n378), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n531), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n538), .B1(new_n531), .B2(new_n537), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n530), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  XOR2_X1   g355(.A(KEYINPUT66), .B(KEYINPUT27), .Z(new_n542));
  NAND2_X1  g356(.A1(new_n210), .A2(G210), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT26), .B(G101), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n359), .A2(new_n347), .B1(new_n536), .B2(new_n378), .ZN(new_n547));
  INV_X1    g361(.A(new_n530), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n541), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT31), .ZN(new_n551));
  INV_X1    g365(.A(new_n546), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n531), .A2(new_n537), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT67), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n530), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n547), .A2(KEYINPUT67), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT28), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT28), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n553), .A2(new_n530), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n559), .B2(new_n549), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n552), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT31), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n541), .A2(new_n562), .A3(new_n546), .A4(new_n549), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n551), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(G472), .A2(G902), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n529), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n565), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n548), .B1(new_n547), .B2(KEYINPUT67), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n553), .A2(new_n554), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n558), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n553), .A2(new_n530), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n547), .A2(new_n548), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT28), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n574), .A2(new_n552), .B1(new_n550), .B2(KEYINPUT31), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n567), .B1(new_n575), .B2(new_n563), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n566), .B1(KEYINPUT32), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n570), .A2(new_n573), .A3(KEYINPUT29), .A4(new_n546), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT29), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n553), .A2(KEYINPUT30), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n547), .A2(new_n538), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n571), .B1(new_n582), .B2(new_n530), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n579), .B1(new_n583), .B2(new_n546), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n557), .A2(new_n560), .A3(new_n552), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n302), .B(new_n578), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G472), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n528), .B1(new_n577), .B2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n324), .A2(KEYINPUT83), .A3(new_n409), .A4(new_n490), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n493), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  INV_X1    g405(.A(new_n410), .ZN(new_n592));
  INV_X1    g406(.A(new_n489), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT84), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n488), .A2(KEYINPUT84), .A3(new_n489), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n301), .A2(new_n598), .A3(new_n304), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n298), .A2(new_n300), .A3(KEYINPUT33), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n306), .A2(G902), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT85), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n305), .A2(new_n306), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT85), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n599), .A2(new_n605), .A3(new_n600), .A4(new_n601), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n264), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT86), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT86), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n607), .A2(new_n264), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n597), .A2(new_n317), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n564), .A2(new_n302), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n576), .B1(G472), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n527), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n408), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT34), .B(G104), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  AOI21_X1  g434(.A(new_n264), .B1(new_n318), .B2(new_n308), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n595), .A2(new_n596), .A3(new_n621), .A4(new_n317), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n622), .A2(new_n616), .A3(new_n408), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT35), .B(G107), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G9));
  NAND2_X1  g439(.A1(new_n614), .A2(G472), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n564), .A2(new_n565), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n514), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n511), .B(new_n629), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n526), .A2(new_n519), .B1(new_n520), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n493), .A2(new_n589), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT37), .B(G110), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G12));
  NAND2_X1  g449(.A1(new_n308), .A2(new_n318), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n311), .B1(new_n315), .B2(G900), .ZN(new_n637));
  AND4_X1   g451(.A1(new_n248), .A2(new_n636), .A3(new_n263), .A4(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n595), .A2(new_n596), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT87), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT87), .A4(new_n638), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n529), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n627), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n564), .A2(KEYINPUT32), .A3(new_n565), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n587), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n631), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(new_n409), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  NOR2_X1   g466(.A1(new_n571), .A2(new_n572), .ZN(new_n653));
  AOI21_X1  g467(.A(G902), .B1(new_n653), .B2(new_n552), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n583), .A2(new_n552), .ZN(new_n656));
  OAI21_X1  g470(.A(G472), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n577), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT40), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n637), .B(KEYINPUT39), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n408), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n659), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n660), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n264), .A2(new_n636), .ZN(new_n666));
  NOR4_X1   g480(.A1(new_n665), .A2(new_n592), .A3(new_n648), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n488), .A2(new_n489), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT38), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n664), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G143), .ZN(G45));
  AND3_X1   g485(.A1(new_n607), .A2(new_n264), .A3(new_n637), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n595), .A2(new_n672), .A3(new_n596), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT88), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n595), .A2(new_n672), .A3(new_n596), .A4(KEYINPUT88), .ZN(new_n676));
  AOI211_X1 g490(.A(KEYINPUT89), .B(new_n649), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT89), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n678), .B1(new_n679), .B2(new_n650), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n205), .ZN(G48));
  NAND3_X1  g496(.A1(new_n597), .A2(new_n317), .A3(new_n612), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n393), .A2(new_n380), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n390), .A2(new_n387), .ZN(new_n685));
  OAI22_X1  g499(.A1(new_n684), .A2(new_n384), .B1(new_n685), .B2(new_n385), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n325), .B1(new_n686), .B2(new_n302), .ZN(new_n687));
  INV_X1    g501(.A(new_n395), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n687), .A2(new_n688), .A3(new_n406), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n647), .A2(new_n527), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n683), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT41), .B(G113), .Z(new_n692));
  XOR2_X1   g506(.A(new_n692), .B(KEYINPUT90), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n691), .B(new_n693), .ZN(G15));
  NOR2_X1   g508(.A1(new_n690), .A2(new_n622), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n278), .ZN(G18));
  NAND2_X1  g510(.A1(new_n597), .A2(new_n689), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n324), .A2(new_n647), .A3(new_n648), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n430), .ZN(G21));
  NAND4_X1  g514(.A1(new_n615), .A2(new_n689), .A3(new_n527), .A4(new_n317), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n595), .A2(new_n596), .A3(new_n264), .A4(new_n636), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n192), .ZN(G24));
  NAND2_X1  g518(.A1(new_n595), .A2(new_n596), .ZN(new_n705));
  INV_X1    g519(.A(new_n689), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT91), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n708), .B1(new_n628), .B2(new_n631), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n615), .A2(new_n648), .A3(KEYINPUT91), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n707), .A2(new_n709), .A3(new_n672), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G125), .ZN(G27));
  INV_X1    g526(.A(KEYINPUT92), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n403), .A2(new_n713), .A3(new_n407), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n488), .A2(new_n489), .A3(new_n410), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n713), .B1(new_n403), .B2(new_n407), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n672), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT42), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI22_X1  g534(.A1(new_n646), .A2(KEYINPUT94), .B1(new_n586), .B2(G472), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT95), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(new_n576), .B2(KEYINPUT32), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT32), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n627), .A2(KEYINPUT95), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT94), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n576), .A2(new_n726), .A3(KEYINPUT32), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n721), .A2(new_n723), .A3(new_n725), .A4(new_n727), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n728), .A2(KEYINPUT96), .A3(new_n527), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT96), .B1(new_n728), .B2(new_n527), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n717), .B(new_n720), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n588), .A2(new_n672), .A3(new_n717), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT93), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n732), .A2(new_n733), .A3(new_n719), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n733), .B1(new_n732), .B2(new_n719), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n731), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G131), .ZN(G33));
  NAND2_X1  g551(.A1(new_n588), .A2(new_n717), .ZN(new_n738));
  INV_X1    g552(.A(new_n638), .ZN(new_n739));
  OR3_X1    g553(.A1(new_n738), .A2(KEYINPUT97), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT97), .B1(new_n738), .B2(new_n739), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  INV_X1    g557(.A(KEYINPUT101), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n264), .B(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(KEYINPUT43), .A3(new_n607), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n265), .A2(new_n607), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n615), .A2(new_n631), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(KEYINPUT102), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n715), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n753), .B(new_n754), .C1(new_n752), .C2(new_n751), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT102), .B1(new_n751), .B2(new_n752), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n399), .A2(new_n384), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n397), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n325), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n759), .A2(KEYINPUT45), .A3(new_n397), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT98), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT98), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n762), .A2(new_n766), .A3(new_n763), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(KEYINPUT99), .B(new_n758), .C1(new_n768), .C2(new_n401), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT99), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n401), .B1(new_n765), .B2(new_n767), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n770), .B1(new_n771), .B2(KEYINPUT46), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n688), .B1(new_n771), .B2(KEYINPUT46), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n769), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n407), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n662), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n757), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(KEYINPUT103), .B(G137), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT104), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n777), .B(new_n779), .ZN(G39));
  NOR4_X1   g594(.A1(new_n647), .A2(new_n718), .A3(new_n527), .A4(new_n715), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n774), .A2(KEYINPUT47), .A3(new_n407), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT47), .B1(new_n774), .B2(new_n407), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  OR2_X1    g600(.A1(G952), .A2(G953), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n732), .A2(new_n719), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT93), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n732), .A2(new_n733), .A3(new_n719), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI22_X1  g605(.A1(new_n791), .A2(new_n731), .B1(new_n740), .B2(new_n741), .ZN(new_n792));
  OAI22_X1  g606(.A1(new_n683), .A2(new_n690), .B1(new_n701), .B2(new_n702), .ZN(new_n793));
  OAI22_X1  g607(.A1(new_n697), .A2(new_n698), .B1(new_n690), .B2(new_n622), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n608), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n490), .A2(new_n317), .A3(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT105), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n308), .A2(KEYINPUT106), .A3(new_n318), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT106), .B1(new_n308), .B2(new_n318), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n490), .A2(new_n265), .A3(new_n317), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n797), .A2(new_n798), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n617), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n493), .B(new_n589), .C1(new_n632), .C2(new_n588), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n248), .A2(new_n263), .A3(new_n637), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT107), .B1(new_n803), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT106), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n636), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n800), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT107), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n814), .A3(new_n265), .A4(new_n637), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n810), .A2(new_n754), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n649), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n709), .A2(new_n672), .A3(new_n710), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n817), .B1(new_n818), .B2(new_n717), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n795), .A2(new_n807), .A3(new_n808), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n822));
  INV_X1    g636(.A(new_n702), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n631), .A2(new_n637), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n409), .A3(new_n658), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n651), .A2(new_n825), .A3(new_n711), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n681), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n679), .A2(new_n650), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT89), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n679), .A2(new_n678), .A3(new_n650), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n651), .A2(new_n711), .A3(new_n825), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n792), .B(new_n821), .C1(new_n827), .C2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n736), .A2(new_n742), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n836), .A2(new_n835), .A3(new_n820), .ZN(new_n837));
  OAI211_X1 g651(.A(KEYINPUT109), .B(new_n822), .C1(new_n681), .C2(new_n826), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT109), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n831), .B2(new_n832), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n838), .B1(new_n840), .B2(new_n822), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n834), .A2(new_n835), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT112), .ZN(new_n843));
  XNOR2_X1  g657(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n843), .B1(new_n842), .B2(new_n844), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT110), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n792), .A2(new_n821), .A3(KEYINPUT108), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT108), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n836), .B2(new_n820), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n841), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n835), .ZN(new_n853));
  INV_X1    g667(.A(new_n834), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT53), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n848), .B1(new_n856), .B2(KEYINPUT54), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  AOI211_X1 g672(.A(KEYINPUT110), .B(new_n858), .C1(new_n853), .C2(new_n855), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n847), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n749), .A2(new_n310), .ZN(new_n861));
  INV_X1    g675(.A(new_n616), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n715), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT113), .ZN(new_n865));
  INV_X1    g679(.A(new_n784), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n782), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n687), .A2(new_n688), .A3(new_n407), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n870), .B(KEYINPUT115), .Z(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n867), .A2(new_n868), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n865), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n706), .A2(new_n715), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n861), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n709), .A2(new_n710), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n659), .A2(new_n875), .A3(new_n527), .A4(new_n310), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n607), .A2(new_n264), .ZN(new_n879));
  OAI22_X1  g693(.A1(new_n876), .A2(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n669), .A2(new_n410), .A3(new_n706), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n863), .A2(new_n882), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n883), .A2(KEYINPUT50), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(KEYINPUT50), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT51), .B1(new_n874), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n865), .B1(new_n867), .B2(new_n870), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n888), .A2(KEYINPUT51), .A3(new_n886), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n729), .A2(new_n730), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n861), .A3(new_n875), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT48), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n863), .A2(new_n697), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n309), .B(KEYINPUT116), .Z(new_n894));
  AOI21_X1  g708(.A(new_n878), .B1(new_n609), .B2(new_n611), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n892), .A2(KEYINPUT117), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT117), .B1(new_n892), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n889), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n887), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n787), .B1(new_n860), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n687), .A2(new_n688), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT49), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n745), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n406), .A2(new_n411), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n527), .A2(new_n607), .A3(new_n905), .ZN(new_n906));
  OR4_X1    g720(.A1(new_n669), .A2(new_n904), .A3(new_n658), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n901), .A2(new_n907), .ZN(G75));
  NOR2_X1   g722(.A1(new_n842), .A2(new_n302), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(G210), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT56), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n479), .A2(new_n483), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT118), .Z(new_n913));
  XNOR2_X1  g727(.A(new_n482), .B(KEYINPUT55), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n910), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n915), .B1(new_n910), .B2(new_n911), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n215), .A2(G952), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(G51));
  XOR2_X1   g733(.A(new_n842), .B(new_n844), .Z(new_n920));
  XOR2_X1   g734(.A(new_n401), .B(KEYINPUT57), .Z(new_n921));
  OAI21_X1  g735(.A(new_n686), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n909), .A2(new_n768), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n918), .B1(new_n922), .B2(new_n923), .ZN(G54));
  INV_X1    g738(.A(new_n918), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n909), .A2(KEYINPUT58), .A3(G475), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(new_n260), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n260), .B2(new_n926), .ZN(G60));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT59), .Z(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n599), .A2(new_n600), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n925), .B1(new_n920), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n860), .A2(new_n931), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n599), .A2(new_n600), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(G63));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT60), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT119), .B1(new_n842), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT119), .ZN(new_n940));
  INV_X1    g754(.A(new_n938), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n837), .A2(new_n841), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n836), .A2(new_n820), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n822), .B1(new_n681), .B2(new_n826), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT52), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT53), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n940), .B(new_n941), .C1(new_n942), .C2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n939), .A2(new_n518), .A3(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n949), .A2(new_n925), .ZN(new_n950));
  INV_X1    g764(.A(new_n630), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n939), .B2(new_n948), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n950), .B(new_n953), .C1(KEYINPUT120), .C2(KEYINPUT61), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n949), .A2(KEYINPUT120), .A3(new_n925), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n949), .A2(new_n925), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n955), .B(new_n956), .C1(new_n957), .C2(new_n952), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n954), .A2(new_n958), .ZN(G66));
  OAI21_X1  g773(.A(G953), .B1(new_n312), .B2(new_n412), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT121), .ZN(new_n961));
  INV_X1    g775(.A(new_n793), .ZN(new_n962));
  INV_X1    g776(.A(new_n794), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n962), .A2(new_n963), .A3(new_n807), .A4(new_n808), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n961), .B1(new_n965), .B2(G953), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n913), .B1(G898), .B2(new_n215), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G69));
  OR2_X1    g782(.A1(new_n250), .A2(new_n251), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n582), .B(new_n969), .Z(new_n970));
  NAND3_X1  g784(.A1(new_n776), .A2(new_n823), .A3(new_n890), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n777), .A2(new_n785), .A3(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n651), .B(new_n711), .C1(new_n677), .C2(new_n680), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT122), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT123), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(new_n836), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n792), .A2(KEYINPUT123), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n972), .A2(new_n976), .A3(KEYINPUT124), .A4(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT124), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n973), .B(KEYINPUT122), .Z(new_n980));
  NAND2_X1  g794(.A1(new_n836), .A2(new_n975), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n980), .A2(new_n977), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n777), .A2(new_n785), .A3(new_n971), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n978), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n215), .ZN(new_n986));
  INV_X1    g800(.A(G227), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n987), .A2(G900), .A3(G953), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n970), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n980), .A2(new_n670), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT62), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT62), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n980), .A2(new_n993), .A3(new_n670), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n608), .B1(new_n813), .B2(new_n264), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n588), .A2(new_n663), .A3(new_n754), .A4(new_n995), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n777), .A2(new_n785), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n992), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n990), .B1(new_n998), .B2(G953), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n989), .B1(new_n970), .B2(new_n999), .ZN(G72));
  NAND4_X1  g814(.A1(new_n992), .A2(new_n965), .A3(new_n994), .A4(new_n997), .ZN(new_n1001));
  XNOR2_X1  g815(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1002));
  NAND2_X1  g816(.A1(G472), .A2(G902), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n656), .ZN(new_n1006));
  INV_X1    g820(.A(new_n656), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n583), .A2(new_n552), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n856), .A2(new_n1007), .A3(new_n1004), .A4(new_n1008), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1006), .A2(new_n925), .A3(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n978), .A2(new_n984), .A3(new_n965), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1011), .A2(KEYINPUT126), .A3(new_n1004), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1008), .B(KEYINPUT127), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1011), .A2(new_n1004), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT126), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1010), .B1(new_n1014), .B2(new_n1017), .ZN(G57));
endmodule


